
module table_parse_engine ( CLK, reset, boot_up, table_parse, input_valid, 
        glob_scen_noc_input_valid, delay_matrix_element, obj_id_element, 
        local_controller_id, calc_global_controller_prefetch_start, 
        calc_glob_dest_addr, tapping_loc_packet, calc_glob_prefetch_stop, 
        scenario_update, hardware_latency1, hardware_latency2, scenario_len, 
        prefetch_bypass_dest_addr_int, prefetch_bypass_cycles, 
        prefetch_bypass_start_addr );
  input [13:0] delay_matrix_element;
  input [1:0] obj_id_element;
  output [5:0] local_controller_id;
  output [7:0] calc_global_controller_prefetch_start;
  output [3:0] calc_glob_dest_addr;
  output [9:0] tapping_loc_packet;
  output [7:0] calc_glob_prefetch_stop;
  input [13:0] hardware_latency1;
  input [13:0] hardware_latency2;
  input [10:0] scenario_len;
  output [3:0] prefetch_bypass_dest_addr_int;
  output [7:0] prefetch_bypass_cycles;
  output [13:0] prefetch_bypass_start_addr;
  input CLK, reset, boot_up, table_parse, input_valid,
         glob_scen_noc_input_valid, scenario_update;
  wire   n2227, n2228, n2229, n2230, n2231, n2232, n2233, done, done2, N3860,
         N3861, N3862, N4190, N4191, N4192, N4193, N4194, N4195, N4196, N4197,
         N4198, N4199, N4200, N4201, N4202, N4203, N4204, N4205, N4206, N4207,
         N4208, N4209, N4210, N4211, N4212, N4213, N4214, N4215, N4216, N4217,
         N4218, N4219, N4220, N4221, N4222, N4223, N4224, N4225, N4226, N4227,
         N4228, N4229, N4230, N4231, N4232, N4233, N4234, N4235, N4236, N4237,
         N4238, N4239, N4240, N4241, N4242, N4243, N4244, N4245, N4246, N4247,
         N4248, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n809, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2220, n2225,
         n2226;
  wire   [1:0] table_ptr;
  wire   [7:0] obj_id;
  wire   [31:0] pointer;
  wire   [55:0] delay_matrix_N_1_next;
  wire   [7:0] obj_id_next;
  wire   [55:0] delay_matrix_N_1;
  wire   [31:0] copy_pointer;
  wire   [55:0] delay_matrix_N_1_next_original;
  wire   [55:0] delay_matrix_N_1_original;
  wire   [31:0] ptr_next;
  wire   [31:0] copy_ptr_next;
  wire   [1:0] group_header;
  wire   [7:0] calc_glob_controller_prefetch_start_int;
  wire   [5:0] local_controller_id_int;
  wire   [3:0] calc_glob_dest_addr_int;
  wire   [7:0] calc_glob_prefetch_stop_int;

  DFQD1BWP30P140LVT pointer_reg_31_ ( .D(n1148), .CP(CLK), .Q(pointer[31]) );
  DFQD1BWP30P140LVT pointer_reg_30_ ( .D(n1149), .CP(CLK), .Q(pointer[30]) );
  DFQD1BWP30P140LVT pointer_reg_29_ ( .D(n1150), .CP(CLK), .Q(pointer[29]) );
  DFQD1BWP30P140LVT pointer_reg_28_ ( .D(n1151), .CP(CLK), .Q(pointer[28]) );
  DFQD1BWP30P140LVT pointer_reg_27_ ( .D(n1152), .CP(CLK), .Q(pointer[27]) );
  DFQD1BWP30P140LVT pointer_reg_26_ ( .D(n1153), .CP(CLK), .Q(pointer[26]) );
  DFQD1BWP30P140LVT pointer_reg_25_ ( .D(n1154), .CP(CLK), .Q(pointer[25]) );
  DFQD1BWP30P140LVT pointer_reg_24_ ( .D(n1155), .CP(CLK), .Q(pointer[24]) );
  DFQD1BWP30P140LVT pointer_reg_23_ ( .D(n1156), .CP(CLK), .Q(pointer[23]) );
  DFQD1BWP30P140LVT pointer_reg_22_ ( .D(n1157), .CP(CLK), .Q(pointer[22]) );
  DFQD1BWP30P140LVT pointer_reg_21_ ( .D(n1158), .CP(CLK), .Q(pointer[21]) );
  DFQD1BWP30P140LVT pointer_reg_20_ ( .D(n1159), .CP(CLK), .Q(pointer[20]) );
  DFQD1BWP30P140LVT pointer_reg_19_ ( .D(n1160), .CP(CLK), .Q(pointer[19]) );
  DFQD1BWP30P140LVT pointer_reg_18_ ( .D(n1161), .CP(CLK), .Q(pointer[18]) );
  DFQD1BWP30P140LVT pointer_reg_17_ ( .D(n1162), .CP(CLK), .Q(pointer[17]) );
  DFQD1BWP30P140LVT pointer_reg_16_ ( .D(n1163), .CP(CLK), .Q(pointer[16]) );
  DFQD1BWP30P140LVT pointer_reg_15_ ( .D(n1164), .CP(CLK), .Q(pointer[15]) );
  DFQD1BWP30P140LVT pointer_reg_14_ ( .D(n1165), .CP(CLK), .Q(pointer[14]) );
  DFQD1BWP30P140LVT pointer_reg_13_ ( .D(n1166), .CP(CLK), .Q(pointer[13]) );
  DFQD1BWP30P140LVT pointer_reg_12_ ( .D(n1167), .CP(CLK), .Q(pointer[12]) );
  DFQD1BWP30P140LVT pointer_reg_11_ ( .D(n1168), .CP(CLK), .Q(pointer[11]) );
  DFQD1BWP30P140LVT pointer_reg_10_ ( .D(n1169), .CP(CLK), .Q(pointer[10]) );
  DFQD1BWP30P140LVT pointer_reg_9_ ( .D(n1170), .CP(CLK), .Q(pointer[9]) );
  DFQD1BWP30P140LVT pointer_reg_8_ ( .D(n1171), .CP(CLK), .Q(pointer[8]) );
  DFQD1BWP30P140LVT pointer_reg_7_ ( .D(n1172), .CP(CLK), .Q(pointer[7]) );
  DFQD1BWP30P140LVT pointer_reg_6_ ( .D(n1173), .CP(CLK), .Q(pointer[6]) );
  DFQD1BWP30P140LVT pointer_reg_5_ ( .D(n1174), .CP(CLK), .Q(pointer[5]) );
  DFQD1BWP30P140LVT pointer_reg_4_ ( .D(n1175), .CP(CLK), .Q(pointer[4]) );
  DFQD1BWP30P140LVT pointer_reg_3_ ( .D(n1176), .CP(CLK), .Q(pointer[3]) );
  DFQD1BWP30P140LVT pointer_reg_2_ ( .D(n1177), .CP(CLK), .Q(pointer[2]) );
  DFQD1BWP30P140LVT pointer_reg_1_ ( .D(n1178), .CP(CLK), .Q(pointer[1]) );
  DFQD1BWP30P140LVT pointer_reg_0_ ( .D(n1179), .CP(CLK), .Q(pointer[0]) );
  DFQD1BWP30P140LVT copy_pointer_reg_31_ ( .D(n1116), .CP(CLK), .Q(
        copy_pointer[31]) );
  DFQD1BWP30P140LVT copy_pointer_reg_30_ ( .D(n1117), .CP(CLK), .Q(
        copy_pointer[30]) );
  DFQD1BWP30P140LVT copy_pointer_reg_29_ ( .D(n1118), .CP(CLK), .Q(
        copy_pointer[29]) );
  DFQD1BWP30P140LVT copy_pointer_reg_28_ ( .D(n1119), .CP(CLK), .Q(
        copy_pointer[28]) );
  DFQD1BWP30P140LVT copy_pointer_reg_27_ ( .D(n1120), .CP(CLK), .Q(
        copy_pointer[27]) );
  DFQD1BWP30P140LVT copy_pointer_reg_26_ ( .D(n1121), .CP(CLK), .Q(
        copy_pointer[26]) );
  DFQD1BWP30P140LVT copy_pointer_reg_25_ ( .D(n1122), .CP(CLK), .Q(
        copy_pointer[25]) );
  DFQD1BWP30P140LVT copy_pointer_reg_24_ ( .D(n1123), .CP(CLK), .Q(
        copy_pointer[24]) );
  DFQD1BWP30P140LVT copy_pointer_reg_23_ ( .D(n1124), .CP(CLK), .Q(
        copy_pointer[23]) );
  DFQD1BWP30P140LVT copy_pointer_reg_22_ ( .D(n1125), .CP(CLK), .Q(
        copy_pointer[22]) );
  DFQD1BWP30P140LVT copy_pointer_reg_21_ ( .D(n1126), .CP(CLK), .Q(
        copy_pointer[21]) );
  DFQD1BWP30P140LVT copy_pointer_reg_20_ ( .D(n1127), .CP(CLK), .Q(
        copy_pointer[20]) );
  DFQD1BWP30P140LVT copy_pointer_reg_19_ ( .D(n1128), .CP(CLK), .Q(
        copy_pointer[19]) );
  DFQD1BWP30P140LVT copy_pointer_reg_18_ ( .D(n1129), .CP(CLK), .Q(
        copy_pointer[18]) );
  DFQD1BWP30P140LVT copy_pointer_reg_17_ ( .D(n1130), .CP(CLK), .Q(
        copy_pointer[17]) );
  DFQD1BWP30P140LVT copy_pointer_reg_16_ ( .D(n1131), .CP(CLK), .Q(
        copy_pointer[16]) );
  DFQD1BWP30P140LVT copy_pointer_reg_15_ ( .D(n1132), .CP(CLK), .Q(
        copy_pointer[15]) );
  DFQD1BWP30P140LVT copy_pointer_reg_14_ ( .D(n1133), .CP(CLK), .Q(
        copy_pointer[14]) );
  DFQD1BWP30P140LVT copy_pointer_reg_13_ ( .D(n1134), .CP(CLK), .Q(
        copy_pointer[13]) );
  DFQD1BWP30P140LVT copy_pointer_reg_12_ ( .D(n1135), .CP(CLK), .Q(
        copy_pointer[12]) );
  DFQD1BWP30P140LVT copy_pointer_reg_11_ ( .D(n1136), .CP(CLK), .Q(
        copy_pointer[11]) );
  DFQD1BWP30P140LVT copy_pointer_reg_10_ ( .D(n1137), .CP(CLK), .Q(
        copy_pointer[10]) );
  DFQD1BWP30P140LVT copy_pointer_reg_9_ ( .D(n1138), .CP(CLK), .Q(
        copy_pointer[9]) );
  DFQD1BWP30P140LVT copy_pointer_reg_8_ ( .D(n1139), .CP(CLK), .Q(
        copy_pointer[8]) );
  DFQD1BWP30P140LVT copy_pointer_reg_7_ ( .D(n1140), .CP(CLK), .Q(
        copy_pointer[7]) );
  DFQD1BWP30P140LVT copy_pointer_reg_6_ ( .D(n1141), .CP(CLK), .Q(
        copy_pointer[6]) );
  DFQD1BWP30P140LVT copy_pointer_reg_5_ ( .D(n1142), .CP(CLK), .Q(
        copy_pointer[5]) );
  DFQD1BWP30P140LVT copy_pointer_reg_4_ ( .D(n1143), .CP(CLK), .Q(
        copy_pointer[4]) );
  DFQD1BWP30P140LVT copy_pointer_reg_3_ ( .D(n1144), .CP(CLK), .Q(
        copy_pointer[3]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_3__13_ ( .D(n1070), .CP(CLK), 
        .Q(delay_matrix_N_1_next[55]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_3__13_ ( .D(n964), .CP(CLK), .Q(
        delay_matrix_N_1[55]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_3__12_ ( .D(n1071), .CP(CLK), 
        .Q(delay_matrix_N_1_next[54]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_3__12_ ( .D(n965), .CP(CLK), .Q(
        delay_matrix_N_1[54]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_3__11_ ( .D(n1072), .CP(CLK), 
        .Q(delay_matrix_N_1_next[53]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_3__11_ ( .D(n966), .CP(CLK), .Q(
        delay_matrix_N_1[53]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_3__10_ ( .D(n1073), .CP(CLK), 
        .Q(delay_matrix_N_1_next[52]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_3__10_ ( .D(n967), .CP(CLK), .Q(
        delay_matrix_N_1[52]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_3__9_ ( .D(n1074), .CP(CLK), .Q(
        delay_matrix_N_1_next[51]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_3__9_ ( .D(n968), .CP(CLK), .Q(
        delay_matrix_N_1[51]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_3__8_ ( .D(n1075), .CP(CLK), .Q(
        delay_matrix_N_1_next[50]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_3__8_ ( .D(n969), .CP(CLK), .Q(
        delay_matrix_N_1[50]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_3__7_ ( .D(n1076), .CP(CLK), .Q(
        delay_matrix_N_1_next[49]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_3__7_ ( .D(n970), .CP(CLK), .Q(
        delay_matrix_N_1[49]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_3__6_ ( .D(n1077), .CP(CLK), .Q(
        delay_matrix_N_1_next[48]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_3__6_ ( .D(n971), .CP(CLK), .Q(
        delay_matrix_N_1[48]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_3__5_ ( .D(n1078), .CP(CLK), .Q(
        delay_matrix_N_1_next[47]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_3__5_ ( .D(n972), .CP(CLK), .Q(
        delay_matrix_N_1[47]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_3__4_ ( .D(n1079), .CP(CLK), .Q(
        delay_matrix_N_1_next[46]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_3__4_ ( .D(n973), .CP(CLK), .Q(
        delay_matrix_N_1[46]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_3__3_ ( .D(n1080), .CP(CLK), .Q(
        delay_matrix_N_1_next[45]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_3__3_ ( .D(n974), .CP(CLK), .Q(
        delay_matrix_N_1[45]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_3__2_ ( .D(n1081), .CP(CLK), .Q(
        delay_matrix_N_1_next[44]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_3__2_ ( .D(n975), .CP(CLK), .Q(
        delay_matrix_N_1[44]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_3__1_ ( .D(n1082), .CP(CLK), .Q(
        delay_matrix_N_1_next[43]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_3__1_ ( .D(n976), .CP(CLK), .Q(
        delay_matrix_N_1[43]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_3__0_ ( .D(n1083), .CP(CLK), .Q(
        delay_matrix_N_1_next[42]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_3__0_ ( .D(n977), .CP(CLK), .Q(
        delay_matrix_N_1[42]) );
  DFQD1BWP30P140LVT obj_id_next_reg_3__1_ ( .D(n1054), .CP(CLK), .Q(
        obj_id_next[7]) );
  DFQD1BWP30P140LVT obj_id_reg_3__1_ ( .D(n956), .CP(CLK), .Q(obj_id[7]) );
  DFQD1BWP30P140LVT obj_id_next_reg_3__0_ ( .D(n1055), .CP(CLK), .Q(
        obj_id_next[6]) );
  DFQD1BWP30P140LVT obj_id_reg_3__0_ ( .D(n957), .CP(CLK), .Q(obj_id[6]) );
  DFQD1BWP30P140LVT ptr_next_reg_31_ ( .D(n1084), .CP(CLK), .Q(ptr_next[31])
         );
  DFQD1BWP30P140LVT ptr_next_reg_30_ ( .D(n1085), .CP(CLK), .Q(ptr_next[30])
         );
  DFQD1BWP30P140LVT ptr_next_reg_29_ ( .D(n1086), .CP(CLK), .Q(ptr_next[29])
         );
  DFQD1BWP30P140LVT ptr_next_reg_28_ ( .D(n1087), .CP(CLK), .Q(ptr_next[28])
         );
  DFQD1BWP30P140LVT ptr_next_reg_27_ ( .D(n1088), .CP(CLK), .Q(ptr_next[27])
         );
  DFQD1BWP30P140LVT ptr_next_reg_26_ ( .D(n1089), .CP(CLK), .Q(ptr_next[26])
         );
  DFQD1BWP30P140LVT ptr_next_reg_25_ ( .D(n1090), .CP(CLK), .Q(ptr_next[25])
         );
  DFQD1BWP30P140LVT ptr_next_reg_24_ ( .D(n1091), .CP(CLK), .Q(ptr_next[24])
         );
  DFQD1BWP30P140LVT ptr_next_reg_23_ ( .D(n1092), .CP(CLK), .Q(ptr_next[23])
         );
  DFQD1BWP30P140LVT ptr_next_reg_22_ ( .D(n1093), .CP(CLK), .Q(ptr_next[22])
         );
  DFQD1BWP30P140LVT ptr_next_reg_21_ ( .D(n1094), .CP(CLK), .Q(ptr_next[21])
         );
  DFQD1BWP30P140LVT ptr_next_reg_20_ ( .D(n1095), .CP(CLK), .Q(ptr_next[20])
         );
  DFQD1BWP30P140LVT ptr_next_reg_19_ ( .D(n1096), .CP(CLK), .Q(ptr_next[19])
         );
  DFQD1BWP30P140LVT ptr_next_reg_18_ ( .D(n1097), .CP(CLK), .Q(ptr_next[18])
         );
  DFQD1BWP30P140LVT ptr_next_reg_17_ ( .D(n1098), .CP(CLK), .Q(ptr_next[17])
         );
  DFQD1BWP30P140LVT ptr_next_reg_16_ ( .D(n1099), .CP(CLK), .Q(ptr_next[16])
         );
  DFQD1BWP30P140LVT ptr_next_reg_15_ ( .D(n1100), .CP(CLK), .Q(ptr_next[15])
         );
  DFQD1BWP30P140LVT ptr_next_reg_14_ ( .D(n1101), .CP(CLK), .Q(ptr_next[14])
         );
  DFQD1BWP30P140LVT ptr_next_reg_13_ ( .D(n1102), .CP(CLK), .Q(ptr_next[13])
         );
  DFQD1BWP30P140LVT ptr_next_reg_12_ ( .D(n1103), .CP(CLK), .Q(ptr_next[12])
         );
  DFQD1BWP30P140LVT ptr_next_reg_11_ ( .D(n1104), .CP(CLK), .Q(ptr_next[11])
         );
  DFQD1BWP30P140LVT ptr_next_reg_10_ ( .D(n1105), .CP(CLK), .Q(ptr_next[10])
         );
  DFQD1BWP30P140LVT ptr_next_reg_9_ ( .D(n1106), .CP(CLK), .Q(ptr_next[9]) );
  DFQD1BWP30P140LVT ptr_next_reg_8_ ( .D(n1107), .CP(CLK), .Q(ptr_next[8]) );
  DFQD1BWP30P140LVT ptr_next_reg_7_ ( .D(n1108), .CP(CLK), .Q(ptr_next[7]) );
  DFQD1BWP30P140LVT ptr_next_reg_6_ ( .D(n1109), .CP(CLK), .Q(ptr_next[6]) );
  DFQD1BWP30P140LVT ptr_next_reg_5_ ( .D(n1110), .CP(CLK), .Q(ptr_next[5]) );
  DFQD1BWP30P140LVT ptr_next_reg_4_ ( .D(n1111), .CP(CLK), .Q(ptr_next[4]) );
  DFQD1BWP30P140LVT ptr_next_reg_3_ ( .D(n1112), .CP(CLK), .Q(ptr_next[3]) );
  DFQD1BWP30P140LVT ptr_next_reg_2_ ( .D(n1113), .CP(CLK), .Q(ptr_next[2]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_2__0_ ( .D(n1069), .CP(CLK), .Q(
        delay_matrix_N_1_next[28]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_2__0_ ( .D(n991), .CP(CLK), .Q(
        delay_matrix_N_1[28]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_2__1_ ( .D(n1068), .CP(CLK), .Q(
        delay_matrix_N_1_next[29]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_2__1_ ( .D(n990), .CP(CLK), .Q(
        delay_matrix_N_1[29]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_2__2_ ( .D(n1067), .CP(CLK), .Q(
        delay_matrix_N_1_next[30]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_2__2_ ( .D(n989), .CP(CLK), .Q(
        delay_matrix_N_1[30]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_2__3_ ( .D(n1066), .CP(CLK), .Q(
        delay_matrix_N_1_next[31]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_2__3_ ( .D(n988), .CP(CLK), .Q(
        delay_matrix_N_1[31]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_2__4_ ( .D(n1065), .CP(CLK), .Q(
        delay_matrix_N_1_next[32]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_2__4_ ( .D(n987), .CP(CLK), .Q(
        delay_matrix_N_1[32]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_2__5_ ( .D(n1064), .CP(CLK), .Q(
        delay_matrix_N_1_next[33]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_2__5_ ( .D(n986), .CP(CLK), .Q(
        delay_matrix_N_1[33]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_2__6_ ( .D(n1063), .CP(CLK), .Q(
        delay_matrix_N_1_next[34]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_2__6_ ( .D(n985), .CP(CLK), .Q(
        delay_matrix_N_1[34]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_2__7_ ( .D(n1062), .CP(CLK), .Q(
        delay_matrix_N_1_next[35]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_2__7_ ( .D(n984), .CP(CLK), .Q(
        delay_matrix_N_1[35]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_2__8_ ( .D(n1061), .CP(CLK), .Q(
        delay_matrix_N_1_next[36]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_2__8_ ( .D(n983), .CP(CLK), .Q(
        delay_matrix_N_1[36]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_2__9_ ( .D(n1060), .CP(CLK), .Q(
        delay_matrix_N_1_next[37]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_2__9_ ( .D(n982), .CP(CLK), .Q(
        delay_matrix_N_1[37]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_2__10_ ( .D(n1059), .CP(CLK), 
        .Q(delay_matrix_N_1_next[38]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_2__10_ ( .D(n981), .CP(CLK), .Q(
        delay_matrix_N_1[38]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_2__11_ ( .D(n1058), .CP(CLK), 
        .Q(delay_matrix_N_1_next[39]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_2__11_ ( .D(n980), .CP(CLK), .Q(
        delay_matrix_N_1[39]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_2__12_ ( .D(n1057), .CP(CLK), 
        .Q(delay_matrix_N_1_next[40]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_2__12_ ( .D(n979), .CP(CLK), .Q(
        delay_matrix_N_1[40]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_2__13_ ( .D(n1056), .CP(CLK), 
        .Q(delay_matrix_N_1_next[41]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_2__13_ ( .D(n978), .CP(CLK), .Q(
        delay_matrix_N_1[41]) );
  DFQD1BWP30P140LVT obj_id_next_reg_2__0_ ( .D(n1053), .CP(CLK), .Q(
        obj_id_next[4]) );
  DFQD1BWP30P140LVT obj_id_reg_2__0_ ( .D(n959), .CP(CLK), .Q(obj_id[4]) );
  DFQD1BWP30P140LVT obj_id_next_reg_2__1_ ( .D(n1052), .CP(CLK), .Q(
        obj_id_next[5]) );
  DFQD1BWP30P140LVT obj_id_reg_2__1_ ( .D(n958), .CP(CLK), .Q(obj_id[5]) );
  DFQD1BWP30P140LVT obj_id_next_reg_0__0_ ( .D(n1051), .CP(CLK), .Q(
        obj_id_next[0]) );
  DFQD1BWP30P140LVT obj_id_reg_0__0_ ( .D(n963), .CP(CLK), .Q(obj_id[0]) );
  DFQD1BWP30P140LVT obj_id_next_reg_0__1_ ( .D(n1050), .CP(CLK), .Q(
        obj_id_next[1]) );
  DFQD1BWP30P140LVT obj_id_reg_0__1_ ( .D(n962), .CP(CLK), .Q(obj_id[1]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_0__0_ ( .D(n1047), .CP(CLK), .Q(
        delay_matrix_N_1_next[0]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_0__0_ ( .D(n1019), .CP(CLK), .Q(
        delay_matrix_N_1[0]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_0__1_ ( .D(n1046), .CP(CLK), .Q(
        delay_matrix_N_1_next[1]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_0__1_ ( .D(n1018), .CP(CLK), .Q(
        delay_matrix_N_1[1]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_0__2_ ( .D(n1045), .CP(CLK), .Q(
        delay_matrix_N_1_next[2]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_0__2_ ( .D(n1017), .CP(CLK), .Q(
        delay_matrix_N_1[2]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_0__3_ ( .D(n1044), .CP(CLK), .Q(
        delay_matrix_N_1_next[3]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_0__3_ ( .D(n1016), .CP(CLK), .Q(
        delay_matrix_N_1[3]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_0__4_ ( .D(n1043), .CP(CLK), .Q(
        delay_matrix_N_1_next[4]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_0__4_ ( .D(n1015), .CP(CLK), .Q(
        delay_matrix_N_1[4]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_0__5_ ( .D(n1042), .CP(CLK), .Q(
        delay_matrix_N_1_next[5]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_0__5_ ( .D(n1014), .CP(CLK), .Q(
        delay_matrix_N_1[5]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_0__6_ ( .D(n1041), .CP(CLK), .Q(
        delay_matrix_N_1_next[6]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_0__6_ ( .D(n1013), .CP(CLK), .Q(
        delay_matrix_N_1[6]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_0__7_ ( .D(n1040), .CP(CLK), .Q(
        delay_matrix_N_1_next[7]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_0__7_ ( .D(n1012), .CP(CLK), .Q(
        delay_matrix_N_1[7]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_0__8_ ( .D(n1039), .CP(CLK), .Q(
        delay_matrix_N_1_next[8]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_0__8_ ( .D(n1011), .CP(CLK), .Q(
        delay_matrix_N_1[8]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_0__9_ ( .D(n1038), .CP(CLK), .Q(
        delay_matrix_N_1_next[9]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_0__9_ ( .D(n1010), .CP(CLK), .Q(
        delay_matrix_N_1[9]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_0__10_ ( .D(n1037), .CP(CLK), 
        .Q(delay_matrix_N_1_next[10]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_0__10_ ( .D(n1009), .CP(CLK), .Q(
        delay_matrix_N_1[10]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_0__11_ ( .D(n1036), .CP(CLK), 
        .Q(delay_matrix_N_1_next[11]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_0__11_ ( .D(n1008), .CP(CLK), .Q(
        delay_matrix_N_1[11]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_0__12_ ( .D(n1035), .CP(CLK), 
        .Q(delay_matrix_N_1_next[12]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_0__12_ ( .D(n1007), .CP(CLK), .Q(
        delay_matrix_N_1[12]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_0__13_ ( .D(n1034), .CP(CLK), 
        .Q(delay_matrix_N_1_next[13]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_0__13_ ( .D(n1006), .CP(CLK), .Q(
        delay_matrix_N_1[13]) );
  DFQD1BWP30P140LVT obj_id_next_reg_1__0_ ( .D(n1049), .CP(CLK), .Q(
        obj_id_next[2]) );
  DFQD1BWP30P140LVT obj_id_reg_1__0_ ( .D(n961), .CP(CLK), .Q(obj_id[2]) );
  DFQD1BWP30P140LVT obj_id_next_reg_1__1_ ( .D(n1048), .CP(CLK), .Q(
        obj_id_next[3]) );
  DFQD1BWP30P140LVT obj_id_reg_1__1_ ( .D(n960), .CP(CLK), .Q(obj_id[3]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_1__0_ ( .D(n1033), .CP(CLK), .Q(
        delay_matrix_N_1_next[14]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_1__0_ ( .D(n1005), .CP(CLK), .Q(
        delay_matrix_N_1[14]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_1__1_ ( .D(n1032), .CP(CLK), .Q(
        delay_matrix_N_1_next[15]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_1__1_ ( .D(n1004), .CP(CLK), .Q(
        delay_matrix_N_1[15]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_1__2_ ( .D(n1031), .CP(CLK), .Q(
        delay_matrix_N_1_next[16]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_1__2_ ( .D(n1003), .CP(CLK), .Q(
        delay_matrix_N_1[16]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_1__3_ ( .D(n1030), .CP(CLK), .Q(
        delay_matrix_N_1_next[17]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_1__3_ ( .D(n1002), .CP(CLK), .Q(
        delay_matrix_N_1[17]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_1__4_ ( .D(n1029), .CP(CLK), .Q(
        delay_matrix_N_1_next[18]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_1__4_ ( .D(n1001), .CP(CLK), .Q(
        delay_matrix_N_1[18]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_1__5_ ( .D(n1028), .CP(CLK), .Q(
        delay_matrix_N_1_next[19]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_1__5_ ( .D(n1000), .CP(CLK), .Q(
        delay_matrix_N_1[19]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_1__6_ ( .D(n1027), .CP(CLK), .Q(
        delay_matrix_N_1_next[20]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_1__6_ ( .D(n999), .CP(CLK), .Q(
        delay_matrix_N_1[20]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_1__7_ ( .D(n1026), .CP(CLK), .Q(
        delay_matrix_N_1_next[21]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_1__7_ ( .D(n998), .CP(CLK), .Q(
        delay_matrix_N_1[21]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_1__8_ ( .D(n1025), .CP(CLK), .Q(
        delay_matrix_N_1_next[22]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_1__8_ ( .D(n997), .CP(CLK), .Q(
        delay_matrix_N_1[22]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_1__9_ ( .D(n1024), .CP(CLK), .Q(
        delay_matrix_N_1_next[23]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_1__9_ ( .D(n996), .CP(CLK), .Q(
        delay_matrix_N_1[23]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_1__10_ ( .D(n1023), .CP(CLK), 
        .Q(delay_matrix_N_1_next[24]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_1__10_ ( .D(n995), .CP(CLK), .Q(
        delay_matrix_N_1[24]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_1__11_ ( .D(n1022), .CP(CLK), 
        .Q(delay_matrix_N_1_next[25]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_1__11_ ( .D(n994), .CP(CLK), .Q(
        delay_matrix_N_1[25]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_1__12_ ( .D(n1021), .CP(CLK), 
        .Q(delay_matrix_N_1_next[26]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_1__12_ ( .D(n993), .CP(CLK), .Q(
        delay_matrix_N_1[26]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_reg_1__13_ ( .D(n1020), .CP(CLK), 
        .Q(delay_matrix_N_1_next[27]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_reg_1__13_ ( .D(n992), .CP(CLK), .Q(
        delay_matrix_N_1[27]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_31_ ( .D(n924), .CP(CLK), .Q(
        copy_ptr_next[31]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_30_ ( .D(n925), .CP(CLK), .Q(
        copy_ptr_next[30]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_29_ ( .D(n926), .CP(CLK), .Q(
        copy_ptr_next[29]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_28_ ( .D(n927), .CP(CLK), .Q(
        copy_ptr_next[28]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_27_ ( .D(n928), .CP(CLK), .Q(
        copy_ptr_next[27]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_26_ ( .D(n929), .CP(CLK), .Q(
        copy_ptr_next[26]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_25_ ( .D(n930), .CP(CLK), .Q(
        copy_ptr_next[25]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_24_ ( .D(n931), .CP(CLK), .Q(
        copy_ptr_next[24]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_23_ ( .D(n932), .CP(CLK), .Q(
        copy_ptr_next[23]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_22_ ( .D(n933), .CP(CLK), .Q(
        copy_ptr_next[22]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_21_ ( .D(n934), .CP(CLK), .Q(
        copy_ptr_next[21]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_20_ ( .D(n935), .CP(CLK), .Q(
        copy_ptr_next[20]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_19_ ( .D(n936), .CP(CLK), .Q(
        copy_ptr_next[19]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_18_ ( .D(n937), .CP(CLK), .Q(
        copy_ptr_next[18]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_17_ ( .D(n938), .CP(CLK), .Q(
        copy_ptr_next[17]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_16_ ( .D(n939), .CP(CLK), .Q(
        copy_ptr_next[16]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_15_ ( .D(n940), .CP(CLK), .Q(
        copy_ptr_next[15]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_14_ ( .D(n941), .CP(CLK), .Q(
        copy_ptr_next[14]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_13_ ( .D(n942), .CP(CLK), .Q(
        copy_ptr_next[13]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_12_ ( .D(n943), .CP(CLK), .Q(
        copy_ptr_next[12]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_11_ ( .D(n944), .CP(CLK), .Q(
        copy_ptr_next[11]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_10_ ( .D(n945), .CP(CLK), .Q(
        copy_ptr_next[10]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_9_ ( .D(n946), .CP(CLK), .Q(
        copy_ptr_next[9]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_8_ ( .D(n947), .CP(CLK), .Q(
        copy_ptr_next[8]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_7_ ( .D(n948), .CP(CLK), .Q(
        copy_ptr_next[7]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_6_ ( .D(n949), .CP(CLK), .Q(
        copy_ptr_next[6]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_5_ ( .D(n950), .CP(CLK), .Q(
        copy_ptr_next[5]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_4_ ( .D(n951), .CP(CLK), .Q(
        copy_ptr_next[4]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_3_ ( .D(n952), .CP(CLK), .Q(
        copy_ptr_next[3]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_2_ ( .D(n953), .CP(CLK), .Q(
        copy_ptr_next[2]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_3__0_ ( .D(n923), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[42]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_3__0_ ( .D(n825), .CP(CLK), 
        .Q(delay_matrix_N_1_original[42]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_3__1_ ( .D(n922), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[43]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_3__1_ ( .D(n824), .CP(CLK), 
        .Q(delay_matrix_N_1_original[43]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_3__2_ ( .D(n921), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[44]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_3__2_ ( .D(n823), .CP(CLK), 
        .Q(delay_matrix_N_1_original[44]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_3__3_ ( .D(n920), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[45]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_3__3_ ( .D(n822), .CP(CLK), 
        .Q(delay_matrix_N_1_original[45]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_3__4_ ( .D(n919), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[46]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_3__4_ ( .D(n821), .CP(CLK), 
        .Q(delay_matrix_N_1_original[46]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_3__5_ ( .D(n918), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[47]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_3__5_ ( .D(n820), .CP(CLK), 
        .Q(delay_matrix_N_1_original[47]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_3__6_ ( .D(n917), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[48]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_3__6_ ( .D(n819), .CP(CLK), 
        .Q(delay_matrix_N_1_original[48]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_3__7_ ( .D(n916), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[49]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_3__7_ ( .D(n818), .CP(CLK), 
        .Q(delay_matrix_N_1_original[49]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_3__8_ ( .D(n915), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[50]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_3__8_ ( .D(n817), .CP(CLK), 
        .Q(delay_matrix_N_1_original[50]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_3__9_ ( .D(n914), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[51]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_3__9_ ( .D(n816), .CP(CLK), 
        .Q(delay_matrix_N_1_original[51]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_3__10_ ( .D(n913), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[52]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_3__10_ ( .D(n815), .CP(CLK), 
        .Q(delay_matrix_N_1_original[52]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_3__11_ ( .D(n912), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[53]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_3__11_ ( .D(n814), .CP(CLK), 
        .Q(delay_matrix_N_1_original[53]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_3__12_ ( .D(n911), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[54]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_3__12_ ( .D(n813), .CP(CLK), 
        .Q(delay_matrix_N_1_original[54]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_3__13_ ( .D(n910), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[55]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_3__13_ ( .D(n812), .CP(CLK), 
        .Q(delay_matrix_N_1_original[55]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_2__0_ ( .D(n909), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[28]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_2__0_ ( .D(n839), .CP(CLK), 
        .Q(delay_matrix_N_1_original[28]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_2__1_ ( .D(n908), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[29]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_2__1_ ( .D(n838), .CP(CLK), 
        .Q(delay_matrix_N_1_original[29]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_2__2_ ( .D(n907), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[30]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_2__2_ ( .D(n837), .CP(CLK), 
        .Q(delay_matrix_N_1_original[30]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_2__3_ ( .D(n906), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[31]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_2__3_ ( .D(n836), .CP(CLK), 
        .Q(delay_matrix_N_1_original[31]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_2__4_ ( .D(n905), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[32]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_2__4_ ( .D(n835), .CP(CLK), 
        .Q(delay_matrix_N_1_original[32]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_2__5_ ( .D(n904), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[33]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_2__5_ ( .D(n834), .CP(CLK), 
        .Q(delay_matrix_N_1_original[33]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_2__6_ ( .D(n903), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[34]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_2__6_ ( .D(n833), .CP(CLK), 
        .Q(delay_matrix_N_1_original[34]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_2__7_ ( .D(n902), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[35]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_2__7_ ( .D(n832), .CP(CLK), 
        .Q(delay_matrix_N_1_original[35]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_2__8_ ( .D(n901), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[36]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_2__8_ ( .D(n831), .CP(CLK), 
        .Q(delay_matrix_N_1_original[36]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_2__9_ ( .D(n900), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[37]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_2__9_ ( .D(n830), .CP(CLK), 
        .Q(delay_matrix_N_1_original[37]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_2__10_ ( .D(n899), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[38]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_2__10_ ( .D(n829), .CP(CLK), 
        .Q(delay_matrix_N_1_original[38]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_2__11_ ( .D(n898), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[39]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_2__11_ ( .D(n828), .CP(CLK), 
        .Q(delay_matrix_N_1_original[39]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_2__12_ ( .D(n897), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[40]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_2__12_ ( .D(n827), .CP(CLK), 
        .Q(delay_matrix_N_1_original[40]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_2__13_ ( .D(n896), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[41]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_2__13_ ( .D(n826), .CP(CLK), 
        .Q(delay_matrix_N_1_original[41]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_0__0_ ( .D(n895), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[0]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_0__0_ ( .D(n867), .CP(CLK), 
        .Q(delay_matrix_N_1_original[0]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_0__1_ ( .D(n894), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[1]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_0__1_ ( .D(n866), .CP(CLK), 
        .Q(delay_matrix_N_1_original[1]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_0__2_ ( .D(n893), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[2]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_0__2_ ( .D(n865), .CP(CLK), 
        .Q(delay_matrix_N_1_original[2]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_0__3_ ( .D(n892), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[3]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_0__3_ ( .D(n864), .CP(CLK), 
        .Q(delay_matrix_N_1_original[3]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_0__4_ ( .D(n891), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[4]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_0__4_ ( .D(n863), .CP(CLK), 
        .Q(delay_matrix_N_1_original[4]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_0__5_ ( .D(n890), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[5]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_0__5_ ( .D(n862), .CP(CLK), 
        .Q(delay_matrix_N_1_original[5]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_0__6_ ( .D(n889), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[6]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_0__6_ ( .D(n861), .CP(CLK), 
        .Q(delay_matrix_N_1_original[6]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_0__7_ ( .D(n888), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[7]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_0__7_ ( .D(n860), .CP(CLK), 
        .Q(delay_matrix_N_1_original[7]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_0__8_ ( .D(n887), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[8]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_0__8_ ( .D(n859), .CP(CLK), 
        .Q(delay_matrix_N_1_original[8]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_0__9_ ( .D(n886), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[9]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_0__9_ ( .D(n858), .CP(CLK), 
        .Q(delay_matrix_N_1_original[9]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_0__10_ ( .D(n885), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[10]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_0__10_ ( .D(n857), .CP(CLK), 
        .Q(delay_matrix_N_1_original[10]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_0__11_ ( .D(n884), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[11]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_0__11_ ( .D(n856), .CP(CLK), 
        .Q(delay_matrix_N_1_original[11]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_0__12_ ( .D(n883), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[12]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_0__12_ ( .D(n855), .CP(CLK), 
        .Q(delay_matrix_N_1_original[12]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_0__13_ ( .D(n882), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[13]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_0__13_ ( .D(n854), .CP(CLK), 
        .Q(delay_matrix_N_1_original[13]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_1__0_ ( .D(n881), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[14]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_1__0_ ( .D(n853), .CP(CLK), 
        .Q(delay_matrix_N_1_original[14]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_1__1_ ( .D(n880), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[15]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_1__1_ ( .D(n852), .CP(CLK), 
        .Q(delay_matrix_N_1_original[15]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_1__2_ ( .D(n879), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[16]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_1__2_ ( .D(n851), .CP(CLK), 
        .Q(delay_matrix_N_1_original[16]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_1__3_ ( .D(n878), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[17]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_1__3_ ( .D(n850), .CP(CLK), 
        .Q(delay_matrix_N_1_original[17]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_1__4_ ( .D(n877), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[18]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_1__4_ ( .D(n849), .CP(CLK), 
        .Q(delay_matrix_N_1_original[18]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_1__5_ ( .D(n876), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[19]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_1__5_ ( .D(n848), .CP(CLK), 
        .Q(delay_matrix_N_1_original[19]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_1__6_ ( .D(n875), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[20]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_1__6_ ( .D(n847), .CP(CLK), 
        .Q(delay_matrix_N_1_original[20]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_1__7_ ( .D(n874), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[21]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_1__7_ ( .D(n846), .CP(CLK), 
        .Q(delay_matrix_N_1_original[21]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_1__8_ ( .D(n873), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[22]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_1__8_ ( .D(n845), .CP(CLK), 
        .Q(delay_matrix_N_1_original[22]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_1__9_ ( .D(n872), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[23]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_1__9_ ( .D(n844), .CP(CLK), 
        .Q(delay_matrix_N_1_original[23]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_1__10_ ( .D(n871), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[24]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_1__10_ ( .D(n843), .CP(CLK), 
        .Q(delay_matrix_N_1_original[24]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_1__11_ ( .D(n870), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[25]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_1__11_ ( .D(n842), .CP(CLK), 
        .Q(delay_matrix_N_1_original[25]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_1__12_ ( .D(n869), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[26]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_1__12_ ( .D(n841), .CP(CLK), 
        .Q(delay_matrix_N_1_original[26]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_next_original_reg_1__13_ ( .D(n868), .CP(
        CLK), .Q(delay_matrix_N_1_next_original[27]) );
  DFQD1BWP30P140LVT delay_matrix_N_1_original_reg_1__13_ ( .D(n840), .CP(CLK), 
        .Q(delay_matrix_N_1_original[27]) );
  DFQD1BWP30P140LVT done2_reg ( .D(n2220), .CP(CLK), .Q(done2) );
  DFQD1BWP30P140LVT done_reg ( .D(N3862), .CP(CLK), .Q(done) );
  DFQD1BWP30P140LVT local_controller_id_int_reg_5_ ( .D(N4214), .CP(CLK), .Q(
        local_controller_id_int[5]) );
  DFQD1BWP30P140LVT local_controller_id_int_reg_4_ ( .D(N4213), .CP(CLK), .Q(
        local_controller_id_int[4]) );
  DFQD1BWP30P140LVT local_controller_id_int_reg_3_ ( .D(N4212), .CP(CLK), .Q(
        local_controller_id_int[3]) );
  DFQD1BWP30P140LVT local_controller_id_int_reg_2_ ( .D(N4211), .CP(CLK), .Q(
        local_controller_id_int[2]) );
  DFQD1BWP30P140LVT local_controller_id_int_reg_1_ ( .D(N4210), .CP(CLK), .Q(
        local_controller_id_int[1]) );
  DFQD1BWP30P140LVT local_controller_id_int_reg_0_ ( .D(N4209), .CP(CLK), .Q(
        local_controller_id_int[0]) );
  DFQD1BWP30P140LVT calc_glob_controller_prefetch_start_int_reg_7_ ( .D(N4208), 
        .CP(CLK), .Q(calc_glob_controller_prefetch_start_int[7]) );
  DFQD1BWP30P140LVT calc_glob_controller_prefetch_start_int_reg_6_ ( .D(N4207), 
        .CP(CLK), .Q(calc_glob_controller_prefetch_start_int[6]) );
  DFQD1BWP30P140LVT calc_glob_controller_prefetch_start_int_reg_5_ ( .D(N4206), 
        .CP(CLK), .Q(calc_glob_controller_prefetch_start_int[5]) );
  DFQD1BWP30P140LVT calc_glob_controller_prefetch_start_int_reg_4_ ( .D(N4205), 
        .CP(CLK), .Q(calc_glob_controller_prefetch_start_int[4]) );
  DFQD1BWP30P140LVT calc_glob_controller_prefetch_start_int_reg_3_ ( .D(N4204), 
        .CP(CLK), .Q(calc_glob_controller_prefetch_start_int[3]) );
  DFQD1BWP30P140LVT calc_glob_controller_prefetch_start_int_reg_2_ ( .D(N4203), 
        .CP(CLK), .Q(calc_glob_controller_prefetch_start_int[2]) );
  DFQD1BWP30P140LVT calc_glob_controller_prefetch_start_int_reg_1_ ( .D(N4202), 
        .CP(CLK), .Q(calc_glob_controller_prefetch_start_int[1]) );
  DFQD1BWP30P140LVT calc_glob_controller_prefetch_start_int_reg_0_ ( .D(N4201), 
        .CP(CLK), .Q(calc_glob_controller_prefetch_start_int[0]) );
  DFQD1BWP30P140LVT tapping_loc_packet_reg_9_ ( .D(N4196), .CP(CLK), .Q(
        tapping_loc_packet[9]) );
  DFQD1BWP30P140LVT tapping_loc_packet_reg_8_ ( .D(N4195), .CP(CLK), .Q(
        tapping_loc_packet[8]) );
  DFQD1BWP30P140LVT tapping_loc_packet_reg_7_ ( .D(N4194), .CP(CLK), .Q(
        tapping_loc_packet[7]) );
  DFQD1BWP30P140LVT tapping_loc_packet_reg_6_ ( .D(N4193), .CP(CLK), .Q(
        tapping_loc_packet[6]) );
  DFQD1BWP30P140LVT tapping_loc_packet_reg_5_ ( .D(N4192), .CP(CLK), .Q(
        tapping_loc_packet[5]) );
  DFQD1BWP30P140LVT tapping_loc_packet_reg_4_ ( .D(N4191), .CP(CLK), .Q(
        tapping_loc_packet[4]) );
  DFQD1BWP30P140LVT tapping_loc_packet_reg_3_ ( .D(N4190), .CP(CLK), .Q(
        tapping_loc_packet[3]) );
  DFQD1BWP30P140LVT tapping_loc_packet_reg_1_ ( .D(n2225), .CP(CLK), .Q(
        tapping_loc_packet[1]) );
  DFQD1BWP30P140LVT tapping_loc_packet_reg_0_ ( .D(n2226), .CP(CLK), .Q(
        tapping_loc_packet[0]) );
  DFQD1BWP30P140LVT calc_global_controller_prefetch_start_reg_7_ ( .D(N4230), 
        .CP(CLK), .Q(calc_global_controller_prefetch_start[7]) );
  DFQD1BWP30P140LVT calc_global_controller_prefetch_start_reg_6_ ( .D(N4229), 
        .CP(CLK), .Q(calc_global_controller_prefetch_start[6]) );
  DFQD1BWP30P140LVT calc_global_controller_prefetch_start_reg_5_ ( .D(N4228), 
        .CP(CLK), .Q(calc_global_controller_prefetch_start[5]) );
  DFQD1BWP30P140LVT calc_global_controller_prefetch_start_reg_4_ ( .D(N4227), 
        .CP(CLK), .Q(calc_global_controller_prefetch_start[4]) );
  DFQD1BWP30P140LVT calc_global_controller_prefetch_start_reg_3_ ( .D(N4226), 
        .CP(CLK), .Q(calc_global_controller_prefetch_start[3]) );
  DFQD1BWP30P140LVT calc_global_controller_prefetch_start_reg_2_ ( .D(N4225), 
        .CP(CLK), .Q(calc_global_controller_prefetch_start[2]) );
  DFQD1BWP30P140LVT calc_global_controller_prefetch_start_reg_1_ ( .D(N4224), 
        .CP(CLK), .Q(calc_global_controller_prefetch_start[1]) );
  DFQD1BWP30P140LVT calc_global_controller_prefetch_start_reg_0_ ( .D(N4223), 
        .CP(CLK), .Q(calc_global_controller_prefetch_start[0]) );
  DFQD1BWP30P140LVT local_controller_id_reg_5_ ( .D(N4236), .CP(CLK), .Q(
        local_controller_id[5]) );
  DFQD1BWP30P140LVT local_controller_id_reg_4_ ( .D(N4235), .CP(CLK), .Q(
        local_controller_id[4]) );
  DFQD1BWP30P140LVT local_controller_id_reg_3_ ( .D(N4234), .CP(CLK), .Q(
        local_controller_id[3]) );
  DFQD1BWP30P140LVT local_controller_id_reg_2_ ( .D(N4233), .CP(CLK), .Q(
        local_controller_id[2]) );
  DFQD1BWP30P140LVT local_controller_id_reg_1_ ( .D(N4232), .CP(CLK), .Q(
        local_controller_id[1]) );
  DFQD1BWP30P140LVT local_controller_id_reg_0_ ( .D(N4231), .CP(CLK), .Q(
        local_controller_id[0]) );
  DFQD1BWP30P140LVT calc_glob_dest_addr_int_reg_3_ ( .D(N4200), .CP(CLK), .Q(
        calc_glob_dest_addr_int[3]) );
  DFQD1BWP30P140LVT calc_glob_dest_addr_reg_3_ ( .D(N4240), .CP(CLK), .Q(
        calc_glob_dest_addr[3]) );
  DFQD1BWP30P140LVT calc_glob_dest_addr_int_reg_2_ ( .D(N4199), .CP(CLK), .Q(
        calc_glob_dest_addr_int[2]) );
  DFQD1BWP30P140LVT calc_glob_dest_addr_reg_2_ ( .D(N4239), .CP(CLK), .Q(
        calc_glob_dest_addr[2]) );
  DFQD1BWP30P140LVT calc_glob_dest_addr_int_reg_1_ ( .D(N4198), .CP(CLK), .Q(
        calc_glob_dest_addr_int[1]) );
  DFQD1BWP30P140LVT calc_glob_dest_addr_reg_1_ ( .D(N4238), .CP(CLK), .Q(
        calc_glob_dest_addr[1]) );
  DFQD1BWP30P140LVT calc_glob_dest_addr_int_reg_0_ ( .D(N4197), .CP(CLK), .Q(
        calc_glob_dest_addr_int[0]) );
  DFQD1BWP30P140LVT calc_glob_dest_addr_reg_0_ ( .D(N4237), .CP(CLK), .Q(
        calc_glob_dest_addr[0]) );
  DFQD1BWP30P140LVT calc_glob_prefetch_stop_int_reg_7_ ( .D(N4222), .CP(CLK), 
        .Q(calc_glob_prefetch_stop_int[7]) );
  DFQD1BWP30P140LVT calc_glob_prefetch_stop_reg_7_ ( .D(N4248), .CP(CLK), .Q(
        calc_glob_prefetch_stop[7]) );
  DFQD1BWP30P140LVT calc_glob_prefetch_stop_int_reg_6_ ( .D(N4221), .CP(CLK), 
        .Q(calc_glob_prefetch_stop_int[6]) );
  DFQD1BWP30P140LVT calc_glob_prefetch_stop_reg_6_ ( .D(N4247), .CP(CLK), .Q(
        calc_glob_prefetch_stop[6]) );
  DFQD1BWP30P140LVT calc_glob_prefetch_stop_int_reg_5_ ( .D(N4220), .CP(CLK), 
        .Q(calc_glob_prefetch_stop_int[5]) );
  DFQD1BWP30P140LVT calc_glob_prefetch_stop_reg_5_ ( .D(N4246), .CP(CLK), .Q(
        calc_glob_prefetch_stop[5]) );
  DFQD1BWP30P140LVT calc_glob_prefetch_stop_int_reg_4_ ( .D(N4219), .CP(CLK), 
        .Q(calc_glob_prefetch_stop_int[4]) );
  DFQD1BWP30P140LVT calc_glob_prefetch_stop_reg_4_ ( .D(N4245), .CP(CLK), .Q(
        calc_glob_prefetch_stop[4]) );
  DFQD1BWP30P140LVT calc_glob_prefetch_stop_int_reg_3_ ( .D(N4218), .CP(CLK), 
        .Q(calc_glob_prefetch_stop_int[3]) );
  DFQD1BWP30P140LVT calc_glob_prefetch_stop_reg_3_ ( .D(N4244), .CP(CLK), .Q(
        calc_glob_prefetch_stop[3]) );
  DFQD1BWP30P140LVT calc_glob_prefetch_stop_int_reg_2_ ( .D(N4217), .CP(CLK), 
        .Q(calc_glob_prefetch_stop_int[2]) );
  DFQD1BWP30P140LVT calc_glob_prefetch_stop_reg_2_ ( .D(N4243), .CP(CLK), .Q(
        calc_glob_prefetch_stop[2]) );
  DFQD1BWP30P140LVT calc_glob_prefetch_stop_int_reg_1_ ( .D(N4216), .CP(CLK), 
        .Q(calc_glob_prefetch_stop_int[1]) );
  DFQD1BWP30P140LVT calc_glob_prefetch_stop_reg_1_ ( .D(N4242), .CP(CLK), .Q(
        calc_glob_prefetch_stop[1]) );
  DFQD1BWP30P140LVT calc_glob_prefetch_stop_int_reg_0_ ( .D(N4215), .CP(CLK), 
        .Q(calc_glob_prefetch_stop_int[0]) );
  DFQD1BWP30P140LVT calc_glob_prefetch_stop_reg_0_ ( .D(N4241), .CP(CLK), .Q(
        calc_glob_prefetch_stop[0]) );
  DFQD1BWP30P140LVT prefetch_bypass_start_addr_reg_12_ ( .D(n784), .CP(CLK), 
        .Q(prefetch_bypass_start_addr[12]) );
  DFQD1BWP30P140LVT prefetch_bypass_start_addr_reg_8_ ( .D(n788), .CP(CLK), 
        .Q(n2232) );
  DFQD1BWP30P140LVT prefetch_bypass_start_addr_reg_5_ ( .D(n791), .CP(CLK), 
        .Q(prefetch_bypass_start_addr[5]) );
  DFQD1BWP30P140LVT prefetch_bypass_start_addr_reg_3_ ( .D(n793), .CP(CLK), 
        .Q(prefetch_bypass_start_addr[3]) );
  DFQD1BWP30P140LVT prefetch_bypass_start_addr_reg_2_ ( .D(n794), .CP(CLK), 
        .Q(prefetch_bypass_start_addr[2]) );
  DFQD1BWP30P140LVT tapping_loc_packet_reg_2_ ( .D(n782), .CP(CLK), .Q(
        tapping_loc_packet[2]) );
  DFQD1BWP30P140LVT prefetch_bypass_start_addr_reg_11_ ( .D(n785), .CP(CLK), 
        .Q(n2231) );
  DFQD1BWP30P140LVT prefetch_bypass_start_addr_reg_1_ ( .D(n795), .CP(CLK), 
        .Q(prefetch_bypass_start_addr[1]) );
  DFQD1BWP30P140LVT prefetch_bypass_cycles_reg_6_ ( .D(n798), .CP(CLK), .Q(
        n2227) );
  DFQD1BWP30P140LVT prefetch_bypass_start_addr_reg_0_ ( .D(n796), .CP(CLK), 
        .Q(n2233) );
  DFQD1BWP30P140LVT prefetch_bypass_cycles_reg_4_ ( .D(n800), .CP(CLK), .Q(
        n2229) );
  DFQD4BWP30P140LVT prefetch_bypass_start_addr_reg_13_ ( .D(n783), .CP(CLK), 
        .Q(prefetch_bypass_start_addr[13]) );
  DFQD4BWP30P140LVT prefetch_bypass_start_addr_reg_6_ ( .D(n790), .CP(CLK), 
        .Q(prefetch_bypass_start_addr[6]) );
  DFQD4BWP30P140LVT table_ptr_reg_0_ ( .D(N3860), .CP(CLK), .Q(table_ptr[0])
         );
  DFQD1BWP30P140LVT prefetch_bypass_cycles_reg_2_ ( .D(n802), .CP(CLK), .Q(
        n2230) );
  DFQD4BWP30P140LVT group_header_reg_1_ ( .D(n811), .CP(CLK), .Q(
        group_header[1]) );
  DFQD1BWP30P140LVT prefetch_bypass_cycles_reg_5_ ( .D(n799), .CP(CLK), .Q(
        n2228) );
  DFQD4BWP30P140LVT group_header_reg_0_ ( .D(n810), .CP(CLK), .Q(
        group_header[0]) );
  DFQD4BWP30P140LVT table_ptr_reg_1_ ( .D(N3861), .CP(CLK), .Q(table_ptr[1])
         );
  DFD1BWP30P140LVT copy_pointer_reg_2_ ( .D(n1145), .CP(CLK), .Q(
        copy_pointer[2]), .QN(n2208) );
  DFQD1BWP30P140LVT ptr_next_reg_1_ ( .D(n1114), .CP(CLK), .Q(ptr_next[1]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_1_ ( .D(n954), .CP(CLK), .Q(
        copy_ptr_next[1]) );
  DFQD2BWP30P140LVT prefetch_bypass_dest_addr_int_reg_3_ ( .D(n805), .CP(CLK), 
        .Q(prefetch_bypass_dest_addr_int[3]) );
  DFQD2BWP30P140LVT prefetch_bypass_dest_addr_int_reg_0_ ( .D(n808), .CP(CLK), 
        .Q(prefetch_bypass_dest_addr_int[0]) );
  DFQD2BWP30P140LVT prefetch_bypass_dest_addr_int_reg_2_ ( .D(n806), .CP(CLK), 
        .Q(prefetch_bypass_dest_addr_int[2]) );
  DFQD2BWP30P140LVT prefetch_bypass_dest_addr_int_reg_1_ ( .D(n807), .CP(CLK), 
        .Q(prefetch_bypass_dest_addr_int[1]) );
  DFQD1BWP30P140LVT copy_pointer_reg_0_ ( .D(n1147), .CP(CLK), .Q(
        copy_pointer[0]) );
  DFQD1BWP30P140LVT copy_pointer_reg_1_ ( .D(n1146), .CP(CLK), .Q(
        copy_pointer[1]) );
  DFQD1BWP30P140LVT copy_ptr_next_reg_0_ ( .D(n955), .CP(CLK), .Q(
        copy_ptr_next[0]) );
  DFQD1BWP30P140LVT ptr_next_reg_0_ ( .D(n1115), .CP(CLK), .Q(ptr_next[0]) );
  DFQD4BWP30P140LVT prefetch_bypass_start_addr_reg_4_ ( .D(n792), .CP(CLK), 
        .Q(prefetch_bypass_start_addr[4]) );
  DFQD4BWP30P140LVT prefetch_bypass_start_addr_reg_7_ ( .D(n789), .CP(CLK), 
        .Q(prefetch_bypass_start_addr[7]) );
  DFQD4BWP30P140LVT prefetch_bypass_start_addr_reg_10_ ( .D(n786), .CP(CLK), 
        .Q(prefetch_bypass_start_addr[10]) );
  DFQD4BWP30P140LVT prefetch_bypass_cycles_reg_7_ ( .D(n797), .CP(CLK), .Q(
        prefetch_bypass_cycles[7]) );
  DFQD4BWP30P140LVT prefetch_bypass_cycles_reg_0_ ( .D(n804), .CP(CLK), .Q(
        prefetch_bypass_cycles[0]) );
  DFQD4BWP30P140LVT prefetch_bypass_cycles_reg_1_ ( .D(n803), .CP(CLK), .Q(
        prefetch_bypass_cycles[1]) );
  DFQD4BWP30P140LVT prefetch_bypass_cycles_reg_3_ ( .D(n801), .CP(CLK), .Q(
        prefetch_bypass_cycles[3]) );
  DFQD4BWP30P140LVT prefetch_bypass_start_addr_reg_9_ ( .D(n787), .CP(CLK), 
        .Q(prefetch_bypass_start_addr[9]) );
  INVD4BWP30P140LVT U3 ( .I(n2176), .ZN(n2124) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(n2174), .A2(n459), .ZN(n460) );
  INVD2BWP30P140LVT U5 ( .I(n517), .ZN(n457) );
  INVD1BWP30P140LVT U6 ( .I(n1241), .ZN(n1751) );
  AOI21OPTREPBD1BWP30P140LVT U7 ( .A1(n1232), .A2(n1231), .B(n1230), .ZN(n1268) );
  NR3OPTPAD2BWP30P140LVT U8 ( .A1(n453), .A2(n452), .A3(n1990), .ZN(n455) );
  CKND2D2BWP30P140LVT U9 ( .A1(n498), .A2(n499), .ZN(n1990) );
  NR2D1BWP30P140LVT U10 ( .A1(n555), .A2(n554), .ZN(n656) );
  INVD1BWP30P140LVT U11 ( .I(n2233), .ZN(n477) );
  INVD2BWP30P140LVT U12 ( .I(delay_matrix_element[5]), .ZN(n1798) );
  NR3D0P7BWP30P140LVT U13 ( .A1(n59), .A2(n58), .A3(n57), .ZN(n2009) );
  NR3D0P7BWP30P140LVT U14 ( .A1(n75), .A2(n74), .A3(n73), .ZN(n2115) );
  NR3D0P7BWP30P140LVT U15 ( .A1(n66), .A2(n65), .A3(n64), .ZN(n2118) );
  INVD1BWP30P140LVT U16 ( .I(n2093), .ZN(n2) );
  INR2D1BWP30P140LVT U17 ( .A1(n79), .B1(n78), .ZN(n239) );
  MOAI22D1BWP30P140LVT U18 ( .A1(n549), .A2(n430), .B1(n56), .B2(n10), .ZN(
        n433) );
  ND2D1BWP30P140LVT U19 ( .A1(n92), .A2(n91), .ZN(n2087) );
  ND2OPTIBD1BWP30P140LVT U20 ( .A1(n149), .A2(n148), .ZN(n2094) );
  ND2D1BWP30P140LVT U21 ( .A1(n104), .A2(n103), .ZN(n2088) );
  ND2OPTIBD1BWP30P140LVT U22 ( .A1(n98), .A2(n97), .ZN(n2156) );
  ND2D1BWP30P140LVT U23 ( .A1(n107), .A2(n106), .ZN(n2092) );
  NR2D1BWP30P140LVT U24 ( .A1(n7), .A2(n715), .ZN(n80) );
  ND2D1BWP30P140LVT U25 ( .A1(n120), .A2(n119), .ZN(n2100) );
  NR2D1BWP30P140LVT U26 ( .A1(n7), .A2(n1987), .ZN(n128) );
  INVD4BWP30P140LVT U27 ( .I(n9), .ZN(n508) );
  INVD4BWP30P140LVT U28 ( .I(n1989), .ZN(n175) );
  INVD3BWP30P140LVT U29 ( .I(n56), .ZN(n9) );
  INVD6BWP30P140LVT U30 ( .I(n373), .ZN(n7) );
  NR2D1BWP30P140LVT U31 ( .A1(table_ptr[1]), .A2(table_ptr[0]), .ZN(n348) );
  INR2D1BWP30P140LVT U32 ( .A1(n2096), .B1(n2098), .ZN(n156) );
  INVD1BWP30P140LVT U33 ( .I(n2104), .ZN(n3) );
  NR2D1BWP30P140LVT U34 ( .A1(n686), .A2(n685), .ZN(n1311) );
  NR2D1BWP30P140LVT U35 ( .A1(n7), .A2(n1977), .ZN(n142) );
  AOI21D1BWP30P140LVT U36 ( .A1(n1553), .A2(n707), .B(n706), .ZN(n1310) );
  NR2D1BWP30P140LVT U37 ( .A1(n9), .A2(n1276), .ZN(n49) );
  INVD1BWP30P140LVT U38 ( .I(n5), .ZN(n1984) );
  INVD2BWP30P140LVT U39 ( .I(n13), .ZN(n6) );
  INVD1BWP30P140LVT U40 ( .I(n1245), .ZN(n1616) );
  OAI21D1BWP30P140LVT U41 ( .A1(n2124), .A2(n1996), .B(n460), .ZN(n783) );
  ND2D1BWP30P140LVT U42 ( .A1(n165), .A2(n185), .ZN(n166) );
  ND2OPTIBD1BWP30P140LVT U43 ( .A1(n1306), .A2(n1821), .ZN(n1073) );
  ND2D1BWP30P140LVT U44 ( .A1(n2100), .A2(n2121), .ZN(n2125) );
  ND2D1BWP30P140LVT U45 ( .A1(n2094), .A2(n2), .ZN(n2160) );
  ND2D1BWP30P140LVT U46 ( .A1(n2100), .A2(n2121), .ZN(n2039) );
  ND2D1BWP30P140LVT U47 ( .A1(n2104), .A2(n2103), .ZN(n2105) );
  ND2D1BWP30P140LVT U48 ( .A1(n239), .A2(n164), .ZN(n165) );
  NR2D1BWP30P140LVT U49 ( .A1(n2100), .A2(n300), .ZN(n250) );
  AOI211OPTREPBD1BWP30P140LVT U50 ( .A1(n8), .A2(delay_matrix_N_1_original[10]), .B(n400), .C(n399), .ZN(n440) );
  ND2D1BWP30P140LVT U51 ( .A1(n8), .A2(delay_matrix_N_1[23]), .ZN(n256) );
  INVD2BWP30P140LVT U52 ( .I(n1994), .ZN(n1) );
  INR2D1BWP30P140LVT U53 ( .A1(n184), .B1(n194), .ZN(n163) );
  AOI21OPTREPBD1BWP30P140LVT U54 ( .A1(n69), .A2(n68), .B(n67), .ZN(n498) );
  ND2D1BWP30P140LVT U55 ( .A1(n2098), .A2(n2097), .ZN(n2045) );
  ND2D1BWP30P140LVT U56 ( .A1(n2098), .A2(n2097), .ZN(n2168) );
  ND2D1BWP30P140LVT U57 ( .A1(n241), .A2(n240), .ZN(n242) );
  XNR2OPTND2BWP30P140LVT U58 ( .A1(n1273), .A2(n1272), .ZN(n1638) );
  INVD1BWP30P140LVT U59 ( .I(n164), .ZN(n2021) );
  ND2D1BWP30P140LVT U60 ( .A1(n268), .A2(n60), .ZN(n181) );
  ND2D1BWP30P140LVT U61 ( .A1(n52), .A2(n51), .ZN(n69) );
  ND2D1BWP30P140LVT U62 ( .A1(n510), .A2(n509), .ZN(n2075) );
  ND2D1BWP30P140LVT U63 ( .A1(n613), .A2(n1748), .ZN(n2188) );
  ND2D1BWP30P140LVT U64 ( .A1(n2088), .A2(n289), .ZN(n293) );
  ND2OPTIBD1BWP30P140LVT U65 ( .A1(n82), .A2(n81), .ZN(n164) );
  ND2D1BWP30P140LVT U66 ( .A1(n636), .A2(n635), .ZN(n2185) );
  INVD1BWP30P140LVT U67 ( .I(n239), .ZN(n241) );
  INVD4BWP30P140LVT U68 ( .I(n1191), .ZN(n4) );
  BUFFD4BWP30P140LVT U69 ( .I(n348), .Z(n1989) );
  NR2D1BWP30P140LVT U70 ( .A1(n168), .A2(n1303), .ZN(n53) );
  NR2D1BWP30P140LVT U71 ( .A1(n168), .A2(n1965), .ZN(n118) );
  NR2D1BWP30P140LVT U72 ( .A1(n168), .A2(n1623), .ZN(n70) );
  AN4D0BWP30P140LVT U73 ( .A1(n482), .A2(n481), .A3(n480), .A4(n479), .Z(n483)
         );
  NR2D1BWP30P140LVT U74 ( .A1(n168), .A2(n1252), .ZN(n61) );
  NR2D1BWP30P140LVT U75 ( .A1(n168), .A2(n1297), .ZN(n43) );
  INVD2BWP30P140LVT U76 ( .I(n561), .ZN(n5) );
  INVD1BWP30P140LVT U77 ( .I(delay_matrix_N_1[45]), .ZN(n1969) );
  INVD1BWP30P140LVT U78 ( .I(delay_matrix_N_1[47]), .ZN(n1961) );
  INVD1BWP30P140LVT U79 ( .I(delay_matrix_N_1[48]), .ZN(n1965) );
  INVD1BWP30P140LVT U80 ( .I(delay_matrix_N_1[49]), .ZN(n1987) );
  INVD1BWP30P140LVT U81 ( .I(delay_matrix_N_1[46]), .ZN(n1977) );
  BUFFD4BWP30P140LVT U82 ( .I(n348), .Z(n8) );
  INVD3BWP30P140LVT U83 ( .I(n1821), .ZN(n1807) );
  NR2OPTPAD2BWP30P140LVT U84 ( .A1(n205), .A2(n1280), .ZN(n561) );
  BUFFD4BWP30P140LVT U85 ( .I(n2230), .Z(prefetch_bypass_cycles[2]) );
  AOI21OPTREPBD1BWP30P140LVT U86 ( .A1(n443), .A2(n442), .B(n441), .ZN(n444)
         );
  OAI211D1BWP30P140LVT U87 ( .A1(n440), .A2(scenario_len[10]), .B(n439), .C(
        n438), .ZN(n441) );
  OR2D1BWP30P140LVT U88 ( .A1(delay_matrix_N_1_original[27]), .A2(
        delay_matrix_N_1_original[26]), .Z(n10) );
  INR2D2BWP30P140LVT U89 ( .A1(table_ptr[0]), .B1(table_ptr[1]), .ZN(n56) );
  INR2D2BWP30P140LVT U90 ( .A1(n86), .B1(n85), .ZN(n499) );
  OAI21D2BWP30P140LVT U91 ( .A1(n1268), .A2(n1267), .B(n1266), .ZN(n1273) );
  OAI211D2BWP30P140LVT U92 ( .A1(n520), .A2(n519), .B(n518), .C(n517), .ZN(
        n530) );
  ND2D3BWP30P140LVT U93 ( .A1(n315), .A2(n1989), .ZN(n517) );
  ND3D1BWP30P140LVT U94 ( .A1(n272), .A2(n325), .A3(n326), .ZN(n287) );
  AOI21D2BWP30P140LVT U95 ( .A1(n2143), .A2(n2141), .B(n2089), .ZN(n2136) );
  OAI21D2BWP30P140LVT U96 ( .A1(n2136), .A2(n2132), .B(n2133), .ZN(n2163) );
  ND4D3BWP30P140LVT U97 ( .A1(n1), .A2(n499), .A3(n498), .A4(n501), .ZN(n2054)
         );
  ND2D1BWP30P140LVT U98 ( .A1(n265), .A2(n264), .ZN(n280) );
  ND2D1BWP30P140LVT U99 ( .A1(n274), .A2(n273), .ZN(n335) );
  ND2D1BWP30P140LVT U100 ( .A1(n270), .A2(n269), .ZN(n339) );
  NR2D1BWP30P140LVT U101 ( .A1(n262), .A2(n263), .ZN(n340) );
  INVD1BWP30P140LVT U102 ( .I(n270), .ZN(n268) );
  OAI21D1BWP30P140LVT U103 ( .A1(n153), .A2(n152), .B(n151), .ZN(n11) );
  INVD1BWP30P140LVT U104 ( .I(n184), .ZN(n195) );
  NR2D1BWP30P140LVT U105 ( .A1(n656), .A2(n659), .ZN(n662) );
  ND2D1BWP30P140LVT U106 ( .A1(copy_ptr_next[16]), .A2(copy_ptr_next[17]), 
        .ZN(n1877) );
  ND2D1BWP30P140LVT U107 ( .A1(ptr_next[16]), .A2(ptr_next[17]), .ZN(n1693) );
  ND2D1BWP30P140LVT U108 ( .A1(pointer[16]), .A2(pointer[17]), .ZN(n1430) );
  ND2D1BWP30P140LVT U109 ( .A1(n268), .A2(n267), .ZN(n276) );
  NR2D1BWP30P140LVT U110 ( .A1(n304), .A2(n250), .ZN(n307) );
  ND2D1BWP30P140LVT U111 ( .A1(n258), .A2(n328), .ZN(n331) );
  ND2OPTIBD1BWP30P140LVT U112 ( .A1(n239), .A2(n238), .ZN(n332) );
  ND2D1BWP30P140LVT U113 ( .A1(n440), .A2(scenario_len[10]), .ZN(n442) );
  ND2D1BWP30P140LVT U114 ( .A1(n72), .A2(n71), .ZN(n327) );
  ND2OPTIBD1BWP30P140LVT U115 ( .A1(n63), .A2(n62), .ZN(n278) );
  ND2OPTIBD1BWP30P140LVT U116 ( .A1(n47), .A2(n46), .ZN(n262) );
  ND2OPTIBD1BWP30P140LVT U117 ( .A1(n55), .A2(n54), .ZN(n270) );
  ND2OPTIBD1BWP30P140LVT U118 ( .A1(n173), .A2(n172), .ZN(n274) );
  INVD1BWP30P140LVT U119 ( .I(n2009), .ZN(n60) );
  ND2D1BWP30P140LVT U120 ( .A1(n707), .A2(n688), .ZN(n690) );
  NR2D1BWP30P140LVT U121 ( .A1(n1309), .A2(n1311), .ZN(n688) );
  ND2OPTIBD1BWP30P140LVT U122 ( .A1(n516), .A2(n518), .ZN(n524) );
  INVD1BWP30P140LVT U123 ( .I(n452), .ZN(n198) );
  ND2D1BWP30P140LVT U124 ( .A1(n586), .A2(n585), .ZN(n590) );
  ND2D1BWP30P140LVT U125 ( .A1(n232), .A2(n1255), .ZN(n716) );
  ND2D1BWP30P140LVT U126 ( .A1(copy_ptr_next[6]), .A2(copy_ptr_next[7]), .ZN(
        n230) );
  ND2D1BWP30P140LVT U127 ( .A1(copy_ptr_next[8]), .A2(copy_ptr_next[9]), .ZN(
        n717) );
  ND2D1BWP30P140LVT U128 ( .A1(copy_ptr_next[18]), .A2(copy_ptr_next[19]), 
        .ZN(n223) );
  ND2D1BWP30P140LVT U129 ( .A1(copy_ptr_next[20]), .A2(copy_ptr_next[21]), 
        .ZN(n1865) );
  ND2D1BWP30P140LVT U130 ( .A1(n604), .A2(n603), .ZN(n608) );
  ND2D1BWP30P140LVT U131 ( .A1(n606), .A2(n605), .ZN(n607) );
  ND2D1BWP30P140LVT U132 ( .A1(n470), .A2(n1470), .ZN(n1701) );
  ND2D1BWP30P140LVT U133 ( .A1(ptr_next[6]), .A2(ptr_next[7]), .ZN(n468) );
  ND2D1BWP30P140LVT U134 ( .A1(ptr_next[8]), .A2(ptr_next[9]), .ZN(n1714) );
  ND2D1BWP30P140LVT U135 ( .A1(ptr_next[18]), .A2(ptr_next[19]), .ZN(n461) );
  ND2D1BWP30P140LVT U136 ( .A1(ptr_next[20]), .A2(ptr_next[21]), .ZN(n1687) );
  INVD1BWP30P140LVT U137 ( .I(n661), .ZN(n640) );
  INVD1BWP30P140LVT U138 ( .I(n2172), .ZN(n700) );
  ND2OPTIBD1BWP30P140LVT U139 ( .A1(n1490), .A2(n1489), .ZN(n1508) );
  ND2D1BWP30P140LVT U140 ( .A1(copy_pointer[6]), .A2(copy_pointer[7]), .ZN(
        n1488) );
  ND2D1BWP30P140LVT U141 ( .A1(copy_pointer[8]), .A2(copy_pointer[9]), .ZN(
        n1524) );
  ND2D1BWP30P140LVT U142 ( .A1(copy_pointer[20]), .A2(copy_pointer[21]), .ZN(
        n1530) );
  ND2D1BWP30P140LVT U143 ( .A1(n216), .A2(n1217), .ZN(n1347) );
  ND2D1BWP30P140LVT U144 ( .A1(pointer[6]), .A2(pointer[7]), .ZN(n214) );
  ND2D1BWP30P140LVT U145 ( .A1(pointer[8]), .A2(pointer[9]), .ZN(n1362) );
  ND2D1BWP30P140LVT U146 ( .A1(pointer[12]), .A2(pointer[13]), .ZN(n1349) );
  ND2D1BWP30P140LVT U147 ( .A1(pointer[18]), .A2(pointer[19]), .ZN(n207) );
  ND2D1BWP30P140LVT U148 ( .A1(pointer[20]), .A2(pointer[21]), .ZN(n1426) );
  ND2D1BWP30P140LVT U149 ( .A1(n276), .A2(n339), .ZN(n271) );
  ND2D1BWP30P140LVT U150 ( .A1(n279), .A2(n278), .ZN(n282) );
  ND2D1BWP30P140LVT U151 ( .A1(n249), .A2(n248), .ZN(n317) );
  NR2D1BWP30P140LVT U152 ( .A1(n292), .A2(n247), .ZN(n248) );
  OA21D1BWP30P140LVT U153 ( .A1(n293), .A2(n292), .B(n291), .Z(n318) );
  ND2D1BWP30P140LVT U154 ( .A1(n307), .A2(n252), .ZN(n316) );
  NR2D1BWP30P140LVT U155 ( .A1(n299), .A2(n251), .ZN(n252) );
  ND2D1BWP30P140LVT U156 ( .A1(n401), .A2(n442), .ZN(n446) );
  ND2D1BWP30P140LVT U157 ( .A1(n409), .A2(n408), .ZN(n418) );
  ND2D1BWP30P140LVT U158 ( .A1(n241), .A2(n2021), .ZN(n185) );
  OAI21D1BWP30P140LVT U159 ( .A1(n153), .A2(n152), .B(n151), .ZN(n196) );
  ND2D1BWP30P140LVT U160 ( .A1(n1231), .A2(n756), .ZN(n764) );
  NR2D1BWP30P140LVT U161 ( .A1(ptr_next[31]), .A2(ptr_next[26]), .ZN(n537) );
  ND2D1BWP30P140LVT U162 ( .A1(n331), .A2(n330), .ZN(n334) );
  ND2OPTIBD1BWP30P140LVT U163 ( .A1(n332), .A2(n242), .ZN(n321) );
  INVD1BWP30P140LVT U164 ( .I(n629), .ZN(n1204) );
  NR2D1BWP30P140LVT U165 ( .A1(n760), .A2(n759), .ZN(n766) );
  INVD1BWP30P140LVT U166 ( .I(n767), .ZN(n757) );
  ND2D1BWP30P140LVT U167 ( .A1(n760), .A2(n759), .ZN(n765) );
  XOR3UD1BWP30P140LVT U168 ( .A1(hardware_latency2[13]), .A2(
        hardware_latency1[13]), .A3(n2203), .Z(n771) );
  ND2D1BWP30P140LVT U169 ( .A1(n181), .A2(n190), .ZN(n68) );
  ND2D1BWP30P140LVT U170 ( .A1(n95), .A2(n94), .ZN(n2085) );
  ND2D1BWP30P140LVT U171 ( .A1(n144), .A2(n143), .ZN(n2093) );
  ND2D1BWP30P140LVT U172 ( .A1(n136), .A2(n135), .ZN(n2096) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n574), .A2(copy_pointer[0]), .Z(n575) );
  NR2D1BWP30P140LVT U174 ( .A1(n559), .A2(copy_pointer[0]), .ZN(n487) );
  ND2D1BWP30P140LVT U175 ( .A1(n1861), .A2(n225), .ZN(n1851) );
  ND2D1BWP30P140LVT U176 ( .A1(copy_ptr_next[22]), .A2(copy_ptr_next[23]), 
        .ZN(n224) );
  NR2D1BWP30P140LVT U177 ( .A1(n233), .A2(n716), .ZN(n742) );
  ND2D1BWP30P140LVT U178 ( .A1(n725), .A2(n229), .ZN(n233) );
  ND2D1BWP30P140LVT U179 ( .A1(copy_ptr_next[14]), .A2(copy_ptr_next[15]), 
        .ZN(n228) );
  AOI21D1BWP30P140LVT U180 ( .A1(n619), .A2(n700), .B(n1245), .ZN(n633) );
  INVD1BWP30P140LVT U181 ( .I(n636), .ZN(n619) );
  INR2D1BWP30P140LVT U182 ( .A1(n699), .B1(pointer[1]), .ZN(n636) );
  ND2D1BWP30P140LVT U183 ( .A1(n699), .A2(n612), .ZN(n1584) );
  ND2D1BWP30P140LVT U184 ( .A1(n1685), .A2(n463), .ZN(n1682) );
  ND2D1BWP30P140LVT U185 ( .A1(ptr_next[22]), .A2(ptr_next[23]), .ZN(n462) );
  NR2D1BWP30P140LVT U186 ( .A1(n471), .A2(n1701), .ZN(n1681) );
  ND2D1BWP30P140LVT U187 ( .A1(n1710), .A2(n467), .ZN(n471) );
  ND2D1BWP30P140LVT U188 ( .A1(ptr_next[14]), .A2(ptr_next[15]), .ZN(n466) );
  AN3D1BWP30P140LVT U189 ( .A1(n629), .A2(ptr_next[0]), .A3(ptr_next[1]), .Z(
        n628) );
  ND2D1BWP30P140LVT U190 ( .A1(n1496), .A2(n1483), .ZN(n1520) );
  NR2D1BWP30P140LVT U191 ( .A1(n1491), .A2(n1508), .ZN(n1495) );
  ND2D1BWP30P140LVT U192 ( .A1(n1509), .A2(n1487), .ZN(n1491) );
  INVD1BWP30P140LVT U193 ( .I(pointer[0]), .ZN(n634) );
  ND2D1BWP30P140LVT U194 ( .A1(pointer[0]), .A2(pointer[1]), .ZN(n1187) );
  ND2D1BWP30P140LVT U195 ( .A1(n1422), .A2(n209), .ZN(n1444) );
  NR2D1BWP30P140LVT U196 ( .A1(n217), .A2(n1347), .ZN(n1343) );
  ND2D1BWP30P140LVT U197 ( .A1(n1348), .A2(n213), .ZN(n217) );
  ND2D1BWP30P140LVT U198 ( .A1(pointer[14]), .A2(pointer[15]), .ZN(n212) );
  ND2D1BWP30P140LVT U199 ( .A1(n524), .A2(n523), .ZN(n528) );
  INR2D1BWP30P140LVT U200 ( .A1(table_parse), .B1(n1280), .ZN(n2000) );
  NR2D1BWP30P140LVT U201 ( .A1(n201), .A2(n1991), .ZN(n2001) );
  OAI21D1BWP30P140LVT U202 ( .A1(n2147), .A2(n2150), .B(n2148), .ZN(n2143) );
  AOI21D1BWP30P140LVT U203 ( .A1(n2128), .A2(n2126), .B(n2101), .ZN(n2108) );
  OAI21D1BWP30P140LVT U204 ( .A1(n2171), .A2(n2167), .B(n2168), .ZN(n2128) );
  ND2OPTIBD6BWP30P140LVT U205 ( .A1(n517), .A2(n458), .ZN(n2174) );
  INR2D2BWP30P140LVT U206 ( .A1(n516), .B1(n515), .ZN(n458) );
  INR2D1BWP30P140LVT U207 ( .A1(n505), .B1(n504), .ZN(n2069) );
  OAI21D1BWP30P140LVT U208 ( .A1(n2034), .A2(n2031), .B(n2032), .ZN(n2038) );
  AOI21D1BWP30P140LVT U209 ( .A1(n2038), .A2(n2037), .B(n2095), .ZN(n2047) );
  ND2D1BWP30P140LVT U210 ( .A1(n89), .A2(n88), .ZN(n2084) );
  ND2OPTIBD2BWP30P140LVT U211 ( .A1(n1), .A2(n513), .ZN(n2023) );
  NR2D1BWP30P140LVT U212 ( .A1(n9), .A2(n1415), .ZN(n74) );
  NR2D1BWP30P140LVT U213 ( .A1(n9), .A2(n1237), .ZN(n65) );
  NR2D1BWP30P140LVT U214 ( .A1(n9), .A2(n1222), .ZN(n58) );
  NR2D1BWP30P140LVT U215 ( .A1(done2), .A2(done), .ZN(n491) );
  ND2OPTIBD1BWP30P140LVT U216 ( .A1(n1197), .A2(n592), .ZN(n1392) );
  ND2OPTIBD1BWP30P140LVT U217 ( .A1(n565), .A2(n4), .ZN(n2196) );
  ND2OPTIBD1BWP30P140LVT U218 ( .A1(n1197), .A2(n596), .ZN(n1404) );
  NR2D1BWP30P140LVT U219 ( .A1(copy_ptr_next[1]), .A2(copy_ptr_next[0]), .ZN(
        n596) );
  ND2OPTIBD1BWP30P140LVT U220 ( .A1(n1197), .A2(n594), .ZN(n1398) );
  INVD1BWP30P140LVT U221 ( .I(delay_matrix_element[9]), .ZN(n1282) );
  INVD1BWP30P140LVT U222 ( .I(delay_matrix_element[3]), .ZN(n1678) );
  INVD1BWP30P140LVT U223 ( .I(delay_matrix_element[2]), .ZN(n1810) );
  INVD1BWP30P140LVT U224 ( .I(n716), .ZN(n1260) );
  INVD1BWP30P140LVT U225 ( .I(n742), .ZN(n1890) );
  INVD1BWP30P140LVT U226 ( .I(n2185), .ZN(n1929) );
  INVD1BWP30P140LVT U227 ( .I(n2183), .ZN(n1933) );
  ND2D1BWP30P140LVT U228 ( .A1(n1205), .A2(glob_scen_noc_input_valid), .ZN(
        n1819) );
  NR2D1BWP30P140LVT U229 ( .A1(n1191), .A2(n634), .ZN(n635) );
  ND2D1BWP30P140LVT U230 ( .A1(n630), .A2(glob_scen_noc_input_valid), .ZN(
        n1815) );
  ND2OPTIBD1BWP30P140LVT U231 ( .A1(n636), .A2(n618), .ZN(n2181) );
  INVD1BWP30P140LVT U232 ( .I(n2191), .ZN(n1953) );
  INVD1BWP30P140LVT U233 ( .I(n2188), .ZN(n1957) );
  ND2D1BWP30P140LVT U234 ( .A1(n610), .A2(n699), .ZN(n2191) );
  NR2D1BWP30P140LVT U235 ( .A1(n1191), .A2(n611), .ZN(n610) );
  ND2D1BWP30P140LVT U236 ( .A1(n4), .A2(n1584), .ZN(n613) );
  ND2D1BWP30P140LVT U237 ( .A1(n780), .A2(glob_scen_noc_input_valid), .ZN(
        n1817) );
  INVD1BWP30P140LVT U238 ( .I(n1701), .ZN(n1716) );
  INVD1BWP30P140LVT U239 ( .I(n1681), .ZN(n1727) );
  HA1D1BWP30P140LVT U240 ( .A(ptr_next[29]), .B(n1914), .CO(n1901), .S(n1915)
         );
  HA1D1BWP30P140LVT U241 ( .A(ptr_next[30]), .B(n1901), .CO(n474), .S(n1902)
         );
  INVD1BWP30P140LVT U242 ( .I(n532), .ZN(n1646) );
  XNR2UD1BWP30P140LVT U243 ( .A1(n546), .A2(n550), .ZN(n1970) );
  INVD1BWP30P140LVT U244 ( .I(n1970), .ZN(n1627) );
  ND2D1BWP30P140LVT U245 ( .A1(n556), .A2(n658), .ZN(n557) );
  INVD1BWP30P140LVT U246 ( .I(n1978), .ZN(n1211) );
  XNR2UD1BWP30P140LVT U247 ( .A1(n646), .A2(n645), .ZN(n1966) );
  ND2D1BWP30P140LVT U248 ( .A1(n644), .A2(n657), .ZN(n645) );
  INVD1BWP30P140LVT U249 ( .I(n1966), .ZN(n1215) );
  XNR2UD1BWP30P140LVT U250 ( .A1(n1553), .A2(n666), .ZN(n1974) );
  ND2D1BWP30P140LVT U251 ( .A1(n1552), .A2(n1550), .ZN(n666) );
  INVD1BWP30P140LVT U252 ( .I(n1974), .ZN(n1254) );
  ND2D1BWP30P140LVT U253 ( .A1(n1556), .A2(n1555), .ZN(n1557) );
  INVD1BWP30P140LVT U254 ( .I(n1958), .ZN(n1692) );
  ND2D1BWP30P140LVT U255 ( .A1(n708), .A2(n1308), .ZN(n709) );
  INVD1BWP30P140LVT U256 ( .I(n1962), .ZN(n1637) );
  ND2D1BWP30P140LVT U257 ( .A1(n1313), .A2(n1312), .ZN(n1314) );
  INVD1BWP30P140LVT U258 ( .I(delay_matrix_N_1[50]), .ZN(n715) );
  ND2D1BWP30P140LVT U259 ( .A1(n694), .A2(n1405), .ZN(n695) );
  INVD1BWP30P140LVT U260 ( .I(n1949), .ZN(n1565) );
  ND2D1BWP30P140LVT U261 ( .A1(n1410), .A2(n1409), .ZN(n1411) );
  INVD1BWP30P140LVT U262 ( .I(delay_matrix_N_1[52]), .ZN(n1252) );
  XOR2UD1BWP30P140LVT U263 ( .A1(n1268), .A2(n1234), .Z(n1631) );
  ND2D1BWP30P140LVT U264 ( .A1(n1233), .A2(n1266), .ZN(n1234) );
  NR2D1BWP30P140LVT U265 ( .A1(n701), .A2(n1191), .ZN(n1982) );
  ND2D1BWP30P140LVT U266 ( .A1(n1271), .A2(n1270), .ZN(n1272) );
  ND2OPTIBD1BWP30P140LVT U267 ( .A1(n628), .A2(glob_scen_noc_input_valid), 
        .ZN(n1813) );
  AOI21D1BWP30P140LVT U268 ( .A1(n701), .A2(n700), .B(n1245), .ZN(n1988) );
  INVD1BWP30P140LVT U269 ( .I(n1495), .ZN(n1540) );
  ND2D1BWP30P140LVT U270 ( .A1(n1364), .A2(n1348), .ZN(n1377) );
  INVD1BWP30P140LVT U271 ( .I(n1343), .ZN(n1445) );
  BUFFD3BWP30P140LVT U272 ( .I(n2229), .Z(prefetch_bypass_cycles[4]) );
  BUFFD3BWP30P140LVT U273 ( .I(n2228), .Z(prefetch_bypass_cycles[5]) );
  BUFFD4BWP30P140LVT U274 ( .I(n2227), .Z(prefetch_bypass_cycles[6]) );
  ND2D1BWP30P140LVT U275 ( .A1(n258), .A2(n257), .ZN(n283) );
  NR2D1BWP30P140LVT U276 ( .A1(n2092), .A2(n290), .ZN(n292) );
  ND2D1BWP30P140LVT U277 ( .A1(n507), .A2(delay_matrix_N_1_original[37]), .ZN(
        n428) );
  NR2D1BWP30P140LVT U278 ( .A1(n1267), .A2(n1269), .ZN(n756) );
  NR2D1BWP30P140LVT U279 ( .A1(n2104), .A2(n301), .ZN(n304) );
  ND2D1BWP30P140LVT U280 ( .A1(n2100), .A2(n300), .ZN(n303) );
  NR2D1BWP30P140LVT U281 ( .A1(n2098), .A2(n295), .ZN(n299) );
  ND2D1BWP30P140LVT U282 ( .A1(n294), .A2(n2094), .ZN(n298) );
  XNR2UD1BWP30P140LVT U283 ( .A1(n329), .A2(n283), .ZN(n284) );
  ND2D1BWP30P140LVT U284 ( .A1(n327), .A2(n255), .ZN(n330) );
  ND2D1BWP30P140LVT U285 ( .A1(n170), .A2(delay_matrix_N_1[5]), .ZN(n137) );
  AOI21D1BWP30P140LVT U286 ( .A1(n113), .A2(n112), .B(n111), .ZN(n153) );
  ND2D1BWP30P140LVT U287 ( .A1(n2086), .A2(n2087), .ZN(n112) );
  ND2D1BWP30P140LVT U288 ( .A1(n12), .A2(n2088), .ZN(n117) );
  NR3D0P7BWP30P140LVT U289 ( .A1(n154), .A2(n156), .A3(n150), .ZN(n151) );
  ND2D1BWP30P140LVT U290 ( .A1(n2121), .A2(n2100), .ZN(n162) );
  ND2OPTIBD1BWP30P140LVT U291 ( .A1(n159), .A2(n158), .ZN(n184) );
  ND2D1BWP30P140LVT U292 ( .A1(n2), .A2(n2094), .ZN(n157) );
  ND2D1BWP30P140LVT U293 ( .A1(n190), .A2(n189), .ZN(n191) );
  ND2D1BWP30P140LVT U294 ( .A1(n188), .A2(n187), .ZN(n192) );
  ND2D1BWP30P140LVT U295 ( .A1(n186), .A2(n185), .ZN(n193) );
  ND2D1BWP30P140LVT U296 ( .A1(n25), .A2(n24), .ZN(n264) );
  ND2D1BWP30P140LVT U297 ( .A1(n405), .A2(delay_matrix_N_1[38]), .ZN(n24) );
  ND2D1BWP30P140LVT U298 ( .A1(n27), .A2(n26), .ZN(n267) );
  ND2D1BWP30P140LVT U299 ( .A1(n405), .A2(delay_matrix_N_1[40]), .ZN(n26) );
  ND2D1BWP30P140LVT U300 ( .A1(n310), .A2(n321), .ZN(n311) );
  ND2D1BWP30P140LVT U301 ( .A1(n254), .A2(n253), .ZN(n308) );
  NR2D1BWP30P140LVT U302 ( .A1(n310), .A2(n321), .ZN(n309) );
  ND2D1BWP30P140LVT U303 ( .A1(n421), .A2(n420), .ZN(n450) );
  INVD1BWP30P140LVT U304 ( .I(n165), .ZN(n83) );
  ND2D1BWP30P140LVT U305 ( .A1(n327), .A2(n2115), .ZN(n186) );
  ND2D1BWP30P140LVT U306 ( .A1(n278), .A2(n2118), .ZN(n187) );
  INVD1BWP30P140LVT U307 ( .I(n2006), .ZN(n51) );
  INVD1BWP30P140LVT U308 ( .I(n262), .ZN(n52) );
  NR2D1BWP30P140LVT U309 ( .A1(n278), .A2(n2118), .ZN(n76) );
  ND2D1BWP30P140LVT U310 ( .A1(n262), .A2(n2006), .ZN(n189) );
  ND2D1BWP30P140LVT U311 ( .A1(n270), .A2(n2009), .ZN(n190) );
  NR2D1BWP30P140LVT U312 ( .A1(n141), .A2(n140), .ZN(n155) );
  OAI21D1BWP30P140LVT U313 ( .A1(n1961), .A2(n168), .B(n139), .ZN(n140) );
  ND2D1BWP30P140LVT U314 ( .A1(n138), .A2(n137), .ZN(n141) );
  ND2D1BWP30P140LVT U315 ( .A1(n125), .A2(delay_matrix_N_1[33]), .ZN(n139) );
  NR2D1BWP30P140LVT U316 ( .A1(n7), .A2(n1961), .ZN(n132) );
  AOI21D1BWP30P140LVT U317 ( .A1(n188), .A2(n183), .B(n182), .ZN(n452) );
  INVD1BWP30P140LVT U318 ( .I(n181), .ZN(n182) );
  ND2D1BWP30P140LVT U319 ( .A1(n180), .A2(n179), .ZN(n183) );
  ND2D1BWP30P140LVT U320 ( .A1(n28), .A2(n256), .ZN(n328) );
  INVD1BWP30P140LVT U321 ( .I(n264), .ZN(n279) );
  AOI21D1BWP30P140LVT U322 ( .A1(n405), .A2(delay_matrix_N_1[39]), .B(n23), 
        .ZN(n263) );
  ND2D1BWP30P140LVT U323 ( .A1(n36), .A2(n35), .ZN(n238) );
  ND2D1BWP30P140LVT U324 ( .A1(n8), .A2(delay_matrix_N_1[22]), .ZN(n35) );
  NR2D1BWP30P140LVT U325 ( .A1(n564), .A2(copy_pointer[1]), .ZN(n574) );
  NR2D1BWP30P140LVT U326 ( .A1(copy_ptr_next[31]), .A2(copy_ptr_next[26]), 
        .ZN(n587) );
  IND2D1BWP30P140LVT U327 ( .A1(n564), .B1(copy_pointer[1]), .ZN(n559) );
  INVD1BWP30P140LVT U328 ( .I(delay_matrix_element[2]), .ZN(n641) );
  OAI21D1BWP30P140LVT U329 ( .A1(n553), .A2(n552), .B(n551), .ZN(n661) );
  INVD1BWP30P140LVT U330 ( .I(delay_matrix_element[3]), .ZN(n663) );
  NR2D1BWP30P140LVT U331 ( .A1(n665), .A2(n664), .ZN(n680) );
  NR2D1BWP30P140LVT U332 ( .A1(n680), .A2(n1554), .ZN(n707) );
  INVD1BWP30P140LVT U333 ( .I(delay_matrix_element[9]), .ZN(n748) );
  NR2D1BWP30P140LVT U334 ( .A1(n1406), .A2(n1408), .ZN(n1231) );
  NR2D1BWP30P140LVT U335 ( .A1(n542), .A2(n541), .ZN(n629) );
  ND2D1BWP30P140LVT U336 ( .A1(table_parse), .A2(n491), .ZN(n521) );
  ND3D2BWP30P140LVT U337 ( .A1(n347), .A2(n346), .A3(n345), .ZN(n516) );
  ND2D1BWP30P140LVT U338 ( .A1(n324), .A2(n19), .ZN(n346) );
  OR2D1BWP30P140LVT U339 ( .A1(n497), .A2(n1280), .Z(n501) );
  ND2D1BWP30P140LVT U340 ( .A1(table_parse), .A2(done), .ZN(n497) );
  INVD2BWP30P140LVT U341 ( .I(n549), .ZN(n503) );
  INVD1BWP30P140LVT U342 ( .I(group_header[0]), .ZN(n44) );
  INVD1BWP30P140LVT U343 ( .I(group_header[1]), .ZN(n45) );
  NR2D1BWP30P140LVT U344 ( .A1(n168), .A2(n1977), .ZN(n147) );
  ND2D1BWP30P140LVT U345 ( .A1(n123), .A2(n122), .ZN(n2099) );
  NR2D1BWP30P140LVT U346 ( .A1(n7), .A2(n1965), .ZN(n121) );
  INVD1BWP30P140LVT U347 ( .I(n1990), .ZN(n511) );
  INR2D1BWP30P140LVT U348 ( .A1(n500), .B1(n1991), .ZN(n512) );
  AOI21D1BWP30P140LVT U349 ( .A1(n405), .A2(delay_matrix_N_1[41]), .B(n29), 
        .ZN(n273) );
  INVD1BWP30P140LVT U350 ( .I(n238), .ZN(n240) );
  ND2OPTIBD1BWP30P140LVT U351 ( .A1(copy_ptr_next[1]), .A2(copy_ptr_next[0]), 
        .ZN(n727) );
  NR2D1BWP30P140LVT U352 ( .A1(n231), .A2(n727), .ZN(n1255) );
  ND2D1BWP30P140LVT U353 ( .A1(copy_ptr_next[2]), .A2(copy_ptr_next[3]), .ZN(
        n231) );
  ND2D1BWP30P140LVT U354 ( .A1(copy_ptr_next[4]), .A2(copy_ptr_next[5]), .ZN(
        n1256) );
  ND2D1BWP30P140LVT U355 ( .A1(copy_ptr_next[10]), .A2(copy_ptr_next[11]), 
        .ZN(n227) );
  ND2D1BWP30P140LVT U356 ( .A1(copy_ptr_next[12]), .A2(copy_ptr_next[13]), 
        .ZN(n733) );
  ND2D1BWP30P140LVT U357 ( .A1(n634), .A2(pointer[1]), .ZN(n611) );
  ND2OPTIBD1BWP30P140LVT U358 ( .A1(ptr_next[1]), .A2(ptr_next[0]), .ZN(n1825)
         );
  NR2D1BWP30P140LVT U359 ( .A1(n469), .A2(n1825), .ZN(n1470) );
  ND2D1BWP30P140LVT U360 ( .A1(ptr_next[2]), .A2(ptr_next[3]), .ZN(n469) );
  ND2D1BWP30P140LVT U361 ( .A1(ptr_next[4]), .A2(ptr_next[5]), .ZN(n1474) );
  ND2D1BWP30P140LVT U362 ( .A1(ptr_next[10]), .A2(ptr_next[11]), .ZN(n465) );
  ND2D1BWP30P140LVT U363 ( .A1(ptr_next[12]), .A2(ptr_next[13]), .ZN(n1711) );
  ND2D1BWP30P140LVT U364 ( .A1(n544), .A2(n1793), .ZN(n551) );
  NR2D1BWP30P140LVT U365 ( .A1(n544), .A2(n1793), .ZN(n553) );
  NR2D1BWP30P140LVT U366 ( .A1(n643), .A2(n642), .ZN(n659) );
  ND2D1BWP30P140LVT U367 ( .A1(n643), .A2(n642), .ZN(n657) );
  ND2D1BWP30P140LVT U368 ( .A1(n665), .A2(n664), .ZN(n1550) );
  NR2D1BWP30P140LVT U369 ( .A1(n682), .A2(n681), .ZN(n1554) );
  ND2D1BWP30P140LVT U370 ( .A1(n684), .A2(n683), .ZN(n1308) );
  NR2D1BWP30P140LVT U371 ( .A1(n684), .A2(n683), .ZN(n1309) );
  NR2D1BWP30P140LVT U372 ( .A1(n750), .A2(n749), .ZN(n1408) );
  ND2D1BWP30P140LVT U373 ( .A1(n693), .A2(n692), .ZN(n1405) );
  NR2D1BWP30P140LVT U374 ( .A1(n693), .A2(n692), .ZN(n1406) );
  ND2D1BWP30P140LVT U375 ( .A1(n750), .A2(n749), .ZN(n1409) );
  NR2D1BWP30P140LVT U376 ( .A1(n754), .A2(n753), .ZN(n1269) );
  ND2D1BWP30P140LVT U377 ( .A1(n752), .A2(n751), .ZN(n1266) );
  NR2D1BWP30P140LVT U378 ( .A1(n752), .A2(n751), .ZN(n1267) );
  ND2D1BWP30P140LVT U379 ( .A1(n754), .A2(n753), .ZN(n1270) );
  ND2D1BWP30P140LVT U380 ( .A1(n761), .A2(n765), .ZN(n762) );
  ND2D1BWP30P140LVT U381 ( .A1(n773), .A2(n772), .ZN(n774) );
  ND2D1BWP30P140LVT U382 ( .A1(n771), .A2(n770), .ZN(n772) );
  ND2OPTIBD1BWP30P140LVT U383 ( .A1(copy_pointer[0]), .A2(copy_pointer[1]), 
        .ZN(n1201) );
  NR2D1BWP30P140LVT U384 ( .A1(n1202), .A2(n1201), .ZN(n1489) );
  ND2D1BWP30P140LVT U385 ( .A1(copy_pointer[2]), .A2(copy_pointer[3]), .ZN(
        n1202) );
  ND2D1BWP30P140LVT U386 ( .A1(copy_pointer[4]), .A2(copy_pointer[5]), .ZN(
        n1535) );
  ND2D1BWP30P140LVT U387 ( .A1(copy_pointer[10]), .A2(copy_pointer[11]), .ZN(
        n1485) );
  ND2D1BWP30P140LVT U388 ( .A1(copy_pointer[12]), .A2(copy_pointer[13]), .ZN(
        n1510) );
  ND2D1BWP30P140LVT U389 ( .A1(copy_pointer[16]), .A2(copy_pointer[17]), .ZN(
        n1501) );
  INVD1BWP30P140LVT U390 ( .I(n204), .ZN(n206) );
  INR2D1BWP30P140LVT U391 ( .A1(boot_up), .B1(n203), .ZN(n204) );
  INVD1BWP30P140LVT U392 ( .I(input_valid), .ZN(n203) );
  ND2D1BWP30P140LVT U393 ( .A1(pointer[2]), .A2(pointer[3]), .ZN(n215) );
  ND2D1BWP30P140LVT U394 ( .A1(pointer[4]), .A2(pointer[5]), .ZN(n1339) );
  ND2D1BWP30P140LVT U395 ( .A1(pointer[10]), .A2(pointer[11]), .ZN(n211) );
  INVD1BWP30P140LVT U396 ( .I(glob_scen_noc_input_valid), .ZN(n222) );
  ND2D1BWP30P140LVT U397 ( .A1(n496), .A2(n494), .ZN(n548) );
  OR2D1BWP30P140LVT U398 ( .A1(n512), .A2(n502), .Z(n2055) );
  INVD1BWP30P140LVT U399 ( .I(n501), .ZN(n502) );
  INVD2BWP30P140LVT U400 ( .I(n2054), .ZN(n2068) );
  INVD1BWP30P140LVT U401 ( .I(n2055), .ZN(n2067) );
  NR2D1BWP30P140LVT U402 ( .A1(n9), .A2(n1243), .ZN(n177) );
  OAI21D2BWP30P140LVT U403 ( .A1(n1994), .A2(n1993), .B(n1992), .ZN(n2079) );
  INVD1BWP30P140LVT U404 ( .I(n1991), .ZN(n1992) );
  ND2D1BWP30P140LVT U405 ( .A1(n1260), .A2(n725), .ZN(n738) );
  ND2D1BWP30P140LVT U406 ( .A1(copy_ptr_next[24]), .A2(copy_ptr_next[25]), 
        .ZN(n226) );
  INVD1BWP30P140LVT U407 ( .I(delay_matrix_N_1[27]), .ZN(n1243) );
  INVD1BWP30P140LVT U408 ( .I(delay_matrix_N_1[25]), .ZN(n1276) );
  ND2D1BWP30P140LVT U409 ( .A1(n1819), .A2(n1821), .ZN(n1227) );
  INVD1BWP30P140LVT U410 ( .I(n1205), .ZN(n1228) );
  INVD1BWP30P140LVT U411 ( .I(n2179), .ZN(n1248) );
  ND2D1BWP30P140LVT U412 ( .A1(n1815), .A2(n1821), .ZN(n776) );
  INVD1BWP30P140LVT U413 ( .I(n630), .ZN(n777) );
  ND2D1BWP30P140LVT U414 ( .A1(n1817), .A2(n1821), .ZN(n1223) );
  INVD1BWP30P140LVT U415 ( .I(n780), .ZN(n1224) );
  ND2D1BWP30P140LVT U416 ( .A1(n1716), .A2(n1710), .ZN(n1729) );
  HA1D1BWP30P140LVT U417 ( .A(ptr_next[26]), .B(n17), .CO(n1908), .S(n1679) );
  ND2D1BWP30P140LVT U418 ( .A1(ptr_next[24]), .A2(ptr_next[25]), .ZN(n464) );
  HA1D1BWP30P140LVT U419 ( .A(ptr_next[27]), .B(n1908), .CO(n1911), .S(n1909)
         );
  ND2D1BWP30P140LVT U420 ( .A1(n6), .A2(obj_id_element[0]), .ZN(n1208) );
  ND2D1BWP30P140LVT U421 ( .A1(n6), .A2(obj_id_element[1]), .ZN(n1206) );
  INVD1BWP30P140LVT U422 ( .I(delay_matrix_N_1[51]), .ZN(n1623) );
  INVD1BWP30P140LVT U423 ( .I(delay_matrix_N_1[53]), .ZN(n1297) );
  INVD1BWP30P140LVT U424 ( .I(delay_matrix_N_1[54]), .ZN(n1303) );
  ND2D1BWP30P140LVT U425 ( .A1(n1219), .A2(n6), .ZN(n1229) );
  INVD1BWP30P140LVT U426 ( .I(delay_matrix_N_1[55]), .ZN(n1462) );
  INVD1BWP30P140LVT U427 ( .I(n1982), .ZN(n1461) );
  ND2D1BWP30P140LVT U428 ( .A1(n1241), .A2(n6), .ZN(n1225) );
  ND2D1BWP30P140LVT U429 ( .A1(n1813), .A2(n1760), .ZN(n778) );
  INVD1BWP30P140LVT U430 ( .I(n628), .ZN(n779) );
  INVD1BWP30P140LVT U431 ( .I(n1508), .ZN(n1614) );
  ND2D1BWP30P140LVT U432 ( .A1(n1614), .A2(n1509), .ZN(n1513) );
  ND2D1BWP30P140LVT U433 ( .A1(copy_pointer[24]), .A2(copy_pointer[25]), .ZN(
        n1484) );
  INVD1BWP30P140LVT U434 ( .I(n1347), .ZN(n1364) );
  ND2D1BWP30P140LVT U435 ( .A1(n1381), .A2(n1350), .ZN(n1354) );
  ND2D1BWP30P140LVT U436 ( .A1(pointer[24]), .A2(pointer[25]), .ZN(n210) );
  ND2D1BWP30P140LVT U437 ( .A1(n528), .A2(prefetch_bypass_dest_addr_int[1]), 
        .ZN(n525) );
  ND2D1BWP30P140LVT U438 ( .A1(n528), .A2(prefetch_bypass_dest_addr_int[2]), 
        .ZN(n526) );
  ND2D1BWP30P140LVT U439 ( .A1(n528), .A2(prefetch_bypass_dest_addr_int[0]), 
        .ZN(n527) );
  ND2D1BWP30P140LVT U440 ( .A1(n528), .A2(prefetch_bypass_dest_addr_int[3]), 
        .ZN(n529) );
  ND2D1BWP30P140LVT U441 ( .A1(n2000), .A2(group_header[0]), .ZN(n202) );
  ND2D1BWP30P140LVT U442 ( .A1(n2174), .A2(n2173), .ZN(n2175) );
  ND2D1BWP30P140LVT U443 ( .A1(n2000), .A2(group_header[1]), .ZN(n2003) );
  ND2D1BWP30P140LVT U444 ( .A1(n2174), .A2(n2144), .ZN(n2145) );
  ND2D1BWP30P140LVT U445 ( .A1(n2112), .A2(n2111), .ZN(n797) );
  ND2D1BWP30P140LVT U446 ( .A1(n2174), .A2(n2110), .ZN(n2111) );
  ND2D1BWP30P140LVT U447 ( .A1(n2109), .A2(n2176), .ZN(n2112) );
  ND2D1BWP30P140LVT U448 ( .A1(n2174), .A2(n2082), .ZN(n2083) );
  ND2D1BWP30P140LVT U449 ( .A1(n2174), .A2(n2137), .ZN(n2138) );
  ND2D1BWP30P140LVT U450 ( .A1(n2174), .A2(n2122), .ZN(n2123) );
  ND2D1BWP30P140LVT U451 ( .A1(n2174), .A2(n2164), .ZN(n2165) );
  ND2D1BWP30P140LVT U452 ( .A1(n2174), .A2(n2113), .ZN(n2114) );
  ND2D1BWP30P140LVT U453 ( .A1(n2174), .A2(n2157), .ZN(n2158) );
  ND2D1BWP30P140LVT U454 ( .A1(n2174), .A2(n2152), .ZN(n2153) );
  ND2D1BWP30P140LVT U455 ( .A1(n2174), .A2(n2116), .ZN(n2117) );
  ND2D1BWP30P140LVT U456 ( .A1(n2174), .A2(n2012), .ZN(n2013) );
  ND2D1BWP30P140LVT U457 ( .A1(n2174), .A2(n2129), .ZN(n2130) );
  ND2D1BWP30P140LVT U458 ( .A1(n2174), .A2(n1998), .ZN(n1999) );
  ND2D1BWP30P140LVT U459 ( .A1(n2174), .A2(n2004), .ZN(n2005) );
  ND2D1BWP30P140LVT U460 ( .A1(n2174), .A2(n2017), .ZN(n2018) );
  ND2D1BWP30P140LVT U461 ( .A1(n2174), .A2(n2010), .ZN(n2011) );
  ND2D1BWP30P140LVT U462 ( .A1(n2174), .A2(n2015), .ZN(n2016) );
  ND2D1BWP30P140LVT U463 ( .A1(n2174), .A2(n2019), .ZN(n2020) );
  ND2D1BWP30P140LVT U464 ( .A1(n2174), .A2(n2007), .ZN(n2008) );
  AN3D1BWP30P140LVT U465 ( .A1(n2054), .A2(calc_glob_prefetch_stop_int[0]), 
        .A3(n2055), .Z(N4241) );
  AN3D1BWP30P140LVT U466 ( .A1(n2054), .A2(calc_glob_prefetch_stop_int[1]), 
        .A3(n2055), .Z(N4242) );
  AN3D1BWP30P140LVT U467 ( .A1(n2054), .A2(calc_glob_prefetch_stop_int[2]), 
        .A3(n2055), .Z(N4243) );
  AN3D1BWP30P140LVT U468 ( .A1(n2054), .A2(calc_glob_prefetch_stop_int[3]), 
        .A3(n2055), .Z(N4244) );
  AN3D1BWP30P140LVT U469 ( .A1(n2054), .A2(calc_glob_prefetch_stop_int[4]), 
        .A3(n2055), .Z(N4245) );
  AN3D1BWP30P140LVT U470 ( .A1(n2054), .A2(calc_glob_prefetch_stop_int[5]), 
        .A3(n2055), .Z(N4246) );
  AN3D1BWP30P140LVT U471 ( .A1(n2054), .A2(calc_glob_prefetch_stop_int[6]), 
        .A3(n2055), .Z(N4247) );
  AN3D1BWP30P140LVT U472 ( .A1(n2054), .A2(calc_glob_prefetch_stop_int[7]), 
        .A3(n2055), .Z(N4248) );
  AN3D1BWP30P140LVT U473 ( .A1(n2054), .A2(calc_glob_dest_addr_int[0]), .A3(
        n2055), .Z(N4237) );
  ND2D1BWP30P140LVT U474 ( .A1(n1995), .A2(calc_glob_dest_addr_int[0]), .ZN(
        n514) );
  NR2D1BWP30P140LVT U475 ( .A1(n1991), .A2(n2069), .ZN(n2226) );
  ND2D1BWP30P140LVT U476 ( .A1(n2149), .A2(n2050), .ZN(n2052) );
  ND2D1BWP30P140LVT U477 ( .A1(n2027), .A2(n2026), .ZN(n2022) );
  ND2D1BWP30P140LVT U478 ( .A1(n2088), .A2(n12), .ZN(n2026) );
  ND2D1BWP30P140LVT U479 ( .A1(n2134), .A2(n2032), .ZN(n2033) );
  ND2D1BWP30P140LVT U480 ( .A1(n2037), .A2(n2036), .ZN(n2029) );
  ND2D1BWP30P140LVT U481 ( .A1(n2094), .A2(n2), .ZN(n2036) );
  ND2D1BWP30P140LVT U482 ( .A1(n2169), .A2(n2045), .ZN(n2046) );
  ND2D1BWP30P140LVT U483 ( .A1(n2040), .A2(n2039), .ZN(n2041) );
  NR2D1BWP30P140LVT U484 ( .A1(n2172), .A2(n493), .ZN(n2220) );
  ND2D1BWP30P140LVT U485 ( .A1(n1392), .A2(delay_matrix_N_1_next_original[27]), 
        .ZN(n626) );
  ND2D1BWP30P140LVT U486 ( .A1(n1392), .A2(delay_matrix_N_1_next_original[26]), 
        .ZN(n624) );
  ND2D1BWP30P140LVT U487 ( .A1(n1392), .A2(delay_matrix_N_1_next_original[25]), 
        .ZN(n672) );
  ND2D1BWP30P140LVT U488 ( .A1(n1392), .A2(delay_matrix_N_1_next_original[24]), 
        .ZN(n673) );
  ND2D1BWP30P140LVT U489 ( .A1(n2200), .A2(delay_matrix_N_1_original[23]), 
        .ZN(n577) );
  ND2D1BWP30P140LVT U490 ( .A1(n1762), .A2(delay_matrix_element[8]), .ZN(n675)
         );
  ND2D1BWP30P140LVT U491 ( .A1(n2200), .A2(delay_matrix_N_1_original[21]), 
        .ZN(n1675) );
  ND2D1BWP30P140LVT U492 ( .A1(n2200), .A2(delay_matrix_N_1_original[20]), 
        .ZN(n1671) );
  ND2D1BWP30P140LVT U493 ( .A1(n2200), .A2(delay_matrix_N_1_original[19]), 
        .ZN(n1785) );
  ND2D1BWP30P140LVT U494 ( .A1(n2200), .A2(delay_matrix_N_1_original[18]), 
        .ZN(n1789) );
  ND2D1BWP30P140LVT U495 ( .A1(n2200), .A2(delay_matrix_N_1_original[17]), 
        .ZN(n1654) );
  ND2D1BWP30P140LVT U496 ( .A1(n2200), .A2(delay_matrix_N_1_original[16]), 
        .ZN(n1800) );
  ND2D1BWP30P140LVT U497 ( .A1(n2200), .A2(delay_matrix_N_1_original[15]), 
        .ZN(n1664) );
  ND2D1BWP30P140LVT U498 ( .A1(n1762), .A2(delay_matrix_element[0]), .ZN(n1763) );
  ND2D1BWP30P140LVT U499 ( .A1(n1404), .A2(delay_matrix_N_1_next_original[13]), 
        .ZN(n623) );
  ND2D1BWP30P140LVT U500 ( .A1(n1404), .A2(delay_matrix_N_1_next_original[12]), 
        .ZN(n622) );
  ND2D1BWP30P140LVT U501 ( .A1(n1404), .A2(delay_matrix_N_1_next_original[11]), 
        .ZN(n671) );
  ND2D1BWP30P140LVT U502 ( .A1(n1404), .A2(delay_matrix_N_1_next_original[10]), 
        .ZN(n669) );
  ND2D1BWP30P140LVT U503 ( .A1(n2194), .A2(delay_matrix_N_1_original[9]), .ZN(
        n569) );
  ND2D1BWP30P140LVT U504 ( .A1(n2194), .A2(delay_matrix_N_1_original[8]), .ZN(
        n567) );
  ND2D1BWP30P140LVT U505 ( .A1(n2194), .A2(delay_matrix_N_1_original[7]), .ZN(
        n1650) );
  ND2D1BWP30P140LVT U506 ( .A1(n2194), .A2(delay_matrix_N_1_original[6]), .ZN(
        n1795) );
  ND2D1BWP30P140LVT U507 ( .A1(n2194), .A2(delay_matrix_N_1_original[5]), .ZN(
        n1783) );
  ND2D1BWP30P140LVT U508 ( .A1(n2194), .A2(delay_matrix_N_1_original[4]), .ZN(
        n1648) );
  ND2D1BWP30P140LVT U509 ( .A1(n2194), .A2(delay_matrix_N_1_original[3]), .ZN(
        n1677) );
  ND2D1BWP30P140LVT U510 ( .A1(n2194), .A2(delay_matrix_N_1_original[2]), .ZN(
        n1772) );
  ND2D1BWP30P140LVT U511 ( .A1(n2194), .A2(delay_matrix_N_1_original[1]), .ZN(
        n1656) );
  ND2D1BWP30P140LVT U512 ( .A1(n2194), .A2(delay_matrix_N_1_original[0]), .ZN(
        n1770) );
  ND2D1BWP30P140LVT U513 ( .A1(n1398), .A2(delay_matrix_N_1_next_original[41]), 
        .ZN(n625) );
  ND2D1BWP30P140LVT U514 ( .A1(n1398), .A2(delay_matrix_N_1_next_original[40]), 
        .ZN(n627) );
  ND2D1BWP30P140LVT U515 ( .A1(n2204), .A2(delay_matrix_N_1_original[39]), 
        .ZN(n617) );
  ND2D1BWP30P140LVT U516 ( .A1(n1398), .A2(delay_matrix_N_1_next_original[39]), 
        .ZN(n670) );
  ND2D1BWP30P140LVT U517 ( .A1(n1398), .A2(delay_matrix_N_1_next_original[38]), 
        .ZN(n674) );
  ND2D1BWP30P140LVT U518 ( .A1(n2204), .A2(delay_matrix_N_1_original[37]), 
        .ZN(n580) );
  ND2D1BWP30P140LVT U519 ( .A1(n2204), .A2(delay_matrix_N_1_original[36]), 
        .ZN(n1775) );
  ND2D1BWP30P140LVT U520 ( .A1(n2204), .A2(delay_matrix_N_1_original[35]), 
        .ZN(n1658) );
  ND2D1BWP30P140LVT U521 ( .A1(n2204), .A2(delay_matrix_N_1_original[34]), 
        .ZN(n1652) );
  ND2D1BWP30P140LVT U522 ( .A1(n2204), .A2(delay_matrix_N_1_original[33]), 
        .ZN(n1787) );
  ND2D1BWP30P140LVT U523 ( .A1(n2204), .A2(delay_matrix_N_1_original[32]), 
        .ZN(n1768) );
  ND2D1BWP30P140LVT U524 ( .A1(n2204), .A2(delay_matrix_N_1_original[31]), 
        .ZN(n1641) );
  ND2D1BWP30P140LVT U525 ( .A1(n2204), .A2(delay_matrix_N_1_original[30]), 
        .ZN(n1809) );
  ND2D1BWP30P140LVT U526 ( .A1(n2204), .A2(delay_matrix_N_1_original[29]), 
        .ZN(n1662) );
  ND2D1BWP30P140LVT U527 ( .A1(n2204), .A2(delay_matrix_N_1_original[28]), 
        .ZN(n1667) );
  ND2D1BWP30P140LVT U528 ( .A1(n1333), .A2(delay_matrix_N_1_next_original[55]), 
        .ZN(n1332) );
  ND2D1BWP30P140LVT U529 ( .A1(n1333), .A2(delay_matrix_N_1_next_original[54]), 
        .ZN(n1334) );
  ND2D1BWP30P140LVT U530 ( .A1(n1801), .A2(delay_matrix_N_1_original[53]), 
        .ZN(n573) );
  ND2D1BWP30P140LVT U531 ( .A1(n1333), .A2(delay_matrix_N_1_next_original[53]), 
        .ZN(n1464) );
  ND2D1BWP30P140LVT U532 ( .A1(n1801), .A2(delay_matrix_N_1_original[52]), 
        .ZN(n571) );
  ND2D1BWP30P140LVT U533 ( .A1(n1333), .A2(delay_matrix_N_1_next_original[52]), 
        .ZN(n1198) );
  ND2D1BWP30P140LVT U534 ( .A1(n1801), .A2(delay_matrix_N_1_original[51]), 
        .ZN(n563) );
  ND2D1BWP30P140LVT U535 ( .A1(n1801), .A2(delay_matrix_N_1_original[50]), 
        .ZN(n1669) );
  ND2D1BWP30P140LVT U536 ( .A1(n1801), .A2(delay_matrix_N_1_original[49]), 
        .ZN(n1778) );
  ND2D1BWP30P140LVT U537 ( .A1(n1801), .A2(delay_matrix_N_1_original[48]), 
        .ZN(n1804) );
  ND2D1BWP30P140LVT U538 ( .A1(n1801), .A2(delay_matrix_N_1_original[47]), 
        .ZN(n1797) );
  ND2D1BWP30P140LVT U539 ( .A1(n1801), .A2(delay_matrix_N_1_original[46]), 
        .ZN(n1673) );
  ND2D1BWP30P140LVT U540 ( .A1(n1801), .A2(delay_matrix_N_1_original[45]), 
        .ZN(n1660) );
  ND2D1BWP30P140LVT U541 ( .A1(n1801), .A2(delay_matrix_N_1_original[44]), 
        .ZN(n1781) );
  ND2D1BWP30P140LVT U542 ( .A1(n1801), .A2(delay_matrix_N_1_original[43]), 
        .ZN(n1643) );
  ND2D1BWP30P140LVT U543 ( .A1(n1801), .A2(delay_matrix_N_1_original[42]), 
        .ZN(n1792) );
  ND2D1BWP30P140LVT U544 ( .A1(n1260), .A2(copy_ptr_next[8]), .ZN(n723) );
  ND2D1BWP30P140LVT U545 ( .A1(n1880), .A2(copy_ptr_next[18]), .ZN(n1882) );
  ND2D1BWP30P140LVT U546 ( .A1(n1873), .A2(copy_ptr_next[20]), .ZN(n1875) );
  ND2D1BWP30P140LVT U547 ( .A1(n1871), .A2(copy_ptr_next[22]), .ZN(n1868) );
  ND2D1BWP30P140LVT U548 ( .A1(n1859), .A2(copy_ptr_next[24]), .ZN(n1853) );
  MOAI22D1BWP30P140LVT U549 ( .A1(n1835), .A2(n235), .B1(n6), .B2(n237), .ZN(
        n924) );
  XNR2UD1BWP30P140LVT U550 ( .A1(n236), .A2(n235), .ZN(n237) );
  ND2D1BWP30P140LVT U551 ( .A1(n1618), .A2(n1760), .ZN(n1022) );
  ND2D1BWP30P140LVT U552 ( .A1(n1631), .A2(n1929), .ZN(n1236) );
  ND2D1BWP30P140LVT U553 ( .A1(n1322), .A2(n1760), .ZN(n1023) );
  ND2D1BWP30P140LVT U554 ( .A1(n1822), .A2(n1821), .ZN(n1024) );
  ND2D1BWP30P140LVT U555 ( .A1(n1949), .A2(n1929), .ZN(n697) );
  ND2D1BWP30P140LVT U556 ( .A1(n1983), .A2(n1929), .ZN(n1317) );
  ND2D1BWP30P140LVT U557 ( .A1(n1812), .A2(n1821), .ZN(n1026) );
  ND2D1BWP30P140LVT U558 ( .A1(n1962), .A2(n1929), .ZN(n711) );
  ND2D1BWP30P140LVT U559 ( .A1(n1958), .A2(n1929), .ZN(n1931) );
  ND2D1BWP30P140LVT U560 ( .A1(n1974), .A2(n1929), .ZN(n1921) );
  ND2D1BWP30P140LVT U561 ( .A1(n1966), .A2(n1929), .ZN(n1918) );
  ND2D1BWP30P140LVT U562 ( .A1(n1978), .A2(n1929), .ZN(n1924) );
  ND2D1BWP30P140LVT U563 ( .A1(n1970), .A2(n1929), .ZN(n1927) );
  ND2D1BWP30P140LVT U564 ( .A1(n2179), .A2(delay_matrix_N_1[11]), .ZN(n1628)
         );
  ND2D1BWP30P140LVT U565 ( .A1(n1624), .A2(n1760), .ZN(n1036) );
  ND2D1BWP30P140LVT U566 ( .A1(n2179), .A2(delay_matrix_N_1[10]), .ZN(n1632)
         );
  ND2D1BWP30P140LVT U567 ( .A1(n1305), .A2(n1760), .ZN(n1037) );
  ND2D1BWP30P140LVT U568 ( .A1(n2179), .A2(delay_matrix_N_1[9]), .ZN(n1757) );
  ND2D1BWP30P140LVT U569 ( .A1(n1816), .A2(n1821), .ZN(n1038) );
  ND2D1BWP30P140LVT U570 ( .A1(n2179), .A2(delay_matrix_N_1[8]), .ZN(n1563) );
  ND2D1BWP30P140LVT U571 ( .A1(n2179), .A2(delay_matrix_N_1[7]), .ZN(n1744) );
  ND2D1BWP30P140LVT U572 ( .A1(n1761), .A2(n1760), .ZN(n1040) );
  ND2D1BWP30P140LVT U573 ( .A1(n2179), .A2(delay_matrix_N_1[6]), .ZN(n1635) );
  ND2D1BWP30P140LVT U574 ( .A1(n2179), .A2(delay_matrix_N_1[5]), .ZN(n1690) );
  ND2D1BWP30P140LVT U575 ( .A1(n2179), .A2(delay_matrix_N_1[4]), .ZN(n678) );
  ND2D1BWP30P140LVT U576 ( .A1(n2179), .A2(delay_matrix_N_1[3]), .ZN(n651) );
  ND2D1BWP30P140LVT U577 ( .A1(n2179), .A2(delay_matrix_N_1[2]), .ZN(n620) );
  ND2D1BWP30P140LVT U578 ( .A1(n2179), .A2(delay_matrix_N_1[1]), .ZN(n1625) );
  ND2D1BWP30P140LVT U579 ( .A1(n2179), .A2(delay_matrix_N_1[0]), .ZN(n1645) );
  ND2D1BWP30P140LVT U580 ( .A1(n1755), .A2(n1754), .ZN(n978) );
  ND2D1BWP30P140LVT U581 ( .A1(n1591), .A2(n1590), .ZN(n979) );
  ND2D1BWP30P140LVT U582 ( .A1(n4), .A2(n1589), .ZN(n1590) );
  ND2D1BWP30P140LVT U583 ( .A1(n1639), .A2(n1760), .ZN(n1058) );
  ND2D1BWP30P140LVT U584 ( .A1(n1631), .A2(n1953), .ZN(n1239) );
  ND2D1BWP30P140LVT U585 ( .A1(n1323), .A2(n1760), .ZN(n1059) );
  ND2D1BWP30P140LVT U586 ( .A1(n1818), .A2(n1821), .ZN(n1060) );
  ND2D1BWP30P140LVT U587 ( .A1(n1949), .A2(n1953), .ZN(n1951) );
  ND2D1BWP30P140LVT U588 ( .A1(n1983), .A2(n1953), .ZN(n1320) );
  ND2D1BWP30P140LVT U589 ( .A1(n1811), .A2(n1821), .ZN(n1062) );
  ND2D1BWP30P140LVT U590 ( .A1(n1962), .A2(n1953), .ZN(n1935) );
  ND2D1BWP30P140LVT U591 ( .A1(n1958), .A2(n1953), .ZN(n1947) );
  ND2D1BWP30P140LVT U592 ( .A1(n1974), .A2(n1953), .ZN(n1955) );
  ND2D1BWP30P140LVT U593 ( .A1(n1966), .A2(n1953), .ZN(n1941) );
  ND2D1BWP30P140LVT U594 ( .A1(n1978), .A2(n1953), .ZN(n1944) );
  ND2D1BWP30P140LVT U595 ( .A1(n1970), .A2(n1953), .ZN(n1938) );
  ND2D1BWP30P140LVT U596 ( .A1(n2188), .A2(delay_matrix_N_1[28]), .ZN(n614) );
  ND2D1BWP30P140LVT U597 ( .A1(n1716), .A2(ptr_next[8]), .ZN(n1705) );
  ND2D1BWP30P140LVT U598 ( .A1(n1721), .A2(ptr_next[18]), .ZN(n1695) );
  ND2D1BWP30P140LVT U599 ( .A1(n1697), .A2(ptr_next[20]), .ZN(n1699) );
  ND2D1BWP30P140LVT U600 ( .A1(n1894), .A2(ptr_next[22]), .ZN(n1896) );
  ND2D1BWP30P140LVT U601 ( .A1(n1904), .A2(ptr_next[24]), .ZN(n1906) );
  MOAI22D1BWP30P140LVT U602 ( .A1(n473), .A2(n1835), .B1(n6), .B2(n475), .ZN(
        n1084) );
  XNR2UD1BWP30P140LVT U603 ( .A1(n474), .A2(n473), .ZN(n475) );
  ND2D1BWP30P140LVT U604 ( .A1(n1970), .A2(n1982), .ZN(n1972) );
  ND2D1BWP30P140LVT U605 ( .A1(n1978), .A2(n1982), .ZN(n1980) );
  ND2D1BWP30P140LVT U606 ( .A1(n1966), .A2(n1982), .ZN(n1968) );
  ND2D1BWP30P140LVT U607 ( .A1(n1974), .A2(n1982), .ZN(n1976) );
  ND2D1BWP30P140LVT U608 ( .A1(n1958), .A2(n1982), .ZN(n1960) );
  ND2D1BWP30P140LVT U609 ( .A1(n1962), .A2(n1982), .ZN(n1964) );
  ND2D1BWP30P140LVT U610 ( .A1(n1983), .A2(n1982), .ZN(n1986) );
  ND2D1BWP30P140LVT U611 ( .A1(n1756), .A2(n1821), .ZN(n1076) );
  ND2D1BWP30P140LVT U612 ( .A1(n1949), .A2(n1982), .ZN(n714) );
  ND2D1BWP30P140LVT U613 ( .A1(n1814), .A2(n1821), .ZN(n1074) );
  ND2D1BWP30P140LVT U614 ( .A1(n1631), .A2(n1982), .ZN(n1251) );
  ND2D1BWP30P140LVT U615 ( .A1(n1617), .A2(n1760), .ZN(n1072) );
  ND2D1BWP30P140LVT U616 ( .A1(n1527), .A2(copy_pointer[20]), .ZN(n1499) );
  ND2D1BWP30P140LVT U617 ( .A1(n1582), .A2(copy_pointer[22]), .ZN(n1533) );
  ND2D1BWP30P140LVT U618 ( .A1(n1545), .A2(copy_pointer[24]), .ZN(n1522) );
  XNR2UD1BWP30P140LVT U619 ( .A1(n1837), .A2(n1839), .ZN(n1838) );
  ND2D1BWP30P140LVT U620 ( .A1(n1454), .A2(pointer[18]), .ZN(n1455) );
  ND2D1BWP30P140LVT U621 ( .A1(n1440), .A2(pointer[20]), .ZN(n1441) );
  ND2D1BWP30P140LVT U622 ( .A1(n1436), .A2(pointer[22]), .ZN(n1437) );
  ND2D1BWP30P140LVT U623 ( .A1(n1449), .A2(pointer[24]), .ZN(n1446) );
  MOAI22D1BWP30P140LVT U624 ( .A1(n221), .A2(n1748), .B1(n4), .B2(n220), .ZN(
        n1148) );
  XNR2UD1BWP30P140LVT U625 ( .A1(n219), .A2(n221), .ZN(n220) );
  XNR2OPTND2BWP30P140LVT U626 ( .A1(n1315), .A2(n1314), .ZN(n1983) );
  NR2D1BWP30P140LVT U627 ( .A1(n2191), .A2(n1751), .ZN(n1752) );
  INVD1BWP30P140LVT U628 ( .I(n154), .ZN(n159) );
  INR2D2BWP30P140LVT U629 ( .A1(group_header[1]), .B1(group_header[0]), .ZN(
        n125) );
  INVD2BWP30P140LVT U630 ( .I(n2084), .ZN(n2086) );
  XNR2UD1BWP30P140LVT U631 ( .A1(n1412), .A2(n1411), .ZN(n1820) );
  INVD1BWP30P140LVT U632 ( .I(n1245), .ZN(n1748) );
  OR2D1BWP30P140LVT U633 ( .A1(n2172), .A2(n206), .Z(n1191) );
  ND2OPTIBD1BWP30P140LVT U634 ( .A1(n110), .A2(n109), .ZN(n2090) );
  INR2D1BWP30P140LVT U635 ( .A1(n206), .B1(n2172), .ZN(n1245) );
  CKAN2D1BWP30P140LVT U636 ( .A1(n101), .A2(n100), .Z(n12) );
  INVD1BWP30P140LVT U637 ( .I(n5), .ZN(n1802) );
  INVD1BWP30P140LVT U638 ( .I(n5), .ZN(n1773) );
  OR2D1BWP30P140LVT U639 ( .A1(n222), .A2(n1280), .Z(n13) );
  ND2OPTIBD1BWP30P140LVT U640 ( .A1(n130), .A2(n129), .ZN(n2102) );
  OR2D1BWP30P140LVT U641 ( .A1(reset), .A2(glob_scen_noc_input_valid), .Z(
        n1835) );
  INVD1BWP30P140LVT U642 ( .I(n2099), .ZN(n2121) );
  CKAN2D1BWP30P140LVT U643 ( .A1(n218), .A2(n1343), .Z(n14) );
  CKAN2D1BWP30P140LVT U644 ( .A1(n1492), .A2(n1495), .Z(n15) );
  CKAN2D1BWP30P140LVT U645 ( .A1(n234), .A2(n742), .Z(n16) );
  CKAN2D1BWP30P140LVT U646 ( .A1(n472), .A2(n1681), .Z(n17) );
  INVD1BWP30P140LVT U647 ( .I(n2085), .ZN(n2014) );
  INVD1BWP30P140LVT U648 ( .I(n2085), .ZN(n2155) );
  OR3D1BWP30P140LVT U649 ( .A1(n193), .A2(n192), .A3(n191), .Z(n18) );
  CKAN2D1BWP30P140LVT U650 ( .A1(n323), .A2(n322), .Z(n19) );
  OR2D1BWP30P140LVT U651 ( .A1(n168), .A2(n1987), .Z(n20) );
  INVD1BWP30P140LVT U652 ( .I(delay_matrix_element[13]), .ZN(n2203) );
  OR2D1BWP30P140LVT U653 ( .A1(group_header[0]), .A2(group_header[1]), .Z(n145) );
  INVD1BWP30P140LVT U654 ( .I(scenario_update), .ZN(n205) );
  INVD1BWP30P140LVT U655 ( .I(delay_matrix_element[0]), .ZN(n1793) );
  INVD1BWP30P140LVT U656 ( .I(reset), .ZN(n1821) );
  INVD1BWP30P140LVT U657 ( .I(delay_matrix_element[12]), .ZN(n2199) );
  INVD1BWP30P140LVT U658 ( .I(ptr_next[1]), .ZN(n1824) );
  TIELBWP30P140LVT U659 ( .ZN(n782) );
  INVD2BWP30P140LVT U660 ( .I(n9), .ZN(n405) );
  INVD2BWP30P140LVT U661 ( .I(table_ptr[1]), .ZN(n133) );
  NR2OPTPAD1BWP30P140LVT U662 ( .A1(n133), .A2(table_ptr[0]), .ZN(n22) );
  INVD2BWP30P140LVT U663 ( .I(n22), .ZN(n549) );
  INVD1BWP30P140LVT U664 ( .I(delay_matrix_N_1[17]), .ZN(n1919) );
  OAI22D1BWP30P140LVT U665 ( .A1(n549), .A2(n1969), .B1(n175), .B2(n1919), 
        .ZN(n21) );
  AOI21D1BWP30P140LVT U666 ( .A1(n405), .A2(delay_matrix_N_1[31]), .B(n21), 
        .ZN(n290) );
  INVD2BWP30P140LVT U667 ( .I(n22), .ZN(n174) );
  INVD3BWP30P140LVT U668 ( .I(n1989), .ZN(n500) );
  OAI22D1BWP30P140LVT U669 ( .A1(n174), .A2(n1297), .B1(n500), .B2(n1276), 
        .ZN(n23) );
  AOI22D1BWP30P140LVT U670 ( .A1(n503), .A2(delay_matrix_N_1[52]), .B1(n8), 
        .B2(delay_matrix_N_1[24]), .ZN(n25) );
  AOI22D1BWP30P140LVT U671 ( .A1(n503), .A2(delay_matrix_N_1[54]), .B1(n8), 
        .B2(delay_matrix_N_1[26]), .ZN(n27) );
  INVD1BWP30P140LVT U672 ( .I(n267), .ZN(n269) );
  OR4D1BWP30P140LVT U673 ( .A1(n290), .A2(n263), .A3(n279), .A4(n269), .Z(n30)
         );
  AOI22D1BWP30P140LVT U674 ( .A1(n503), .A2(delay_matrix_N_1[51]), .B1(n508), 
        .B2(delay_matrix_N_1[37]), .ZN(n28) );
  INVD1BWP30P140LVT U675 ( .I(n328), .ZN(n255) );
  OAI22D1BWP30P140LVT U676 ( .A1(n174), .A2(n1462), .B1(n175), .B2(n1243), 
        .ZN(n29) );
  NR3D0P7BWP30P140LVT U677 ( .A1(n30), .A2(n255), .A3(n273), .ZN(n42) );
  INVD1BWP30P140LVT U678 ( .I(delay_matrix_N_1[18]), .ZN(n1922) );
  OAI22D1BWP30P140LVT U679 ( .A1(n174), .A2(n1977), .B1(n175), .B2(n1922), 
        .ZN(n31) );
  AOI21D1BWP30P140LVT U680 ( .A1(n405), .A2(delay_matrix_N_1[32]), .B(n31), 
        .ZN(n294) );
  INVD1BWP30P140LVT U681 ( .I(delay_matrix_N_1[44]), .ZN(n1981) );
  INVD1BWP30P140LVT U682 ( .I(delay_matrix_N_1[16]), .ZN(n1925) );
  OAI22D1BWP30P140LVT U683 ( .A1(n174), .A2(n1981), .B1(n175), .B2(n1925), 
        .ZN(n32) );
  AOI21D1BWP30P140LVT U684 ( .A1(n405), .A2(delay_matrix_N_1[30]), .B(n32), 
        .ZN(n289) );
  INVD1BWP30P140LVT U685 ( .I(delay_matrix_N_1[43]), .ZN(n1973) );
  INVD1BWP30P140LVT U686 ( .I(delay_matrix_N_1[15]), .ZN(n1928) );
  OAI22D1BWP30P140LVT U687 ( .A1(n174), .A2(n1973), .B1(n175), .B2(n1928), 
        .ZN(n33) );
  AOI21D1BWP30P140LVT U688 ( .A1(n405), .A2(delay_matrix_N_1[29]), .B(n33), 
        .ZN(n244) );
  INVD1BWP30P140LVT U689 ( .I(delay_matrix_N_1[42]), .ZN(n702) );
  INVD1BWP30P140LVT U690 ( .I(delay_matrix_N_1[14]), .ZN(n639) );
  OAI22D1BWP30P140LVT U691 ( .A1(n174), .A2(n702), .B1(n175), .B2(n639), .ZN(
        n34) );
  AOI21D1BWP30P140LVT U692 ( .A1(n405), .A2(delay_matrix_N_1[28]), .B(n34), 
        .ZN(n243) );
  NR4D0BWP30P140LVT U693 ( .A1(n294), .A2(n289), .A3(n244), .A4(n243), .ZN(n41) );
  AOI22D1BWP30P140LVT U694 ( .A1(n503), .A2(delay_matrix_N_1[50]), .B1(n508), 
        .B2(delay_matrix_N_1[36]), .ZN(n36) );
  INVD1BWP30P140LVT U695 ( .I(delay_matrix_N_1[20]), .ZN(n712) );
  OAI22D1BWP30P140LVT U696 ( .A1(n174), .A2(n1965), .B1(n175), .B2(n712), .ZN(
        n37) );
  AOI21D1BWP30P140LVT U697 ( .A1(delay_matrix_N_1[34]), .A2(n405), .B(n37), 
        .ZN(n300) );
  INVD1BWP30P140LVT U698 ( .I(delay_matrix_N_1[21]), .ZN(n1318) );
  OAI22D1BWP30P140LVT U699 ( .A1(n174), .A2(n1987), .B1(n175), .B2(n1318), 
        .ZN(n38) );
  AOI21D1BWP30P140LVT U700 ( .A1(n405), .A2(delay_matrix_N_1[35]), .B(n38), 
        .ZN(n301) );
  INVD1BWP30P140LVT U701 ( .I(delay_matrix_N_1[19]), .ZN(n1932) );
  OAI22D1BWP30P140LVT U702 ( .A1(n174), .A2(n1961), .B1(n175), .B2(n1932), 
        .ZN(n39) );
  AOI21D1BWP30P140LVT U703 ( .A1(n405), .A2(delay_matrix_N_1[33]), .B(n39), 
        .ZN(n295) );
  NR4D0BWP30P140LVT U704 ( .A1(n240), .A2(n300), .A3(n301), .A4(n295), .ZN(n40) );
  AN2D2BWP30P140LVT U705 ( .A1(table_ptr[1]), .A2(table_ptr[0]), .Z(n373) );
  AOI31D1BWP30P140LVT U706 ( .A1(n42), .A2(n41), .A3(n40), .B(n373), .ZN(n496)
         );
  INVD2BWP30P140LVT U707 ( .I(reset), .ZN(n1760) );
  INVD2BWP30P140LVT U708 ( .I(n1760), .ZN(n1280) );
  ND2OPTIBD2BWP30P140LVT U709 ( .A1(n2000), .A2(n491), .ZN(n1991) );
  INR2D1BWP30P140LVT U710 ( .A1(n205), .B1(n1991), .ZN(n494) );
  NR2D1BWP30P140LVT U711 ( .A1(n548), .A2(table_ptr[0]), .ZN(N3860) );
  ND2OPTIBD2BWP30P140LVT U712 ( .A1(group_header[0]), .A2(group_header[1]), 
        .ZN(n168) );
  AOI21D1BWP30P140LVT U713 ( .A1(delay_matrix_N_1[39]), .A2(n125), .B(n43), 
        .ZN(n47) );
  INR2D2BWP30P140LVT U714 ( .A1(n45), .B1(n44), .ZN(n171) );
  INVD2BWP30P140LVT U715 ( .I(n145), .ZN(n170) );
  AOI22D1BWP30P140LVT U716 ( .A1(n171), .A2(delay_matrix_N_1[25]), .B1(n170), 
        .B2(delay_matrix_N_1[11]), .ZN(n46) );
  INVD1BWP30P140LVT U717 ( .I(delay_matrix_N_1[39]), .ZN(n1279) );
  OAI22D1BWP30P140LVT U718 ( .A1(n174), .A2(n1279), .B1(n1297), .B2(n7), .ZN(
        n50) );
  INR2D1BWP30P140LVT U719 ( .A1(delay_matrix_N_1[11]), .B1(n175), .ZN(n48) );
  NR3D0P7BWP30P140LVT U720 ( .A1(n50), .A2(n49), .A3(n48), .ZN(n2006) );
  AOI21D1BWP30P140LVT U721 ( .A1(delay_matrix_N_1[40]), .A2(n125), .B(n53), 
        .ZN(n55) );
  AOI22D1BWP30P140LVT U722 ( .A1(n171), .A2(delay_matrix_N_1[26]), .B1(n170), 
        .B2(delay_matrix_N_1[12]), .ZN(n54) );
  INVD1BWP30P140LVT U723 ( .I(delay_matrix_N_1[40]), .ZN(n1585) );
  OAI22D1BWP30P140LVT U724 ( .A1(n174), .A2(n1585), .B1(n1303), .B2(n7), .ZN(
        n59) );
  INVD1BWP30P140LVT U725 ( .I(delay_matrix_N_1[26]), .ZN(n1222) );
  INR2D1BWP30P140LVT U726 ( .A1(delay_matrix_N_1[12]), .B1(n175), .ZN(n57) );
  AOI21D1BWP30P140LVT U727 ( .A1(delay_matrix_N_1[38]), .A2(n125), .B(n61), 
        .ZN(n63) );
  AOI22D1BWP30P140LVT U728 ( .A1(n171), .A2(delay_matrix_N_1[24]), .B1(n170), 
        .B2(delay_matrix_N_1[10]), .ZN(n62) );
  INVD1BWP30P140LVT U729 ( .I(delay_matrix_N_1[38]), .ZN(n1240) );
  OAI22D1BWP30P140LVT U730 ( .A1(n174), .A2(n1240), .B1(n1252), .B2(n7), .ZN(
        n66) );
  INVD1BWP30P140LVT U731 ( .I(delay_matrix_N_1[24]), .ZN(n1237) );
  INR2D1BWP30P140LVT U732 ( .A1(delay_matrix_N_1[10]), .B1(n175), .ZN(n64) );
  AOI21D1BWP30P140LVT U733 ( .A1(n69), .A2(n189), .B(n76), .ZN(n67) );
  INVD1BWP30P140LVT U734 ( .I(n187), .ZN(n77) );
  AOI21D1BWP30P140LVT U735 ( .A1(delay_matrix_N_1[37]), .A2(n125), .B(n70), 
        .ZN(n72) );
  AOI22D1BWP30P140LVT U736 ( .A1(n171), .A2(delay_matrix_N_1[23]), .B1(n170), 
        .B2(delay_matrix_N_1[9]), .ZN(n71) );
  INVD1BWP30P140LVT U737 ( .I(delay_matrix_N_1[37]), .ZN(n1418) );
  OAI22D1BWP30P140LVT U738 ( .A1(n174), .A2(n1418), .B1(n1623), .B2(n7), .ZN(
        n75) );
  INVD1BWP30P140LVT U739 ( .I(delay_matrix_N_1[23]), .ZN(n1415) );
  INR2D1BWP30P140LVT U740 ( .A1(delay_matrix_N_1[9]), .B1(n175), .ZN(n73) );
  OR2D1BWP30P140LVT U741 ( .A1(n327), .A2(n2115), .Z(n84) );
  OAI21D1BWP30P140LVT U742 ( .A1(n77), .A2(n76), .B(n84), .ZN(n86) );
  AOI22D1BWP30P140LVT U743 ( .A1(n171), .A2(delay_matrix_N_1[22]), .B1(n170), 
        .B2(delay_matrix_N_1[8]), .ZN(n79) );
  MOAI22D1BWP30P140LVT U744 ( .A1(n168), .A2(n715), .B1(delay_matrix_N_1[36]), 
        .B2(n125), .ZN(n78) );
  INVD2BWP30P140LVT U745 ( .I(n549), .ZN(n507) );
  AOI21D1BWP30P140LVT U746 ( .A1(delay_matrix_N_1[36]), .A2(n507), .B(n80), 
        .ZN(n82) );
  AOI22D1BWP30P140LVT U747 ( .A1(n508), .A2(delay_matrix_N_1[22]), .B1(n8), 
        .B2(delay_matrix_N_1[8]), .ZN(n81) );
  AOI21D1BWP30P140LVT U748 ( .A1(n84), .A2(n186), .B(n83), .ZN(n85) );
  NR2D1BWP30P140LVT U749 ( .A1(n7), .A2(n1973), .ZN(n87) );
  AOI21D1BWP30P140LVT U750 ( .A1(delay_matrix_N_1[29]), .A2(n507), .B(n87), 
        .ZN(n89) );
  AOI22D1BWP30P140LVT U751 ( .A1(n508), .A2(delay_matrix_N_1[15]), .B1(n8), 
        .B2(delay_matrix_N_1[1]), .ZN(n88) );
  NR2D1BWP30P140LVT U752 ( .A1(n168), .A2(n1973), .ZN(n90) );
  AOI21D1BWP30P140LVT U753 ( .A1(delay_matrix_N_1[29]), .A2(n125), .B(n90), 
        .ZN(n92) );
  AOI22D1BWP30P140LVT U754 ( .A1(n171), .A2(delay_matrix_N_1[15]), .B1(n170), 
        .B2(delay_matrix_N_1[1]), .ZN(n91) );
  NR2D1BWP30P140LVT U755 ( .A1(n7), .A2(n702), .ZN(n93) );
  AOI21D1BWP30P140LVT U756 ( .A1(delay_matrix_N_1[28]), .A2(n507), .B(n93), 
        .ZN(n95) );
  AOI22D1BWP30P140LVT U757 ( .A1(n508), .A2(delay_matrix_N_1[14]), .B1(n8), 
        .B2(delay_matrix_N_1[0]), .ZN(n94) );
  NR2D1BWP30P140LVT U758 ( .A1(n168), .A2(n702), .ZN(n96) );
  AOI21D1BWP30P140LVT U759 ( .A1(delay_matrix_N_1[28]), .A2(n125), .B(n96), 
        .ZN(n98) );
  AOI22D1BWP30P140LVT U760 ( .A1(n171), .A2(delay_matrix_N_1[14]), .B1(n170), 
        .B2(delay_matrix_N_1[0]), .ZN(n97) );
  OAI22D1BWP30P140LVT U761 ( .A1(n2086), .A2(n2087), .B1(n2014), .B2(n2156), 
        .ZN(n113) );
  NR2D1BWP30P140LVT U762 ( .A1(n7), .A2(n1981), .ZN(n99) );
  AOI21D1BWP30P140LVT U763 ( .A1(delay_matrix_N_1[30]), .A2(n507), .B(n99), 
        .ZN(n101) );
  AOI22D1BWP30P140LVT U764 ( .A1(n508), .A2(delay_matrix_N_1[16]), .B1(n8), 
        .B2(delay_matrix_N_1[2]), .ZN(n100) );
  NR2D1BWP30P140LVT U765 ( .A1(n168), .A2(n1981), .ZN(n102) );
  AOI21D1BWP30P140LVT U766 ( .A1(delay_matrix_N_1[30]), .A2(n125), .B(n102), 
        .ZN(n104) );
  AOI22D1BWP30P140LVT U767 ( .A1(n171), .A2(delay_matrix_N_1[16]), .B1(n170), 
        .B2(delay_matrix_N_1[2]), .ZN(n103) );
  NR2D1BWP30P140LVT U768 ( .A1(n168), .A2(n1969), .ZN(n105) );
  AOI21D1BWP30P140LVT U769 ( .A1(delay_matrix_N_1[31]), .A2(n125), .B(n105), 
        .ZN(n107) );
  AOI22D1BWP30P140LVT U770 ( .A1(n171), .A2(delay_matrix_N_1[17]), .B1(n170), 
        .B2(delay_matrix_N_1[3]), .ZN(n106) );
  INVD2BWP30P140LVT U771 ( .I(n2092), .ZN(n115) );
  NR2D1BWP30P140LVT U772 ( .A1(n7), .A2(n1969), .ZN(n108) );
  AOI21D1BWP30P140LVT U773 ( .A1(delay_matrix_N_1[31]), .A2(n507), .B(n108), 
        .ZN(n110) );
  AOI22D1BWP30P140LVT U774 ( .A1(n508), .A2(delay_matrix_N_1[17]), .B1(n8), 
        .B2(delay_matrix_N_1[3]), .ZN(n109) );
  ND2OPTIBD1BWP30P140LVT U775 ( .A1(n115), .A2(n2090), .ZN(n114) );
  OAI21D1BWP30P140LVT U776 ( .A1(n12), .A2(n2088), .B(n114), .ZN(n111) );
  INVD1BWP30P140LVT U777 ( .I(n114), .ZN(n116) );
  OAI22D1BWP30P140LVT U778 ( .A1(n117), .A2(n116), .B1(n115), .B2(n2090), .ZN(
        n152) );
  AOI21D1BWP30P140LVT U779 ( .A1(delay_matrix_N_1[34]), .A2(n125), .B(n118), 
        .ZN(n120) );
  AOI22D1BWP30P140LVT U780 ( .A1(n171), .A2(delay_matrix_N_1[20]), .B1(n170), 
        .B2(delay_matrix_N_1[6]), .ZN(n119) );
  INVD1BWP30P140LVT U781 ( .I(n2100), .ZN(n124) );
  AOI21D1BWP30P140LVT U782 ( .A1(delay_matrix_N_1[34]), .A2(n507), .B(n121), 
        .ZN(n123) );
  AOI22D1BWP30P140LVT U783 ( .A1(n508), .A2(delay_matrix_N_1[20]), .B1(n8), 
        .B2(delay_matrix_N_1[6]), .ZN(n122) );
  ND2OPTIBD1BWP30P140LVT U784 ( .A1(n124), .A2(n2099), .ZN(n131) );
  AOI22D1BWP30P140LVT U785 ( .A1(n170), .A2(delay_matrix_N_1[7]), .B1(n125), 
        .B2(delay_matrix_N_1[35]), .ZN(n127) );
  ND2OPTIBD1BWP30P140LVT U786 ( .A1(n171), .A2(delay_matrix_N_1[21]), .ZN(n126) );
  ND3D2BWP30P140LVT U787 ( .A1(n20), .A2(n127), .A3(n126), .ZN(n2104) );
  AOI21D1BWP30P140LVT U788 ( .A1(delay_matrix_N_1[35]), .A2(n507), .B(n128), 
        .ZN(n130) );
  AOI22D1BWP30P140LVT U789 ( .A1(n508), .A2(delay_matrix_N_1[21]), .B1(n8), 
        .B2(delay_matrix_N_1[7]), .ZN(n129) );
  ND2OPTIBD1BWP30P140LVT U790 ( .A1(n3), .A2(n2102), .ZN(n160) );
  ND2OPTIBD1BWP30P140LVT U791 ( .A1(n131), .A2(n160), .ZN(n154) );
  AOI21D1BWP30P140LVT U792 ( .A1(delay_matrix_N_1[33]), .A2(n507), .B(n132), 
        .ZN(n136) );
  INR2D1BWP30P140LVT U793 ( .A1(delay_matrix_N_1[5]), .B1(table_ptr[0]), .ZN(
        n134) );
  AOI22D1BWP30P140LVT U794 ( .A1(n508), .A2(delay_matrix_N_1[19]), .B1(n134), 
        .B2(n133), .ZN(n135) );
  ND2OPTIBD1BWP30P140LVT U795 ( .A1(n171), .A2(delay_matrix_N_1[19]), .ZN(n138) );
  INVD2BWP30P140LVT U796 ( .I(n155), .ZN(n2098) );
  AOI21D1BWP30P140LVT U797 ( .A1(delay_matrix_N_1[32]), .A2(n507), .B(n142), 
        .ZN(n144) );
  AOI22D1BWP30P140LVT U798 ( .A1(n508), .A2(delay_matrix_N_1[18]), .B1(n8), 
        .B2(delay_matrix_N_1[4]), .ZN(n143) );
  INR2D1BWP30P140LVT U799 ( .A1(delay_matrix_N_1[4]), .B1(n145), .ZN(n146) );
  AOI21D1BWP30P140LVT U800 ( .A1(delay_matrix_N_1[32]), .A2(n125), .B(n146), 
        .ZN(n149) );
  AOI21D1BWP30P140LVT U801 ( .A1(n171), .A2(delay_matrix_N_1[18]), .B(n147), 
        .ZN(n148) );
  INR2D1BWP30P140LVT U802 ( .A1(n2093), .B1(n2094), .ZN(n150) );
  OAI22D1BWP30P140LVT U803 ( .A1(n157), .A2(n156), .B1(n155), .B2(n2096), .ZN(
        n158) );
  INVD1BWP30P140LVT U804 ( .I(n160), .ZN(n161) );
  OAI22D1BWP30P140LVT U805 ( .A1(n162), .A2(n161), .B1(n3), .B2(n2102), .ZN(
        n194) );
  ND2OPTIBD1BWP30P140LVT U806 ( .A1(n196), .A2(n163), .ZN(n167) );
  ND2OPTIBD2BWP30P140LVT U807 ( .A1(n167), .A2(n166), .ZN(n456) );
  NR2D1BWP30P140LVT U808 ( .A1(n168), .A2(n1462), .ZN(n169) );
  AOI21D1BWP30P140LVT U809 ( .A1(delay_matrix_N_1[41]), .A2(n125), .B(n169), 
        .ZN(n173) );
  AOI22D1BWP30P140LVT U810 ( .A1(n171), .A2(delay_matrix_N_1[27]), .B1(n170), 
        .B2(delay_matrix_N_1[13]), .ZN(n172) );
  INVD1BWP30P140LVT U811 ( .I(delay_matrix_N_1[41]), .ZN(n1747) );
  OAI22D1BWP30P140LVT U812 ( .A1(n174), .A2(n1747), .B1(n1462), .B2(n7), .ZN(
        n178) );
  INR2D1BWP30P140LVT U813 ( .A1(delay_matrix_N_1[13]), .B1(n175), .ZN(n176) );
  NR3D0P7BWP30P140LVT U814 ( .A1(n178), .A2(n177), .A3(n176), .ZN(n1996) );
  ND2OPTIBD1BWP30P140LVT U815 ( .A1(n274), .A2(n1996), .ZN(n188) );
  INVD1BWP30P140LVT U816 ( .I(n274), .ZN(n180) );
  INVD1BWP30P140LVT U817 ( .I(n1996), .ZN(n179) );
  NR3D0P7BWP30P140LVT U818 ( .A1(n195), .A2(n194), .A3(n18), .ZN(n197) );
  ND2OPTIBD2BWP30P140LVT U819 ( .A1(n197), .A2(n11), .ZN(n454) );
  ND3OPTPAD2BWP30P140LVT U820 ( .A1(n456), .A2(n198), .A3(n454), .ZN(n1994) );
  INR2D1BWP30P140LVT U821 ( .A1(n511), .B1(n1994), .ZN(n201) );
  INVD1BWP30P140LVT U822 ( .I(done2), .ZN(n199) );
  INR2D1BWP30P140LVT U823 ( .A1(n199), .B1(n1989), .ZN(n200) );
  AOI21D1BWP30P140LVT U824 ( .A1(n201), .A2(n200), .B(done), .ZN(n2002) );
  IOA22D2BWP30P140LVT U825 ( .B1(n202), .B2(n2002), .A1(n2001), .A2(
        table_ptr[0]), .ZN(n810) );
  INVD1BWP30P140LVT U826 ( .I(pointer[31]), .ZN(n221) );
  ND2D3BWP30P140LVT U827 ( .A1(n1760), .A2(n205), .ZN(n2172) );
  NR2D1BWP30P140LVT U828 ( .A1(n1430), .A2(n207), .ZN(n1422) );
  ND2D1BWP30P140LVT U829 ( .A1(pointer[22]), .A2(pointer[23]), .ZN(n208) );
  NR2D1BWP30P140LVT U830 ( .A1(n1426), .A2(n208), .ZN(n209) );
  NR2D1BWP30P140LVT U831 ( .A1(n1444), .A2(n210), .ZN(n218) );
  NR2D1BWP30P140LVT U832 ( .A1(n1362), .A2(n211), .ZN(n1348) );
  NR2D1BWP30P140LVT U833 ( .A1(n1349), .A2(n212), .ZN(n213) );
  NR2D1BWP30P140LVT U834 ( .A1(n1339), .A2(n214), .ZN(n216) );
  NR2D1BWP30P140LVT U835 ( .A1(n1187), .A2(n215), .ZN(n1217) );
  BUFFD6BWP30P140LVT U836 ( .I(n2232), .Z(prefetch_bypass_start_addr[8]) );
  NR2D1BWP30P140LVT U837 ( .A1(n1877), .A2(n223), .ZN(n1861) );
  NR2D1BWP30P140LVT U838 ( .A1(n1865), .A2(n224), .ZN(n225) );
  NR2D1BWP30P140LVT U839 ( .A1(n1851), .A2(n226), .ZN(n234) );
  NR2D1BWP30P140LVT U840 ( .A1(n717), .A2(n227), .ZN(n725) );
  NR2D1BWP30P140LVT U841 ( .A1(n733), .A2(n228), .ZN(n229) );
  NR2D1BWP30P140LVT U842 ( .A1(n1256), .A2(n230), .ZN(n232) );
  INVD1BWP30P140LVT U843 ( .I(copy_ptr_next[31]), .ZN(n235) );
  NR2D1BWP30P140LVT U844 ( .A1(n2087), .A2(n244), .ZN(n246) );
  NR2D1BWP30P140LVT U845 ( .A1(n2156), .A2(n243), .ZN(n245) );
  MOAI22D1BWP30P140LVT U846 ( .A1(n246), .A2(n245), .B1(n244), .B2(n2087), 
        .ZN(n249) );
  NR2D1BWP30P140LVT U847 ( .A1(n2088), .A2(n289), .ZN(n247) );
  INVD1BWP30P140LVT U848 ( .I(n317), .ZN(n254) );
  NR2D1BWP30P140LVT U849 ( .A1(n2094), .A2(n294), .ZN(n251) );
  INVD1BWP30P140LVT U850 ( .I(n316), .ZN(n253) );
  INR2D1BWP30P140LVT U851 ( .A1(n321), .B1(n308), .ZN(n288) );
  INVD1BWP30P140LVT U852 ( .I(n330), .ZN(n260) );
  INVD1BWP30P140LVT U853 ( .I(n327), .ZN(n258) );
  INVD1BWP30P140LVT U854 ( .I(n256), .ZN(n257) );
  INVD1BWP30P140LVT U855 ( .I(n283), .ZN(n259) );
  NR2D1BWP30P140LVT U856 ( .A1(n260), .A2(n259), .ZN(n261) );
  XNR2UD1BWP30P140LVT U857 ( .A1(n261), .A2(n332), .ZN(n272) );
  AOI21D1BWP30P140LVT U858 ( .A1(n263), .A2(n262), .B(n340), .ZN(n266) );
  INVD1BWP30P140LVT U859 ( .I(n278), .ZN(n265) );
  XNR2UD1BWP30P140LVT U860 ( .A1(n266), .A2(n280), .ZN(n325) );
  XNR2UD1BWP30P140LVT U861 ( .A1(n271), .A2(n340), .ZN(n326) );
  NR2D1BWP30P140LVT U862 ( .A1(n274), .A2(n273), .ZN(n275) );
  INR2D1BWP30P140LVT U863 ( .A1(n335), .B1(n275), .ZN(n338) );
  INVD1BWP30P140LVT U864 ( .I(n338), .ZN(n277) );
  MUX2NUD1BWP30P140LVT U865 ( .I0(n335), .I1(n277), .S(n276), .ZN(n285) );
  INVD1BWP30P140LVT U866 ( .I(n280), .ZN(n281) );
  INR2D1BWP30P140LVT U867 ( .A1(n282), .B1(n281), .ZN(n329) );
  ND2OPTIBD1BWP30P140LVT U868 ( .A1(n285), .A2(n284), .ZN(n286) );
  NR3D1P5BWP30P140LVT U869 ( .A1(n288), .A2(n287), .A3(n286), .ZN(n314) );
  ND2OPTIBD1BWP30P140LVT U870 ( .A1(n2092), .A2(n290), .ZN(n291) );
  NR2D1BWP30P140LVT U871 ( .A1(n316), .A2(n318), .ZN(n310) );
  INVD1BWP30P140LVT U872 ( .I(n2098), .ZN(n297) );
  INVD1BWP30P140LVT U873 ( .I(n295), .ZN(n296) );
  OAI22D1BWP30P140LVT U874 ( .A1(n299), .A2(n298), .B1(n297), .B2(n296), .ZN(
        n306) );
  INVD1BWP30P140LVT U875 ( .I(n301), .ZN(n302) );
  OAI22D1BWP30P140LVT U876 ( .A1(n304), .A2(n303), .B1(n302), .B2(n3), .ZN(
        n305) );
  AOI21D1BWP30P140LVT U877 ( .A1(n307), .A2(n306), .B(n305), .ZN(n323) );
  ND3D1BWP30P140LVT U878 ( .A1(n309), .A2(n323), .A3(n308), .ZN(n313) );
  INR2D1BWP30P140LVT U879 ( .A1(n321), .B1(n323), .ZN(n319) );
  INR2D1BWP30P140LVT U880 ( .A1(n311), .B1(n319), .ZN(n312) );
  ND3OPTPAD2BWP30P140LVT U881 ( .A1(n314), .A2(n313), .A3(n312), .ZN(n315) );
  AOI21D1BWP30P140LVT U882 ( .A1(n318), .A2(n317), .B(n316), .ZN(n320) );
  AOI21D1BWP30P140LVT U883 ( .A1(n320), .A2(n321), .B(n319), .ZN(n347) );
  INVD1BWP30P140LVT U884 ( .I(n320), .ZN(n324) );
  INVD1BWP30P140LVT U885 ( .I(n321), .ZN(n322) );
  ND2OPTIBD1BWP30P140LVT U886 ( .A1(n326), .A2(n325), .ZN(n344) );
  XOR2UD1BWP30P140LVT U887 ( .A1(n329), .A2(n331), .Z(n343) );
  INVD1BWP30P140LVT U888 ( .I(n332), .ZN(n333) );
  XNR2UD1BWP30P140LVT U889 ( .A1(n334), .A2(n333), .ZN(n337) );
  AOI31D1BWP30P140LVT U890 ( .A1(n340), .A2(n339), .A3(n335), .B(n500), .ZN(
        n336) );
  ND2OPTIBD1BWP30P140LVT U891 ( .A1(n337), .A2(n336), .ZN(n342) );
  AOI21D1BWP30P140LVT U892 ( .A1(n340), .A2(n339), .B(n338), .ZN(n341) );
  NR4D1BWP30P140LVT U893 ( .A1(n344), .A2(n343), .A3(n342), .A4(n341), .ZN(
        n345) );
  INVD1BWP30P140LVT U894 ( .I(scenario_len[1]), .ZN(n356) );
  AOI22D1BWP30P140LVT U895 ( .A1(n373), .A2(delay_matrix_N_1_original[43]), 
        .B1(n508), .B2(delay_matrix_N_1_original[15]), .ZN(n350) );
  AOI22D1BWP30P140LVT U896 ( .A1(n503), .A2(delay_matrix_N_1_original[29]), 
        .B1(n8), .B2(delay_matrix_N_1_original[1]), .ZN(n349) );
  ND2D1BWP30P140LVT U897 ( .A1(n350), .A2(n349), .ZN(n357) );
  INVD1BWP30P140LVT U898 ( .I(delay_matrix_N_1_original[42]), .ZN(n351) );
  NR2D1BWP30P140LVT U899 ( .A1(n7), .A2(n351), .ZN(n352) );
  AOI21D1BWP30P140LVT U900 ( .A1(n8), .A2(delay_matrix_N_1_original[0]), .B(
        n352), .ZN(n355) );
  INVD1BWP30P140LVT U901 ( .I(delay_matrix_N_1_original[14]), .ZN(n1765) );
  OAI21D1BWP30P140LVT U902 ( .A1(n9), .A2(n1765), .B(scenario_len[0]), .ZN(
        n353) );
  AOI21D1BWP30P140LVT U903 ( .A1(n507), .A2(delay_matrix_N_1_original[28]), 
        .B(n353), .ZN(n354) );
  MOAI22D1BWP30P140LVT U904 ( .A1(n356), .A2(n357), .B1(n355), .B2(n354), .ZN(
        n368) );
  ND2D1BWP30P140LVT U905 ( .A1(n357), .A2(n356), .ZN(n361) );
  AOI22D1BWP30P140LVT U906 ( .A1(n373), .A2(delay_matrix_N_1_original[45]), 
        .B1(n508), .B2(delay_matrix_N_1_original[17]), .ZN(n359) );
  AOI22D1BWP30P140LVT U907 ( .A1(n503), .A2(delay_matrix_N_1_original[31]), 
        .B1(n8), .B2(delay_matrix_N_1_original[3]), .ZN(n358) );
  ND2D1BWP30P140LVT U908 ( .A1(n359), .A2(n358), .ZN(n372) );
  INVD1BWP30P140LVT U909 ( .I(scenario_len[3]), .ZN(n371) );
  NR2D1BWP30P140LVT U910 ( .A1(n372), .A2(n371), .ZN(n360) );
  AOI31D1BWP30P140LVT U911 ( .A1(n368), .A2(scenario_len[2]), .A3(n361), .B(
        n360), .ZN(n384) );
  INVD1BWP30P140LVT U912 ( .I(n361), .ZN(n366) );
  INVD1BWP30P140LVT U913 ( .I(scenario_len[2]), .ZN(n365) );
  AOI22D1BWP30P140LVT U914 ( .A1(n373), .A2(delay_matrix_N_1_original[44]), 
        .B1(n508), .B2(delay_matrix_N_1_original[16]), .ZN(n363) );
  AOI22D1BWP30P140LVT U915 ( .A1(n503), .A2(delay_matrix_N_1_original[30]), 
        .B1(n8), .B2(delay_matrix_N_1_original[2]), .ZN(n362) );
  ND2D1BWP30P140LVT U916 ( .A1(n363), .A2(n362), .ZN(n364) );
  AOI21D1BWP30P140LVT U917 ( .A1(n366), .A2(n365), .B(n364), .ZN(n367) );
  OAI21D1BWP30P140LVT U918 ( .A1(scenario_len[2]), .A2(n368), .B(n367), .ZN(
        n383) );
  INVD1BWP30P140LVT U919 ( .I(scenario_len[4]), .ZN(n415) );
  AOI22D1BWP30P140LVT U920 ( .A1(n373), .A2(delay_matrix_N_1_original[46]), 
        .B1(n503), .B2(delay_matrix_N_1_original[32]), .ZN(n370) );
  AOI22D1BWP30P140LVT U921 ( .A1(n508), .A2(delay_matrix_N_1_original[18]), 
        .B1(n8), .B2(delay_matrix_N_1_original[4]), .ZN(n369) );
  ND2D1BWP30P140LVT U922 ( .A1(n370), .A2(n369), .ZN(n416) );
  AOI22D1BWP30P140LVT U923 ( .A1(n415), .A2(n416), .B1(n372), .B2(n371), .ZN(
        n381) );
  AOI22D1BWP30P140LVT U924 ( .A1(n373), .A2(delay_matrix_N_1_original[48]), 
        .B1(n503), .B2(delay_matrix_N_1_original[34]), .ZN(n375) );
  AOI22D1BWP30P140LVT U925 ( .A1(n508), .A2(delay_matrix_N_1_original[20]), 
        .B1(n8), .B2(delay_matrix_N_1_original[6]), .ZN(n374) );
  ND2D1BWP30P140LVT U926 ( .A1(n375), .A2(n374), .ZN(n409) );
  INVD1BWP30P140LVT U927 ( .I(scenario_len[6]), .ZN(n408) );
  INVD1BWP30P140LVT U928 ( .I(delay_matrix_N_1_original[47]), .ZN(n376) );
  NR2D1BWP30P140LVT U929 ( .A1(n7), .A2(n376), .ZN(n377) );
  AOI21D1BWP30P140LVT U930 ( .A1(n8), .A2(delay_matrix_N_1_original[5]), .B(
        n377), .ZN(n379) );
  ND2D1BWP30P140LVT U931 ( .A1(n405), .A2(delay_matrix_N_1_original[19]), .ZN(
        n378) );
  ND2D1BWP30P140LVT U932 ( .A1(n379), .A2(n378), .ZN(n414) );
  INR2D1BWP30P140LVT U933 ( .A1(delay_matrix_N_1_original[33]), .B1(n549), 
        .ZN(n411) );
  INVD1BWP30P140LVT U934 ( .I(scenario_len[5]), .ZN(n380) );
  OAI21D1BWP30P140LVT U935 ( .A1(n414), .A2(n411), .B(n380), .ZN(n417) );
  ND3D1BWP30P140LVT U936 ( .A1(n381), .A2(n418), .A3(n417), .ZN(n382) );
  AOI21D1BWP30P140LVT U937 ( .A1(n384), .A2(n383), .B(n382), .ZN(n451) );
  INVD1BWP30P140LVT U938 ( .I(delay_matrix_N_1_original[36]), .ZN(n386) );
  INVD1BWP30P140LVT U939 ( .I(delay_matrix_N_1_original[50]), .ZN(n385) );
  OAI22D1BWP30P140LVT U940 ( .A1(n549), .A2(n386), .B1(n7), .B2(n385), .ZN(
        n388) );
  INVD1BWP30P140LVT U941 ( .I(delay_matrix_N_1_original[22]), .ZN(n677) );
  NR2D1BWP30P140LVT U942 ( .A1(n9), .A2(n677), .ZN(n387) );
  AOI211D1BWP30P140LVT U943 ( .A1(n1989), .A2(delay_matrix_N_1_original[8]), 
        .B(n388), .C(n387), .ZN(n422) );
  INVD1BWP30P140LVT U944 ( .I(delay_matrix_N_1_original[9]), .ZN(n390) );
  INVD1BWP30P140LVT U945 ( .I(delay_matrix_N_1_original[51]), .ZN(n389) );
  OAI22D1BWP30P140LVT U946 ( .A1(n500), .A2(n390), .B1(n7), .B2(n389), .ZN(
        n391) );
  AOI21OPTREPBD1BWP30P140LVT U947 ( .A1(n405), .A2(
        delay_matrix_N_1_original[23]), .B(n391), .ZN(n429) );
  INVD1BWP30P140LVT U948 ( .I(n429), .ZN(n394) );
  INVD1BWP30P140LVT U949 ( .I(n428), .ZN(n393) );
  INVD1BWP30P140LVT U950 ( .I(scenario_len[9]), .ZN(n392) );
  NR3D0P7BWP30P140LVT U951 ( .A1(n394), .A2(n393), .A3(n392), .ZN(n395) );
  AOI21D1BWP30P140LVT U952 ( .A1(n422), .A2(scenario_len[8]), .B(n395), .ZN(
        n401) );
  INVD1BWP30P140LVT U953 ( .I(delay_matrix_N_1_original[38]), .ZN(n397) );
  INVD1BWP30P140LVT U954 ( .I(delay_matrix_N_1_original[52]), .ZN(n396) );
  OAI22D1BWP30P140LVT U955 ( .A1(n549), .A2(n397), .B1(n7), .B2(n396), .ZN(
        n400) );
  INVD1BWP30P140LVT U956 ( .I(delay_matrix_N_1_original[24]), .ZN(n398) );
  NR2D1BWP30P140LVT U957 ( .A1(n9), .A2(n398), .ZN(n399) );
  INVD1BWP30P140LVT U958 ( .I(delay_matrix_N_1_original[7]), .ZN(n403) );
  INVD1BWP30P140LVT U959 ( .I(delay_matrix_N_1_original[49]), .ZN(n402) );
  OAI22D1BWP30P140LVT U960 ( .A1(n500), .A2(n403), .B1(n7), .B2(n402), .ZN(
        n404) );
  AOI21D1BWP30P140LVT U961 ( .A1(n405), .A2(delay_matrix_N_1_original[21]), 
        .B(n404), .ZN(n424) );
  INVD1BWP30P140LVT U962 ( .I(n424), .ZN(n407) );
  ND2D1BWP30P140LVT U963 ( .A1(n503), .A2(delay_matrix_N_1_original[35]), .ZN(
        n423) );
  ND2D1BWP30P140LVT U964 ( .A1(n423), .A2(scenario_len[7]), .ZN(n406) );
  OAI22D1BWP30P140LVT U965 ( .A1(n409), .A2(n408), .B1(n407), .B2(n406), .ZN(
        n410) );
  NR2D1BWP30P140LVT U966 ( .A1(n446), .A2(n410), .ZN(n421) );
  INVD1BWP30P140LVT U967 ( .I(n411), .ZN(n412) );
  ND2D1BWP30P140LVT U968 ( .A1(n412), .A2(scenario_len[5]), .ZN(n413) );
  OAI22D1BWP30P140LVT U969 ( .A1(n416), .A2(n415), .B1(n414), .B2(n413), .ZN(
        n419) );
  ND3D1BWP30P140LVT U970 ( .A1(n419), .A2(n418), .A3(n417), .ZN(n420) );
  INVD1BWP30P140LVT U971 ( .I(scenario_len[8]), .ZN(n427) );
  INVD1BWP30P140LVT U972 ( .I(n422), .ZN(n426) );
  AOI21D1BWP30P140LVT U973 ( .A1(n424), .A2(n423), .B(scenario_len[7]), .ZN(
        n425) );
  AOI21D1BWP30P140LVT U974 ( .A1(n427), .A2(n426), .B(n425), .ZN(n445) );
  AOI21D1BWP30P140LVT U975 ( .A1(n429), .A2(n428), .B(scenario_len[9]), .ZN(
        n443) );
  NR2D1BWP30P140LVT U976 ( .A1(delay_matrix_N_1_original[40]), .A2(
        delay_matrix_N_1_original[41]), .ZN(n430) );
  INVD1BWP30P140LVT U977 ( .I(delay_matrix_N_1_original[25]), .ZN(n431) );
  NR2D1BWP30P140LVT U978 ( .A1(n9), .A2(n431), .ZN(n432) );
  AOI211D1BWP30P140LVT U979 ( .A1(n1989), .A2(delay_matrix_N_1_original[11]), 
        .B(n433), .C(n432), .ZN(n439) );
  IAO21D1BWP30P140LVT U980 ( .A1(delay_matrix_N_1_original[13]), .A2(
        delay_matrix_N_1_original[12]), .B(n500), .ZN(n437) );
  NR2D1BWP30P140LVT U981 ( .A1(delay_matrix_N_1_original[55]), .A2(
        delay_matrix_N_1_original[54]), .ZN(n435) );
  INVD1BWP30P140LVT U982 ( .I(delay_matrix_N_1_original[53]), .ZN(n434) );
  AOI21D1BWP30P140LVT U983 ( .A1(n435), .A2(n434), .B(n7), .ZN(n436) );
  AOI211D1BWP30P140LVT U984 ( .A1(n507), .A2(delay_matrix_N_1_original[39]), 
        .B(n437), .C(n436), .ZN(n438) );
  OAI21D1BWP30P140LVT U985 ( .A1(n446), .A2(n445), .B(n444), .ZN(n448) );
  INVD1BWP30P140LVT U986 ( .I(n448), .ZN(n447) );
  OAI21D1BWP30P140LVT U987 ( .A1(n451), .A2(n450), .B(n447), .ZN(n522) );
  INR2D1BWP30P140LVT U988 ( .A1(n494), .B1(n522), .ZN(n518) );
  NR2OPTPAD1BWP30P140LVT U989 ( .A1(n448), .A2(n521), .ZN(n449) );
  OAI21OPTREPBD1BWP30P140LVT U990 ( .A1(n451), .A2(n450), .B(n449), .ZN(n453)
         );
  ND3OPTPAD2BWP30P140LVT U991 ( .A1(n456), .A2(n455), .A3(n454), .ZN(n515) );
  NR3D3BWP30P140LVT U992 ( .A1(n457), .A2(n524), .A3(n515), .ZN(n2176) );
  INR2D1BWP30P140LVT U993 ( .A1(prefetch_bypass_start_addr[13]), .B1(n2172), 
        .ZN(n459) );
  NR2D1BWP30P140LVT U994 ( .A1(n1693), .A2(n461), .ZN(n1685) );
  NR2D1BWP30P140LVT U995 ( .A1(n1687), .A2(n462), .ZN(n463) );
  NR2D1BWP30P140LVT U996 ( .A1(n1682), .A2(n464), .ZN(n472) );
  NR2D1BWP30P140LVT U997 ( .A1(n1714), .A2(n465), .ZN(n1710) );
  NR2D1BWP30P140LVT U998 ( .A1(n1711), .A2(n466), .ZN(n467) );
  NR2D1BWP30P140LVT U999 ( .A1(n1474), .A2(n468), .ZN(n470) );
  INVD1BWP30P140LVT U1000 ( .I(ptr_next[31]), .ZN(n473) );
  INVD2BWP30P140LVT U1001 ( .I(n2231), .ZN(n476) );
  INVD9BWP30P140LVT U1002 ( .I(n476), .ZN(prefetch_bypass_start_addr[11]) );
  INVD9BWP30P140LVT U1003 ( .I(n477), .ZN(prefetch_bypass_start_addr[0]) );
  NR4D0BWP30P140LVT U1004 ( .A1(copy_pointer[2]), .A2(copy_pointer[6]), .A3(
        copy_pointer[8]), .A4(copy_pointer[18]), .ZN(n478) );
  INVD1BWP30P140LVT U1005 ( .I(copy_pointer[31]), .ZN(n1839) );
  INVD1BWP30P140LVT U1006 ( .I(copy_pointer[30]), .ZN(n1507) );
  ND3D1BWP30P140LVT U1007 ( .A1(n478), .A2(n1839), .A3(n1507), .ZN(n486) );
  NR4D0BWP30P140LVT U1008 ( .A1(copy_pointer[22]), .A2(copy_pointer[20]), .A3(
        copy_pointer[3]), .A4(copy_pointer[24]), .ZN(n485) );
  NR4D0BWP30P140LVT U1009 ( .A1(copy_pointer[5]), .A2(copy_pointer[7]), .A3(
        copy_pointer[9]), .A4(copy_pointer[11]), .ZN(n484) );
  NR4D0BWP30P140LVT U1010 ( .A1(copy_pointer[15]), .A2(copy_pointer[13]), .A3(
        copy_pointer[17]), .A4(copy_pointer[19]), .ZN(n482) );
  NR4D0BWP30P140LVT U1011 ( .A1(copy_pointer[10]), .A2(copy_pointer[12]), .A3(
        copy_pointer[14]), .A4(copy_pointer[16]), .ZN(n481) );
  NR4D0BWP30P140LVT U1012 ( .A1(copy_pointer[29]), .A2(copy_pointer[28]), .A3(
        copy_pointer[27]), .A4(copy_pointer[26]), .ZN(n480) );
  NR4D0BWP30P140LVT U1013 ( .A1(copy_pointer[23]), .A2(copy_pointer[21]), .A3(
        copy_pointer[4]), .A4(copy_pointer[25]), .ZN(n479) );
  IND4D1BWP30P140LVT U1014 ( .A1(n486), .B1(n485), .B2(n484), .B3(n483), .ZN(
        n564) );
  OAI21D1BWP30P140LVT U1015 ( .A1(n487), .A2(n1191), .B(n1748), .ZN(n2204) );
  ND2OPTIBD2BWP30P140LVT U1016 ( .A1(n487), .A2(n4), .ZN(n2207) );
  INVD1BWP30P140LVT U1017 ( .I(n2207), .ZN(n489) );
  AOI22D1BWP30P140LVT U1018 ( .A1(n489), .A2(delay_matrix_element[12]), .B1(
        n1984), .B2(delay_matrix_N_1_next_original[40]), .ZN(n488) );
  IOA21D1BWP30P140LVT U1019 ( .A1(delay_matrix_N_1_original[40]), .A2(n2204), 
        .B(n488), .ZN(n827) );
  AOI22D1BWP30P140LVT U1020 ( .A1(n489), .A2(delay_matrix_element[13]), .B1(
        n1984), .B2(delay_matrix_N_1_next_original[41]), .ZN(n490) );
  IOA21D1BWP30P140LVT U1021 ( .A1(delay_matrix_N_1_original[41]), .A2(n2204), 
        .B(n490), .ZN(n826) );
  INVD1BWP30P140LVT U1022 ( .I(n491), .ZN(n492) );
  ND2D1BWP30P140LVT U1023 ( .A1(n492), .A2(table_parse), .ZN(n493) );
  NR2D1BWP30P140LVT U1024 ( .A1(n2121), .A2(n1991), .ZN(N4221) );
  NR2D1BWP30P140LVT U1025 ( .A1(n2086), .A2(n1991), .ZN(N4216) );
  NR2D1BWP30P140LVT U1026 ( .A1(n2103), .A2(n1991), .ZN(N4222) );
  NR2D1BWP30P140LVT U1027 ( .A1(n2097), .A2(n1991), .ZN(N4220) );
  NR2D1BWP30P140LVT U1028 ( .A1(n2), .A2(n1991), .ZN(N4219) );
  NR2D1BWP30P140LVT U1029 ( .A1(n2091), .A2(n1991), .ZN(N4218) );
  NR2D1BWP30P140LVT U1030 ( .A1(n2014), .A2(n1991), .ZN(N4215) );
  NR2D1BWP30P140LVT U1031 ( .A1(n12), .A2(n1991), .ZN(N4217) );
  INVD1BWP30P140LVT U1032 ( .I(n494), .ZN(n495) );
  NR2D1BWP30P140LVT U1033 ( .A1(n496), .A2(n495), .ZN(N3862) );
  AOI22D1BWP30P140LVT U1034 ( .A1(n508), .A2(obj_id[2]), .B1(n8), .B2(
        obj_id[0]), .ZN(n505) );
  INVD1BWP30P140LVT U1035 ( .I(obj_id[6]), .ZN(n744) );
  MOAI22D1BWP30P140LVT U1036 ( .A1(n7), .A2(n744), .B1(obj_id[4]), .B2(n503), 
        .ZN(n504) );
  INVD1BWP30P140LVT U1037 ( .I(n2069), .ZN(n2072) );
  INVD1BWP30P140LVT U1038 ( .I(obj_id[7]), .ZN(n746) );
  NR2D1BWP30P140LVT U1039 ( .A1(n7), .A2(n746), .ZN(n506) );
  AOI21D1BWP30P140LVT U1040 ( .A1(obj_id[5]), .A2(n507), .B(n506), .ZN(n510)
         );
  AOI22D1BWP30P140LVT U1041 ( .A1(n508), .A2(obj_id[3]), .B1(n8), .B2(
        obj_id[1]), .ZN(n509) );
  CKAN2D1BWP30P140LVT U1042 ( .A1(n512), .A2(n511), .Z(n513) );
  INVD2BWP30P140LVT U1043 ( .I(n2023), .ZN(n1995) );
  OAI31D1BWP30P140LVT U1044 ( .A1(n1991), .A2(n2072), .A3(n2075), .B(n514), 
        .ZN(N4197) );
  INR2D1BWP30P140LVT U1045 ( .A1(n2075), .B1(n1991), .ZN(n2225) );
  INVD1BWP30P140LVT U1046 ( .I(n515), .ZN(n520) );
  INVD1BWP30P140LVT U1047 ( .I(n516), .ZN(n519) );
  OAI21D1BWP30P140LVT U1048 ( .A1(n522), .A2(n521), .B(n700), .ZN(n523) );
  OAI31D1BWP30P140LVT U1049 ( .A1(n2069), .A2(n2075), .A3(n530), .B(n525), 
        .ZN(n807) );
  INVD1BWP30P140LVT U1050 ( .I(n2075), .ZN(n531) );
  OAI31D1BWP30P140LVT U1051 ( .A1(n531), .A2(n2072), .A3(n530), .B(n526), .ZN(
        n806) );
  OAI31D1BWP30P140LVT U1052 ( .A1(n2075), .A2(n2072), .A3(n530), .B(n527), 
        .ZN(n808) );
  OAI31D1BWP30P140LVT U1053 ( .A1(n2069), .A2(n531), .A3(n530), .B(n529), .ZN(
        n805) );
  NR4D0BWP30P140LVT U1054 ( .A1(ptr_next[15]), .A2(ptr_next[13]), .A3(
        ptr_next[11]), .A4(ptr_next[9]), .ZN(n536) );
  NR4D0BWP30P140LVT U1055 ( .A1(ptr_next[14]), .A2(ptr_next[12]), .A3(
        ptr_next[10]), .A4(ptr_next[4]), .ZN(n535) );
  NR4D0BWP30P140LVT U1056 ( .A1(ptr_next[29]), .A2(ptr_next[30]), .A3(
        ptr_next[27]), .A4(ptr_next[28]), .ZN(n534) );
  NR4D0BWP30P140LVT U1057 ( .A1(ptr_next[7]), .A2(ptr_next[5]), .A3(
        ptr_next[16]), .A4(ptr_next[3]), .ZN(n533) );
  ND4D1BWP30P140LVT U1058 ( .A1(n536), .A2(n535), .A3(n534), .A4(n533), .ZN(
        n542) );
  NR4D0BWP30P140LVT U1059 ( .A1(ptr_next[24]), .A2(ptr_next[22]), .A3(
        ptr_next[20]), .A4(ptr_next[18]), .ZN(n540) );
  NR4D0BWP30P140LVT U1060 ( .A1(ptr_next[23]), .A2(ptr_next[21]), .A3(
        ptr_next[19]), .A4(ptr_next[17]), .ZN(n539) );
  NR4D0BWP30P140LVT U1061 ( .A1(ptr_next[8]), .A2(ptr_next[6]), .A3(
        ptr_next[25]), .A4(ptr_next[2]), .ZN(n538) );
  ND4D1BWP30P140LVT U1062 ( .A1(n540), .A2(n539), .A3(n538), .A4(n537), .ZN(
        n541) );
  AOI21D1BWP30P140LVT U1063 ( .A1(n1813), .A2(delay_matrix_N_1_next[42]), .B(
        n1807), .ZN(n543) );
  OAI21D1BWP30P140LVT U1064 ( .A1(n1646), .A2(n1813), .B(n543), .ZN(n1083) );
  INVD1BWP30P140LVT U1065 ( .I(n553), .ZN(n545) );
  ND2OPTIBD1BWP30P140LVT U1066 ( .A1(n545), .A2(n551), .ZN(n546) );
  FA1D1BWP30P140LVT U1067 ( .A(hardware_latency2[0]), .B(hardware_latency1[0]), 
        .CI(delay_matrix_element[0]), .CO(n550), .S(n532) );
  AOI21D1BWP30P140LVT U1068 ( .A1(n1813), .A2(delay_matrix_N_1_next[43]), .B(
        n1807), .ZN(n547) );
  OAI21D1BWP30P140LVT U1069 ( .A1(n1627), .A2(n1813), .B(n547), .ZN(n1082) );
  MUX2NUD1BWP30P140LVT U1070 ( .I0(n1191), .I1(n1748), .S(copy_pointer[0]), 
        .ZN(n1147) );
  AOI21D1BWP30P140LVT U1071 ( .A1(n9), .A2(n549), .B(n548), .ZN(N3861) );
  INR2D1BWP30P140LVT U1072 ( .A1(n634), .B1(n1191), .ZN(n618) );
  AO21D1BWP30P140LVT U1073 ( .A1(n1245), .A2(pointer[0]), .B(n618), .Z(n1179)
         );
  INVD1BWP30P140LVT U1074 ( .I(n550), .ZN(n552) );
  FA1D1BWP30P140LVT U1075 ( .A(hardware_latency2[1]), .B(hardware_latency1[1]), 
        .CI(n1665), .CO(n554), .S(n544) );
  INVD1BWP30P140LVT U1076 ( .I(n656), .ZN(n556) );
  ND2OPTIBD1BWP30P140LVT U1077 ( .A1(n555), .A2(n554), .ZN(n658) );
  XOR2UD1BWP30P140LVT U1078 ( .A1(n640), .A2(n557), .Z(n1978) );
  AOI21D1BWP30P140LVT U1079 ( .A1(n1813), .A2(delay_matrix_N_1_next[44]), .B(
        n1807), .ZN(n558) );
  OAI21D1BWP30P140LVT U1080 ( .A1(n1211), .A2(n1813), .B(n558), .ZN(n1081) );
  INR2D1BWP30P140LVT U1081 ( .A1(copy_pointer[0]), .B1(n559), .ZN(n560) );
  ND2OPTIBD2BWP30P140LVT U1082 ( .A1(n560), .A2(n4), .ZN(n1806) );
  OAI21D1BWP30P140LVT U1083 ( .A1(n560), .A2(n1191), .B(n1748), .ZN(n1801) );
  AOI21D1BWP30P140LVT U1084 ( .A1(n1773), .A2(
        delay_matrix_N_1_next_original[51]), .B(n1280), .ZN(n562) );
  OAI211D1BWP30P140LVT U1085 ( .A1(n1806), .A2(n1282), .B(n563), .C(n562), 
        .ZN(n816) );
  INVD2BWP30P140LVT U1086 ( .I(delay_matrix_element[8]), .ZN(n1776) );
  INR2D1BWP30P140LVT U1087 ( .A1(n574), .B1(copy_pointer[0]), .ZN(n565) );
  OAI21D1BWP30P140LVT U1088 ( .A1(n565), .A2(n2172), .B(n1748), .ZN(n2194) );
  AOI21D1BWP30P140LVT U1089 ( .A1(scenario_update), .A2(
        delay_matrix_N_1_next_original[8]), .B(n1280), .ZN(n566) );
  OAI211D1BWP30P140LVT U1090 ( .A1(n1776), .A2(n2196), .B(n567), .C(n566), 
        .ZN(n859) );
  AOI21D1BWP30P140LVT U1091 ( .A1(n1773), .A2(
        delay_matrix_N_1_next_original[9]), .B(n1280), .ZN(n568) );
  OAI211D1BWP30P140LVT U1092 ( .A1(n1282), .A2(n2196), .B(n569), .C(n568), 
        .ZN(n858) );
  INVD2BWP30P140LVT U1093 ( .I(delay_matrix_element[10]), .ZN(n2206) );
  AOI21D1BWP30P140LVT U1094 ( .A1(n1773), .A2(
        delay_matrix_N_1_next_original[52]), .B(n1280), .ZN(n570) );
  OAI211D1BWP30P140LVT U1095 ( .A1(n2206), .A2(n1806), .B(n571), .C(n570), 
        .ZN(n815) );
  INVD2BWP30P140LVT U1096 ( .I(delay_matrix_element[11]), .ZN(n1465) );
  AOI21D1BWP30P140LVT U1097 ( .A1(n1773), .A2(
        delay_matrix_N_1_next_original[53]), .B(n1280), .ZN(n572) );
  OAI211D1BWP30P140LVT U1098 ( .A1(n1465), .A2(n1806), .B(n573), .C(n572), 
        .ZN(n814) );
  ND2OPTIBD2BWP30P140LVT U1099 ( .A1(n575), .A2(n4), .ZN(n2202) );
  OAI21D1BWP30P140LVT U1100 ( .A1(n575), .A2(n2172), .B(n1748), .ZN(n2200) );
  AOI21D1BWP30P140LVT U1101 ( .A1(n1773), .A2(
        delay_matrix_N_1_next_original[23]), .B(n1280), .ZN(n576) );
  OAI211D1BWP30P140LVT U1102 ( .A1(n2202), .A2(n1282), .B(n577), .C(n576), 
        .ZN(n844) );
  AOI22D1BWP30P140LVT U1103 ( .A1(delay_matrix_N_1_original[25]), .A2(n2200), 
        .B1(n561), .B2(delay_matrix_N_1_next_original[25]), .ZN(n578) );
  OAI211D1BWP30P140LVT U1104 ( .A1(n2202), .A2(n1465), .B(n578), .C(n1821), 
        .ZN(n842) );
  AOI21D1BWP30P140LVT U1105 ( .A1(n1773), .A2(
        delay_matrix_N_1_next_original[37]), .B(n1280), .ZN(n579) );
  OAI211D1BWP30P140LVT U1106 ( .A1(n2207), .A2(n1282), .B(n580), .C(n579), 
        .ZN(n830) );
  NR4D0BWP30P140LVT U1107 ( .A1(copy_ptr_next[22]), .A2(copy_ptr_next[20]), 
        .A3(copy_ptr_next[24]), .A4(copy_ptr_next[18]), .ZN(n584) );
  NR4D0BWP30P140LVT U1108 ( .A1(copy_ptr_next[23]), .A2(copy_ptr_next[19]), 
        .A3(copy_ptr_next[21]), .A4(copy_ptr_next[17]), .ZN(n583) );
  NR4D0BWP30P140LVT U1109 ( .A1(copy_ptr_next[15]), .A2(copy_ptr_next[11]), 
        .A3(copy_ptr_next[13]), .A4(copy_ptr_next[9]), .ZN(n582) );
  NR4D0BWP30P140LVT U1110 ( .A1(copy_ptr_next[25]), .A2(copy_ptr_next[8]), 
        .A3(copy_ptr_next[6]), .A4(copy_ptr_next[2]), .ZN(n581) );
  ND4D1BWP30P140LVT U1111 ( .A1(n584), .A2(n583), .A3(n582), .A4(n581), .ZN(
        n591) );
  NR4D0BWP30P140LVT U1112 ( .A1(copy_ptr_next[14]), .A2(copy_ptr_next[12]), 
        .A3(copy_ptr_next[10]), .A4(copy_ptr_next[4]), .ZN(n586) );
  NR4D0BWP30P140LVT U1113 ( .A1(copy_ptr_next[16]), .A2(copy_ptr_next[7]), 
        .A3(copy_ptr_next[5]), .A4(copy_ptr_next[3]), .ZN(n585) );
  NR4D0BWP30P140LVT U1114 ( .A1(copy_ptr_next[30]), .A2(copy_ptr_next[29]), 
        .A3(copy_ptr_next[28]), .A4(copy_ptr_next[27]), .ZN(n588) );
  ND3D1BWP30P140LVT U1115 ( .A1(n588), .A2(glob_scen_noc_input_valid), .A3(
        n587), .ZN(n589) );
  NR3D0P7BWP30P140LVT U1116 ( .A1(n591), .A2(n590), .A3(n589), .ZN(n1197) );
  INR2D1BWP30P140LVT U1117 ( .A1(copy_ptr_next[0]), .B1(copy_ptr_next[1]), 
        .ZN(n592) );
  AOI21D1BWP30P140LVT U1118 ( .A1(n1392), .A2(
        delay_matrix_N_1_next_original[23]), .B(n1280), .ZN(n593) );
  OAI21D1BWP30P140LVT U1119 ( .A1(n1282), .A2(n1392), .B(n593), .ZN(n872) );
  INR2D1BWP30P140LVT U1120 ( .A1(copy_ptr_next[1]), .B1(copy_ptr_next[0]), 
        .ZN(n594) );
  AOI21D1BWP30P140LVT U1121 ( .A1(n1398), .A2(
        delay_matrix_N_1_next_original[37]), .B(n1280), .ZN(n595) );
  OAI21D1BWP30P140LVT U1122 ( .A1(n1282), .A2(n1398), .B(n595), .ZN(n900) );
  AOI21D1BWP30P140LVT U1123 ( .A1(n1404), .A2(
        delay_matrix_N_1_next_original[8]), .B(n1280), .ZN(n597) );
  OAI21D1BWP30P140LVT U1124 ( .A1(n1776), .A2(n1404), .B(n597), .ZN(n887) );
  AOI21D1BWP30P140LVT U1125 ( .A1(n1404), .A2(
        delay_matrix_N_1_next_original[9]), .B(n1280), .ZN(n598) );
  OAI21D1BWP30P140LVT U1126 ( .A1(n1282), .A2(n1404), .B(n598), .ZN(n886) );
  NR4D0BWP30P140LVT U1127 ( .A1(pointer[2]), .A2(pointer[6]), .A3(pointer[8]), 
        .A4(pointer[18]), .ZN(n602) );
  NR4D0BWP30P140LVT U1128 ( .A1(pointer[5]), .A2(pointer[7]), .A3(pointer[9]), 
        .A4(pointer[11]), .ZN(n601) );
  NR4D0BWP30P140LVT U1129 ( .A1(pointer[20]), .A2(pointer[22]), .A3(pointer[3]), .A4(pointer[24]), .ZN(n600) );
  NR2D1BWP30P140LVT U1130 ( .A1(pointer[31]), .A2(pointer[30]), .ZN(n599) );
  ND4D1BWP30P140LVT U1131 ( .A1(n602), .A2(n601), .A3(n600), .A4(n599), .ZN(
        n609) );
  NR4D0BWP30P140LVT U1132 ( .A1(pointer[13]), .A2(pointer[15]), .A3(
        pointer[17]), .A4(pointer[19]), .ZN(n604) );
  NR4D0BWP30P140LVT U1133 ( .A1(pointer[21]), .A2(pointer[23]), .A3(pointer[4]), .A4(pointer[25]), .ZN(n603) );
  NR4D0BWP30P140LVT U1134 ( .A1(pointer[26]), .A2(pointer[27]), .A3(
        pointer[28]), .A4(pointer[29]), .ZN(n606) );
  NR4D0BWP30P140LVT U1135 ( .A1(pointer[10]), .A2(pointer[12]), .A3(
        pointer[14]), .A4(pointer[16]), .ZN(n605) );
  NR3D0P7BWP30P140LVT U1136 ( .A1(n609), .A2(n608), .A3(n607), .ZN(n699) );
  AOI21D1BWP30P140LVT U1137 ( .A1(n561), .A2(delay_matrix_N_1_next[28]), .B(
        n1807), .ZN(n615) );
  INVD1BWP30P140LVT U1138 ( .I(n611), .ZN(n612) );
  OAI211D1BWP30P140LVT U1139 ( .A1(n1646), .A2(n2191), .B(n615), .C(n614), 
        .ZN(n991) );
  AOI21D1BWP30P140LVT U1140 ( .A1(n1773), .A2(
        delay_matrix_N_1_next_original[39]), .B(n1280), .ZN(n616) );
  OAI211D1BWP30P140LVT U1141 ( .A1(n1465), .A2(n2207), .B(n617), .C(n616), 
        .ZN(n828) );
  AOI21D1BWP30P140LVT U1142 ( .A1(n561), .A2(delay_matrix_N_1_next[2]), .B(
        n1807), .ZN(n621) );
  OAI21D1BWP30P140LVT U1143 ( .A1(n2172), .A2(n634), .B(n633), .ZN(n2179) );
  OAI211D1BWP30P140LVT U1144 ( .A1(n1211), .A2(n2181), .B(n621), .C(n620), 
        .ZN(n1017) );
  OAI211D1BWP30P140LVT U1145 ( .A1(n2199), .A2(n1404), .B(n622), .C(n1821), 
        .ZN(n883) );
  OAI211D1BWP30P140LVT U1146 ( .A1(n2203), .A2(n1404), .B(n623), .C(n1821), 
        .ZN(n882) );
  OAI211D1BWP30P140LVT U1147 ( .A1(n2199), .A2(n1392), .B(n624), .C(n1821), 
        .ZN(n869) );
  OAI211D1BWP30P140LVT U1148 ( .A1(n2203), .A2(n1398), .B(n625), .C(n1821), 
        .ZN(n896) );
  OAI211D1BWP30P140LVT U1149 ( .A1(n2203), .A2(n1392), .B(n626), .C(n1821), 
        .ZN(n868) );
  OAI211D1BWP30P140LVT U1150 ( .A1(n2199), .A2(n1398), .B(n627), .C(n1821), 
        .ZN(n897) );
  INVD1BWP30P140LVT U1151 ( .I(obj_id_next[6]), .ZN(n745) );
  OAI22D1BWP30P140LVT U1152 ( .A1(n778), .A2(n745), .B1(n779), .B2(n1208), 
        .ZN(n1055) );
  INVD1BWP30P140LVT U1153 ( .I(obj_id_next[7]), .ZN(n747) );
  OAI22D1BWP30P140LVT U1154 ( .A1(n778), .A2(n747), .B1(n779), .B2(n1206), 
        .ZN(n1054) );
  NR3D0P7BWP30P140LVT U1155 ( .A1(n1204), .A2(ptr_next[0]), .A3(ptr_next[1]), 
        .ZN(n630) );
  INVD1BWP30P140LVT U1156 ( .I(obj_id_next[0]), .ZN(n631) );
  OAI22D1BWP30P140LVT U1157 ( .A1(n776), .A2(n631), .B1(n777), .B2(n1208), 
        .ZN(n1051) );
  INVD1BWP30P140LVT U1158 ( .I(obj_id_next[1]), .ZN(n632) );
  OAI22D1BWP30P140LVT U1159 ( .A1(n776), .A2(n632), .B1(n777), .B2(n1206), 
        .ZN(n1050) );
  OAI21D1BWP30P140LVT U1160 ( .A1(pointer[0]), .A2(n2172), .B(n633), .ZN(n2183) );
  NR2D1BWP30P140LVT U1161 ( .A1(n1646), .A2(n2185), .ZN(n637) );
  AOI211D1BWP30P140LVT U1162 ( .A1(n1773), .A2(delay_matrix_N_1_next[14]), .B(
        n637), .C(n1280), .ZN(n638) );
  OAI21D1BWP30P140LVT U1163 ( .A1(n1933), .A2(n639), .B(n638), .ZN(n1005) );
  OAI21D1BWP30P140LVT U1164 ( .A1(n640), .A2(n656), .B(n658), .ZN(n646) );
  FA1D1BWP30P140LVT U1165 ( .A(hardware_latency2[2]), .B(hardware_latency1[2]), 
        .CI(n641), .CO(n642), .S(n555) );
  INVD1BWP30P140LVT U1166 ( .I(n659), .ZN(n644) );
  AOI21D1BWP30P140LVT U1167 ( .A1(n1813), .A2(delay_matrix_N_1_next[45]), .B(
        n1807), .ZN(n647) );
  OAI21D1BWP30P140LVT U1168 ( .A1(n1215), .A2(n1813), .B(n647), .ZN(n1080) );
  INVD1BWP30P140LVT U1169 ( .I(n1806), .ZN(n649) );
  AOI22D1BWP30P140LVT U1170 ( .A1(n649), .A2(delay_matrix_element[12]), .B1(
        n561), .B2(delay_matrix_N_1_next_original[54]), .ZN(n648) );
  IOA21D1BWP30P140LVT U1171 ( .A1(delay_matrix_N_1_original[54]), .A2(n1801), 
        .B(n648), .ZN(n813) );
  AOI22D1BWP30P140LVT U1172 ( .A1(n649), .A2(delay_matrix_element[13]), .B1(
        n561), .B2(delay_matrix_N_1_next_original[55]), .ZN(n650) );
  IOA21D1BWP30P140LVT U1173 ( .A1(delay_matrix_N_1_original[55]), .A2(n1801), 
        .B(n650), .ZN(n812) );
  AOI21D1BWP30P140LVT U1174 ( .A1(n561), .A2(delay_matrix_N_1_next[3]), .B(
        n1807), .ZN(n652) );
  OAI211D1BWP30P140LVT U1175 ( .A1(n1215), .A2(n2181), .B(n652), .C(n651), 
        .ZN(n1016) );
  AOI21D1BWP30P140LVT U1176 ( .A1(n1815), .A2(delay_matrix_N_1_next[2]), .B(
        n1807), .ZN(n653) );
  OAI21D1BWP30P140LVT U1177 ( .A1(n1211), .A2(n1815), .B(n653), .ZN(n1045) );
  AOI21D1BWP30P140LVT U1178 ( .A1(n1815), .A2(delay_matrix_N_1_next[1]), .B(
        n1807), .ZN(n654) );
  OAI21D1BWP30P140LVT U1179 ( .A1(n1627), .A2(n1815), .B(n654), .ZN(n1046) );
  AOI21D1BWP30P140LVT U1180 ( .A1(n1815), .A2(delay_matrix_N_1_next[3]), .B(
        n1807), .ZN(n655) );
  OAI21D1BWP30P140LVT U1181 ( .A1(n1215), .A2(n1815), .B(n655), .ZN(n1044) );
  OAI21D1BWP30P140LVT U1182 ( .A1(n659), .A2(n658), .B(n657), .ZN(n660) );
  AOI21D2BWP30P140LVT U1183 ( .A1(n662), .A2(n661), .B(n660), .ZN(n691) );
  INVD2BWP30P140LVT U1184 ( .I(n691), .ZN(n1553) );
  FA1D1BWP30P140LVT U1185 ( .A(hardware_latency2[3]), .B(hardware_latency1[3]), 
        .CI(n663), .CO(n664), .S(n643) );
  INVD1BWP30P140LVT U1186 ( .I(n680), .ZN(n1552) );
  AOI21D1BWP30P140LVT U1187 ( .A1(n1813), .A2(delay_matrix_N_1_next[46]), .B(
        n1807), .ZN(n667) );
  OAI21D1BWP30P140LVT U1188 ( .A1(n1254), .A2(n1813), .B(n667), .ZN(n1079) );
  AOI21D1BWP30P140LVT U1189 ( .A1(n1815), .A2(delay_matrix_N_1_next[4]), .B(
        n1807), .ZN(n668) );
  OAI21D1BWP30P140LVT U1190 ( .A1(n1254), .A2(n1815), .B(n668), .ZN(n1043) );
  OAI211D1BWP30P140LVT U1191 ( .A1(n1404), .A2(n2206), .B(n669), .C(n1821), 
        .ZN(n885) );
  OAI211D1BWP30P140LVT U1192 ( .A1(n1398), .A2(n1465), .B(n670), .C(n1821), 
        .ZN(n898) );
  OAI211D1BWP30P140LVT U1193 ( .A1(n1404), .A2(n1465), .B(n671), .C(n1821), 
        .ZN(n884) );
  OAI211D1BWP30P140LVT U1194 ( .A1(n1392), .A2(n1465), .B(n672), .C(n1821), 
        .ZN(n870) );
  OAI211D1BWP30P140LVT U1195 ( .A1(n1392), .A2(n2206), .B(n673), .C(n1821), 
        .ZN(n871) );
  OAI211D1BWP30P140LVT U1196 ( .A1(n1398), .A2(n2206), .B(n674), .C(n1821), 
        .ZN(n899) );
  INVD1BWP30P140LVT U1197 ( .I(n2200), .ZN(n1766) );
  AOI21D1BWP30P140LVT U1198 ( .A1(n1773), .A2(
        delay_matrix_N_1_next_original[22]), .B(n1280), .ZN(n676) );
  INVD1BWP30P140LVT U1199 ( .I(n2202), .ZN(n1762) );
  OAI211D1BWP30P140LVT U1200 ( .A1(n1766), .A2(n677), .B(n676), .C(n675), .ZN(
        n845) );
  AOI21D1BWP30P140LVT U1201 ( .A1(n561), .A2(delay_matrix_N_1_next[4]), .B(
        n1807), .ZN(n679) );
  OAI211D1BWP30P140LVT U1202 ( .A1(n1254), .A2(n2181), .B(n679), .C(n678), 
        .ZN(n1015) );
  INVD1BWP30P140LVT U1203 ( .I(delay_matrix_N_1[22]), .ZN(n698) );
  FA1D1BWP30P140LVT U1204 ( .A(hardware_latency2[4]), .B(hardware_latency1[4]), 
        .CI(n1790), .CO(n681), .S(n665) );
  FA1D1BWP30P140LVT U1205 ( .A(hardware_latency2[5]), .B(hardware_latency1[5]), 
        .CI(n1798), .CO(n683), .S(n682) );
  FA1D1BWP30P140LVT U1206 ( .A(hardware_latency2[6]), .B(hardware_latency1[6]), 
        .CI(n1805), .CO(n685), .S(n684) );
  ND2OPTIBD1BWP30P140LVT U1207 ( .A1(n682), .A2(n681), .ZN(n1555) );
  OAI21D1BWP30P140LVT U1208 ( .A1(n1554), .A2(n1550), .B(n1555), .ZN(n706) );
  ND2OPTIBD1BWP30P140LVT U1209 ( .A1(n686), .A2(n685), .ZN(n1312) );
  OAI21D1BWP30P140LVT U1210 ( .A1(n1311), .A2(n1308), .B(n1312), .ZN(n687) );
  AOI21D1BWP30P140LVT U1211 ( .A1(n688), .A2(n706), .B(n687), .ZN(n689) );
  OAI21OPTREPBD2BWP30P140LVT U1212 ( .A1(n691), .A2(n690), .B(n689), .ZN(n1232) );
  INVD2BWP30P140LVT U1213 ( .I(n1232), .ZN(n1407) );
  FA1D1BWP30P140LVT U1214 ( .A(hardware_latency2[7]), .B(hardware_latency1[7]), 
        .CI(n1779), .CO(n692), .S(n686) );
  INVD1BWP30P140LVT U1215 ( .I(n1406), .ZN(n694) );
  XOR2UD1BWP30P140LVT U1216 ( .A1(n1407), .A2(n695), .Z(n1949) );
  AOI21D1BWP30P140LVT U1217 ( .A1(n561), .A2(delay_matrix_N_1_next[22]), .B(
        n1807), .ZN(n696) );
  OAI211D1BWP30P140LVT U1218 ( .A1(n1933), .A2(n698), .B(n697), .C(n696), .ZN(
        n997) );
  ND3D1BWP30P140LVT U1219 ( .A1(n699), .A2(pointer[0]), .A3(pointer[1]), .ZN(
        n701) );
  NR2D1BWP30P140LVT U1220 ( .A1(n1988), .A2(n702), .ZN(n703) );
  AOI211D1BWP30P140LVT U1221 ( .A1(n1773), .A2(delay_matrix_N_1_next[42]), .B(
        n703), .C(n1280), .ZN(n704) );
  OAI21D1BWP30P140LVT U1222 ( .A1(n1646), .A2(n1461), .B(n704), .ZN(n977) );
  AOI22D1BWP30P140LVT U1223 ( .A1(delay_matrix_N_1_original[11]), .A2(n2194), 
        .B1(n1802), .B2(delay_matrix_N_1_next_original[11]), .ZN(n705) );
  OAI211D1BWP30P140LVT U1224 ( .A1(n2196), .A2(n1465), .B(n705), .C(n1821), 
        .ZN(n856) );
  INVD1BWP30P140LVT U1225 ( .I(n1309), .ZN(n708) );
  XOR2UD1BWP30P140LVT U1226 ( .A1(n1310), .A2(n709), .Z(n1962) );
  AOI21D1BWP30P140LVT U1227 ( .A1(n561), .A2(delay_matrix_N_1_next[20]), .B(
        n1807), .ZN(n710) );
  OAI211D1BWP30P140LVT U1228 ( .A1(n1933), .A2(n712), .B(n711), .C(n710), .ZN(
        n999) );
  AOI21D1BWP30P140LVT U1229 ( .A1(n561), .A2(delay_matrix_N_1_next[50]), .B(
        n1807), .ZN(n713) );
  OAI211D1BWP30P140LVT U1230 ( .A1(n1988), .A2(n715), .B(n714), .C(n713), .ZN(
        n969) );
  MUX2NUD1BWP30P140LVT U1231 ( .I0(n13), .I1(n1835), .S(copy_ptr_next[0]), 
        .ZN(n955) );
  MUX2NUD1BWP30P140LVT U1232 ( .I0(n13), .I1(n1835), .S(ptr_next[0]), .ZN(
        n1115) );
  INVD1BWP30P140LVT U1233 ( .I(n717), .ZN(n718) );
  ND2D1BWP30P140LVT U1234 ( .A1(n1260), .A2(n718), .ZN(n731) );
  INVD1BWP30P140LVT U1235 ( .I(copy_ptr_next[10]), .ZN(n730) );
  NR2D1BWP30P140LVT U1236 ( .A1(n731), .A2(n730), .ZN(n720) );
  INVD1BWP30P140LVT U1237 ( .I(copy_ptr_next[11]), .ZN(n719) );
  XNR2UD1BWP30P140LVT U1238 ( .A1(n720), .A2(n719), .ZN(n721) );
  MOAI22D1BWP30P140LVT U1239 ( .A1(n1835), .A2(n719), .B1(n6), .B2(n721), .ZN(
        n944) );
  INVD1BWP30P140LVT U1240 ( .I(copy_ptr_next[9]), .ZN(n722) );
  XOR2UD1BWP30P140LVT U1241 ( .A1(n723), .A2(n722), .Z(n724) );
  MOAI22D1BWP30P140LVT U1242 ( .A1(n1835), .A2(n722), .B1(n6), .B2(n724), .ZN(
        n946) );
  INVD1BWP30P140LVT U1243 ( .I(n738), .ZN(n735) );
  INVD1BWP30P140LVT U1244 ( .I(copy_ptr_next[12]), .ZN(n737) );
  XNR2UD1BWP30P140LVT U1245 ( .A1(n735), .A2(n737), .ZN(n726) );
  MOAI22D1BWP30P140LVT U1246 ( .A1(n1835), .A2(n737), .B1(n6), .B2(n726), .ZN(
        n943) );
  INVD1BWP30P140LVT U1247 ( .I(n727), .ZN(n1262) );
  INVD1BWP30P140LVT U1248 ( .I(copy_ptr_next[2]), .ZN(n728) );
  XNR2UD1BWP30P140LVT U1249 ( .A1(n1262), .A2(n728), .ZN(n729) );
  MOAI22D1BWP30P140LVT U1250 ( .A1(n1835), .A2(n728), .B1(n6), .B2(n729), .ZN(
        n953) );
  XOR2UD1BWP30P140LVT U1251 ( .A1(n731), .A2(n730), .Z(n732) );
  MOAI22D1BWP30P140LVT U1252 ( .A1(n1835), .A2(n730), .B1(n6), .B2(n732), .ZN(
        n945) );
  INVD1BWP30P140LVT U1253 ( .I(n733), .ZN(n734) );
  ND2D1BWP30P140LVT U1254 ( .A1(n735), .A2(n734), .ZN(n1885) );
  INVD1BWP30P140LVT U1255 ( .I(copy_ptr_next[14]), .ZN(n1884) );
  XOR2UD1BWP30P140LVT U1256 ( .A1(n1885), .A2(n1884), .Z(n736) );
  MOAI22D1BWP30P140LVT U1257 ( .A1(n1835), .A2(n1884), .B1(n6), .B2(n736), 
        .ZN(n941) );
  NR2D1BWP30P140LVT U1258 ( .A1(n738), .A2(n737), .ZN(n740) );
  INVD1BWP30P140LVT U1259 ( .I(copy_ptr_next[13]), .ZN(n739) );
  XNR2UD1BWP30P140LVT U1260 ( .A1(n740), .A2(n739), .ZN(n741) );
  MOAI22D1BWP30P140LVT U1261 ( .A1(n1835), .A2(n739), .B1(n6), .B2(n741), .ZN(
        n942) );
  INVD1BWP30P140LVT U1262 ( .I(copy_ptr_next[16]), .ZN(n1889) );
  XOR2UD1BWP30P140LVT U1263 ( .A1(n1890), .A2(n1889), .Z(n743) );
  MOAI22D1BWP30P140LVT U1264 ( .A1(n1835), .A2(n1889), .B1(n6), .B2(n743), 
        .ZN(n939) );
  INVD1BWP30P140LVT U1265 ( .I(obj_id_element[0]), .ZN(n2187) );
  OAI222D1BWP30P140LVT U1266 ( .A1(n5), .A2(n745), .B1(n744), .B2(n1988), .C1(
        n1461), .C2(n2187), .ZN(n957) );
  INVD1BWP30P140LVT U1267 ( .I(obj_id_element[1]), .ZN(n2190) );
  OAI222D1BWP30P140LVT U1268 ( .A1(n5), .A2(n747), .B1(n746), .B2(n1988), .C1(
        n1461), .C2(n2190), .ZN(n956) );
  FA1D1BWP30P140LVT U1269 ( .A(hardware_latency2[8]), .B(hardware_latency1[8]), 
        .CI(n1776), .CO(n749), .S(n693) );
  FA1D1BWP30P140LVT U1270 ( .A(hardware_latency2[9]), .B(hardware_latency1[9]), 
        .CI(n748), .CO(n751), .S(n750) );
  FA1D1BWP30P140LVT U1271 ( .A(hardware_latency2[10]), .B(
        hardware_latency1[10]), .CI(n2206), .CO(n753), .S(n752) );
  INVD1BWP30P140LVT U1272 ( .I(n764), .ZN(n758) );
  OAI21D1BWP30P140LVT U1273 ( .A1(n1408), .A2(n1405), .B(n1409), .ZN(n1230) );
  OAI21D1BWP30P140LVT U1274 ( .A1(n1269), .A2(n1266), .B(n1270), .ZN(n755) );
  AOI21D1BWP30P140LVT U1275 ( .A1(n756), .A2(n1230), .B(n755), .ZN(n767) );
  AOI21D1BWP30P140LVT U1276 ( .A1(n1232), .A2(n758), .B(n757), .ZN(n763) );
  FA1D1BWP30P140LVT U1277 ( .A(hardware_latency2[11]), .B(
        hardware_latency1[11]), .CI(n1465), .CO(n759), .S(n754) );
  INVD1BWP30P140LVT U1278 ( .I(n766), .ZN(n761) );
  XOR2UD1BWP30P140LVT U1279 ( .A1(n763), .A2(n762), .Z(n1219) );
  INVD1BWP30P140LVT U1280 ( .I(delay_matrix_N_1_next[12]), .ZN(n1220) );
  OAI22D1BWP30P140LVT U1281 ( .A1(n1229), .A2(n777), .B1(n776), .B2(n1220), 
        .ZN(n1035) );
  INVD1BWP30P140LVT U1282 ( .I(delay_matrix_N_1_next[54]), .ZN(n1304) );
  OAI22D1BWP30P140LVT U1283 ( .A1(n1229), .A2(n779), .B1(n778), .B2(n1304), 
        .ZN(n1071) );
  NR2D1BWP30P140LVT U1284 ( .A1(n764), .A2(n766), .ZN(n769) );
  OAI21D1BWP30P140LVT U1285 ( .A1(n767), .A2(n766), .B(n765), .ZN(n768) );
  AOI21D1BWP30P140LVT U1286 ( .A1(n1232), .A2(n769), .B(n768), .ZN(n775) );
  FA1D1BWP30P140LVT U1287 ( .A(hardware_latency2[12]), .B(
        hardware_latency1[12]), .CI(n2199), .CO(n770), .S(n760) );
  OR2D1BWP30P140LVT U1288 ( .A1(n771), .A2(n770), .Z(n773) );
  XOR2UD1BWP30P140LVT U1289 ( .A1(n775), .A2(n774), .Z(n1241) );
  INVD1BWP30P140LVT U1290 ( .I(delay_matrix_N_1_next[13]), .ZN(n1247) );
  OAI22D1BWP30P140LVT U1291 ( .A1(n1225), .A2(n777), .B1(n776), .B2(n1247), 
        .ZN(n1034) );
  INVD1BWP30P140LVT U1292 ( .I(delay_matrix_N_1_next[55]), .ZN(n1463) );
  OAI22D1BWP30P140LVT U1293 ( .A1(n1225), .A2(n779), .B1(n778), .B2(n1463), 
        .ZN(n1070) );
  NR3D0P7BWP30P140LVT U1294 ( .A1(n1204), .A2(ptr_next[0]), .A3(n1824), .ZN(
        n780) );
  INVD1BWP30P140LVT U1295 ( .I(obj_id_next[4]), .ZN(n781) );
  OAI22D1BWP30P140LVT U1296 ( .A1(n1223), .A2(n781), .B1(n1224), .B2(n1208), 
        .ZN(n1053) );
  INVD1BWP30P140LVT U1297 ( .I(obj_id_next[5]), .ZN(n809) );
  OAI22D1BWP30P140LVT U1298 ( .A1(n1223), .A2(n809), .B1(n1224), .B2(n1206), 
        .ZN(n1052) );
  AOI21D1BWP30P140LVT U1299 ( .A1(n1817), .A2(delay_matrix_N_1_next[31]), .B(
        n1807), .ZN(n1180) );
  OAI21D1BWP30P140LVT U1300 ( .A1(n1215), .A2(n1817), .B(n1180), .ZN(n1066) );
  AOI21D1BWP30P140LVT U1301 ( .A1(n1817), .A2(delay_matrix_N_1_next[30]), .B(
        n1807), .ZN(n1181) );
  OAI21D1BWP30P140LVT U1302 ( .A1(n1211), .A2(n1817), .B(n1181), .ZN(n1067) );
  AOI21D1BWP30P140LVT U1303 ( .A1(n1817), .A2(delay_matrix_N_1_next[29]), .B(
        n1807), .ZN(n1182) );
  OAI21D1BWP30P140LVT U1304 ( .A1(n1627), .A2(n1817), .B(n1182), .ZN(n1068) );
  AOI21D1BWP30P140LVT U1305 ( .A1(n1817), .A2(delay_matrix_N_1_next[28]), .B(
        n1807), .ZN(n1183) );
  OAI21D1BWP30P140LVT U1306 ( .A1(n1646), .A2(n1817), .B(n1183), .ZN(n1069) );
  INVD1BWP30P140LVT U1307 ( .I(n1201), .ZN(n1190) );
  ND2D1BWP30P140LVT U1308 ( .A1(n1190), .A2(copy_pointer[2]), .ZN(n1185) );
  INVD1BWP30P140LVT U1309 ( .I(copy_pointer[3]), .ZN(n1184) );
  XOR2UD1BWP30P140LVT U1310 ( .A1(n1185), .A2(n1184), .Z(n1186) );
  MOAI22D1BWP30P140LVT U1311 ( .A1(n1184), .A2(n1748), .B1(n1186), .B2(n4), 
        .ZN(n1144) );
  INVD1BWP30P140LVT U1312 ( .I(pointer[2]), .ZN(n1189) );
  INVD1BWP30P140LVT U1313 ( .I(n1187), .ZN(n1193) );
  XNR2UD1BWP30P140LVT U1314 ( .A1(n1193), .A2(n1189), .ZN(n1188) );
  MOAI22D1BWP30P140LVT U1315 ( .A1(n1189), .A2(n1748), .B1(n1188), .B2(n4), 
        .ZN(n1177) );
  XNR2UD1BWP30P140LVT U1316 ( .A1(n1190), .A2(n2208), .ZN(n1192) );
  MOAI22D1BWP30P140LVT U1317 ( .A1(n2208), .A2(n1748), .B1(n1192), .B2(n4), 
        .ZN(n1145) );
  INVD1BWP30P140LVT U1318 ( .I(pointer[3]), .ZN(n1196) );
  ND2D1BWP30P140LVT U1319 ( .A1(n1193), .A2(pointer[2]), .ZN(n1194) );
  XOR2UD1BWP30P140LVT U1320 ( .A1(n1194), .A2(n1196), .Z(n1195) );
  MOAI22D1BWP30P140LVT U1321 ( .A1(n1196), .A2(n1748), .B1(n1195), .B2(n4), 
        .ZN(n1176) );
  ND3D1BWP30P140LVT U1322 ( .A1(n1197), .A2(copy_ptr_next[1]), .A3(
        copy_ptr_next[0]), .ZN(n1333) );
  OAI211D1BWP30P140LVT U1323 ( .A1(n2206), .A2(n1333), .B(n1198), .C(n1821), 
        .ZN(n913) );
  INVD1BWP30P140LVT U1324 ( .I(pointer[1]), .ZN(n1200) );
  XNR2UD1BWP30P140LVT U1325 ( .A1(n1200), .A2(pointer[0]), .ZN(n1199) );
  MOAI22D1BWP30P140LVT U1326 ( .A1(n1200), .A2(n1748), .B1(n1199), .B2(n4), 
        .ZN(n1178) );
  INVD1BWP30P140LVT U1327 ( .I(n1489), .ZN(n1593) );
  INVD1BWP30P140LVT U1328 ( .I(copy_pointer[4]), .ZN(n1592) );
  XOR2UD1BWP30P140LVT U1329 ( .A1(n1593), .A2(n1592), .Z(n1203) );
  MOAI22D1BWP30P140LVT U1330 ( .A1(n1592), .A2(n1748), .B1(n4), .B2(n1203), 
        .ZN(n1143) );
  INR3D0BWP30P140LVT U1331 ( .A1(ptr_next[0]), .B1(ptr_next[1]), .B2(n1204), 
        .ZN(n1205) );
  INVD1BWP30P140LVT U1332 ( .I(obj_id_next[3]), .ZN(n1207) );
  OAI22D1BWP30P140LVT U1333 ( .A1(n1227), .A2(n1207), .B1(n1228), .B2(n1206), 
        .ZN(n1048) );
  INVD1BWP30P140LVT U1334 ( .I(obj_id_next[2]), .ZN(n1209) );
  OAI22D1BWP30P140LVT U1335 ( .A1(n1227), .A2(n1209), .B1(n1228), .B2(n1208), 
        .ZN(n1049) );
  AOI21D1BWP30P140LVT U1336 ( .A1(n1819), .A2(delay_matrix_N_1_next[16]), .B(
        n1807), .ZN(n1210) );
  OAI21D1BWP30P140LVT U1337 ( .A1(n1211), .A2(n1819), .B(n1210), .ZN(n1031) );
  AOI21D1BWP30P140LVT U1338 ( .A1(n1819), .A2(delay_matrix_N_1_next[14]), .B(
        n1807), .ZN(n1212) );
  OAI21D1BWP30P140LVT U1339 ( .A1(n1646), .A2(n1819), .B(n1212), .ZN(n1033) );
  AOI21D1BWP30P140LVT U1340 ( .A1(n1819), .A2(delay_matrix_N_1_next[18]), .B(
        n1807), .ZN(n1213) );
  OAI21D1BWP30P140LVT U1341 ( .A1(n1254), .A2(n1819), .B(n1213), .ZN(n1029) );
  AOI21D1BWP30P140LVT U1342 ( .A1(n1819), .A2(delay_matrix_N_1_next[17]), .B(
        n1807), .ZN(n1214) );
  OAI21D1BWP30P140LVT U1343 ( .A1(n1215), .A2(n1819), .B(n1214), .ZN(n1030) );
  AOI21D1BWP30P140LVT U1344 ( .A1(n1819), .A2(delay_matrix_N_1_next[15]), .B(
        n1807), .ZN(n1216) );
  OAI21D1BWP30P140LVT U1345 ( .A1(n1627), .A2(n1819), .B(n1216), .ZN(n1032) );
  INVD1BWP30P140LVT U1346 ( .I(pointer[4]), .ZN(n1335) );
  INVD1BWP30P140LVT U1347 ( .I(n1217), .ZN(n1340) );
  XOR2UD1BWP30P140LVT U1348 ( .A1(n1340), .A2(n1335), .Z(n1218) );
  MOAI22D1BWP30P140LVT U1349 ( .A1(n1335), .A2(n1748), .B1(n1218), .B2(n4), 
        .ZN(n1175) );
  INVD2BWP30P140LVT U1350 ( .I(n1219), .ZN(n1587) );
  INVD1BWP30P140LVT U1351 ( .I(delay_matrix_N_1[12]), .ZN(n1221) );
  OAI222D1BWP30P140LVT U1352 ( .A1(n1587), .A2(n2181), .B1(n1221), .B2(n1248), 
        .C1(n5), .C2(n1220), .ZN(n1007) );
  INVD1BWP30P140LVT U1353 ( .I(delay_matrix_N_1_next[26]), .ZN(n1226) );
  OAI222D1BWP30P140LVT U1354 ( .A1(n1587), .A2(n2185), .B1(n1222), .B2(n1933), 
        .C1(n5), .C2(n1226), .ZN(n993) );
  INVD1BWP30P140LVT U1355 ( .I(delay_matrix_N_1_next[41]), .ZN(n1753) );
  OAI22D1BWP30P140LVT U1356 ( .A1(n1225), .A2(n1224), .B1(n1223), .B2(n1753), 
        .ZN(n1056) );
  INVD1BWP30P140LVT U1357 ( .I(delay_matrix_N_1_next[40]), .ZN(n1586) );
  OAI22D1BWP30P140LVT U1358 ( .A1(n1229), .A2(n1224), .B1(n1223), .B2(n1586), 
        .ZN(n1057) );
  INVD1BWP30P140LVT U1359 ( .I(delay_matrix_N_1_next[27]), .ZN(n1242) );
  OAI22D1BWP30P140LVT U1360 ( .A1(n1225), .A2(n1228), .B1(n1227), .B2(n1242), 
        .ZN(n1020) );
  OAI22D1BWP30P140LVT U1361 ( .A1(n1229), .A2(n1228), .B1(n1227), .B2(n1226), 
        .ZN(n1021) );
  INVD1BWP30P140LVT U1362 ( .I(n1267), .ZN(n1233) );
  AOI21D1BWP30P140LVT U1363 ( .A1(n561), .A2(delay_matrix_N_1_next[24]), .B(
        n1807), .ZN(n1235) );
  OAI211D1BWP30P140LVT U1364 ( .A1(n1933), .A2(n1237), .B(n1236), .C(n1235), 
        .ZN(n995) );
  AOI21D1BWP30P140LVT U1365 ( .A1(n561), .A2(delay_matrix_N_1_next[38]), .B(
        n1807), .ZN(n1238) );
  OAI211D1BWP30P140LVT U1366 ( .A1(n1957), .A2(n1240), .B(n1239), .C(n1238), 
        .ZN(n981) );
  OAI222D1BWP30P140LVT U1367 ( .A1(n1751), .A2(n2185), .B1(n1243), .B2(n1933), 
        .C1(n5), .C2(n1242), .ZN(n992) );
  INVD1BWP30P140LVT U1368 ( .I(copy_pointer[1]), .ZN(n1244) );
  XNR2UD1BWP30P140LVT U1369 ( .A1(n1244), .A2(copy_pointer[0]), .ZN(n1246) );
  AO22D1BWP30P140LVT U1370 ( .A1(n4), .A2(n1246), .B1(n1245), .B2(
        copy_pointer[1]), .Z(n1146) );
  INVD1BWP30P140LVT U1371 ( .I(delay_matrix_N_1[13]), .ZN(n1249) );
  OAI222D1BWP30P140LVT U1372 ( .A1(n1751), .A2(n2181), .B1(n1249), .B2(n1248), 
        .C1(n5), .C2(n1247), .ZN(n1006) );
  AOI21D1BWP30P140LVT U1373 ( .A1(n561), .A2(delay_matrix_N_1_next[52]), .B(
        n1807), .ZN(n1250) );
  OAI211D1BWP30P140LVT U1374 ( .A1(n1988), .A2(n1252), .B(n1251), .C(n1250), 
        .ZN(n967) );
  AOI21D1BWP30P140LVT U1375 ( .A1(n1817), .A2(delay_matrix_N_1_next[32]), .B(
        n1807), .ZN(n1253) );
  OAI21D1BWP30P140LVT U1376 ( .A1(n1254), .A2(n1817), .B(n1253), .ZN(n1065) );
  INVD1BWP30P140LVT U1377 ( .I(n1255), .ZN(n1899) );
  NR2D1BWP30P140LVT U1378 ( .A1(n1899), .A2(n1256), .ZN(n1324) );
  INVD1BWP30P140LVT U1379 ( .I(copy_ptr_next[6]), .ZN(n1257) );
  XNR2UD1BWP30P140LVT U1380 ( .A1(n1324), .A2(n1257), .ZN(n1258) );
  MOAI22D1BWP30P140LVT U1381 ( .A1(n1835), .A2(n1257), .B1(n6), .B2(n1258), 
        .ZN(n949) );
  INVD1BWP30P140LVT U1382 ( .I(copy_ptr_next[8]), .ZN(n1259) );
  XNR2UD1BWP30P140LVT U1383 ( .A1(n1260), .A2(n1259), .ZN(n1261) );
  MOAI22D1BWP30P140LVT U1384 ( .A1(n1835), .A2(n1259), .B1(n6), .B2(n1261), 
        .ZN(n947) );
  ND2D1BWP30P140LVT U1385 ( .A1(n1262), .A2(copy_ptr_next[2]), .ZN(n1264) );
  INVD1BWP30P140LVT U1386 ( .I(copy_ptr_next[3]), .ZN(n1263) );
  XOR2UD1BWP30P140LVT U1387 ( .A1(n1264), .A2(n1263), .Z(n1265) );
  MOAI22D1BWP30P140LVT U1388 ( .A1(n1835), .A2(n1263), .B1(n6), .B2(n1265), 
        .ZN(n952) );
  INVD1BWP30P140LVT U1389 ( .I(n1269), .ZN(n1271) );
  ND2OPTIBD1BWP30P140LVT U1390 ( .A1(n1638), .A2(n1929), .ZN(n1275) );
  AOI21D1BWP30P140LVT U1391 ( .A1(n561), .A2(delay_matrix_N_1_next[25]), .B(
        n1807), .ZN(n1274) );
  OAI211D1BWP30P140LVT U1392 ( .A1(n1933), .A2(n1276), .B(n1275), .C(n1274), 
        .ZN(n994) );
  ND2OPTIBD1BWP30P140LVT U1393 ( .A1(n1638), .A2(n1953), .ZN(n1278) );
  AOI21D1BWP30P140LVT U1394 ( .A1(n561), .A2(delay_matrix_N_1_next[39]), .B(
        n1807), .ZN(n1277) );
  OAI211D1BWP30P140LVT U1395 ( .A1(n1957), .A2(n1279), .B(n1278), .C(n1277), 
        .ZN(n980) );
  AOI21D1BWP30P140LVT U1396 ( .A1(n1333), .A2(
        delay_matrix_N_1_next_original[51]), .B(n1280), .ZN(n1281) );
  OAI21D1BWP30P140LVT U1397 ( .A1(n1282), .A2(n1333), .B(n1281), .ZN(n914) );
  AOI21D1BWP30P140LVT U1398 ( .A1(n1815), .A2(delay_matrix_N_1_next[0]), .B(
        n1807), .ZN(n1283) );
  OAI21D1BWP30P140LVT U1399 ( .A1(n1646), .A2(n1815), .B(n1283), .ZN(n1047) );
  AOI21D1BWP30P140LVT U1400 ( .A1(n1392), .A2(
        delay_matrix_N_1_next_original[22]), .B(n1807), .ZN(n1284) );
  OAI21D1BWP30P140LVT U1401 ( .A1(n1776), .A2(n1392), .B(n1284), .ZN(n873) );
  INVD2BWP30P140LVT U1402 ( .I(delay_matrix_element[1]), .ZN(n1665) );
  AOI21D1BWP30P140LVT U1403 ( .A1(n1392), .A2(
        delay_matrix_N_1_next_original[15]), .B(n1807), .ZN(n1285) );
  OAI21D1BWP30P140LVT U1404 ( .A1(n1665), .A2(n1392), .B(n1285), .ZN(n880) );
  AOI21D1BWP30P140LVT U1405 ( .A1(n1392), .A2(
        delay_matrix_N_1_next_original[17]), .B(n1807), .ZN(n1286) );
  OAI21D1BWP30P140LVT U1406 ( .A1(n1678), .A2(n1392), .B(n1286), .ZN(n878) );
  INVD2BWP30P140LVT U1407 ( .I(delay_matrix_element[4]), .ZN(n1790) );
  AOI21D1BWP30P140LVT U1408 ( .A1(n1392), .A2(
        delay_matrix_N_1_next_original[18]), .B(n1807), .ZN(n1287) );
  OAI21D1BWP30P140LVT U1409 ( .A1(n1790), .A2(n1392), .B(n1287), .ZN(n877) );
  AOI21D1BWP30P140LVT U1410 ( .A1(n1398), .A2(
        delay_matrix_N_1_next_original[28]), .B(n1807), .ZN(n1288) );
  OAI21D1BWP30P140LVT U1411 ( .A1(n1793), .A2(n1398), .B(n1288), .ZN(n909) );
  AOI21D1BWP30P140LVT U1412 ( .A1(n1398), .A2(
        delay_matrix_N_1_next_original[31]), .B(n1807), .ZN(n1289) );
  OAI21D1BWP30P140LVT U1413 ( .A1(n1678), .A2(n1398), .B(n1289), .ZN(n906) );
  INVD2BWP30P140LVT U1414 ( .I(delay_matrix_element[7]), .ZN(n1779) );
  AOI21D1BWP30P140LVT U1415 ( .A1(n1398), .A2(
        delay_matrix_N_1_next_original[35]), .B(n1807), .ZN(n1290) );
  OAI21D1BWP30P140LVT U1416 ( .A1(n1779), .A2(n1398), .B(n1290), .ZN(n902) );
  AOI21D1BWP30P140LVT U1417 ( .A1(n1398), .A2(
        delay_matrix_N_1_next_original[29]), .B(n1807), .ZN(n1291) );
  OAI21D1BWP30P140LVT U1418 ( .A1(n1665), .A2(n1398), .B(n1291), .ZN(n908) );
  AOI21D1BWP30P140LVT U1419 ( .A1(n1404), .A2(
        delay_matrix_N_1_next_original[1]), .B(n1807), .ZN(n1292) );
  OAI21D1BWP30P140LVT U1420 ( .A1(n1665), .A2(n1404), .B(n1292), .ZN(n894) );
  AOI21D1BWP30P140LVT U1421 ( .A1(n1404), .A2(
        delay_matrix_N_1_next_original[4]), .B(n1807), .ZN(n1293) );
  OAI21D1BWP30P140LVT U1422 ( .A1(n1790), .A2(n1404), .B(n1293), .ZN(n891) );
  AOI21D1BWP30P140LVT U1423 ( .A1(n1404), .A2(
        delay_matrix_N_1_next_original[3]), .B(n1807), .ZN(n1294) );
  OAI21D1BWP30P140LVT U1424 ( .A1(n1678), .A2(n1404), .B(n1294), .ZN(n892) );
  ND2OPTIBD1BWP30P140LVT U1425 ( .A1(n1638), .A2(n1982), .ZN(n1296) );
  AOI21D1BWP30P140LVT U1426 ( .A1(n561), .A2(delay_matrix_N_1_next[53]), .B(
        n1807), .ZN(n1295) );
  OAI211D1BWP30P140LVT U1427 ( .A1(n1988), .A2(n1297), .B(n1296), .C(n1295), 
        .ZN(n966) );
  AOI21D1BWP30P140LVT U1428 ( .A1(n1333), .A2(
        delay_matrix_N_1_next_original[45]), .B(n1807), .ZN(n1298) );
  OAI21D1BWP30P140LVT U1429 ( .A1(n1678), .A2(n1333), .B(n1298), .ZN(n920) );
  AOI21D1BWP30P140LVT U1430 ( .A1(n1333), .A2(
        delay_matrix_N_1_next_original[49]), .B(n1807), .ZN(n1299) );
  OAI21D1BWP30P140LVT U1431 ( .A1(n1779), .A2(n1333), .B(n1299), .ZN(n916) );
  AOI21D1BWP30P140LVT U1432 ( .A1(n1333), .A2(
        delay_matrix_N_1_next_original[43]), .B(n1807), .ZN(n1300) );
  OAI21D1BWP30P140LVT U1433 ( .A1(n1665), .A2(n1333), .B(n1300), .ZN(n922) );
  AOI21D1BWP30P140LVT U1434 ( .A1(n1819), .A2(delay_matrix_N_1_next[22]), .B(
        n1807), .ZN(n1301) );
  OAI21D1BWP30P140LVT U1435 ( .A1(n1565), .A2(n1819), .B(n1301), .ZN(n1025) );
  AOI21D1BWP30P140LVT U1436 ( .A1(n1813), .A2(delay_matrix_N_1_next[50]), .B(
        n1807), .ZN(n1302) );
  OAI21D1BWP30P140LVT U1437 ( .A1(n1565), .A2(n1813), .B(n1302), .ZN(n1075) );
  OAI222D1BWP30P140LVT U1438 ( .A1(n1304), .A2(n5), .B1(n1303), .B2(n1988), 
        .C1(n1461), .C2(n1587), .ZN(n965) );
  MUX2NUD1BWP30P140LVT U1439 ( .I0(n1631), .I1(delay_matrix_N_1_next[10]), .S(
        n1815), .ZN(n1305) );
  MUX2NUD1BWP30P140LVT U1440 ( .I0(n1631), .I1(delay_matrix_N_1_next[52]), .S(
        n1813), .ZN(n1306) );
  AOI21D1BWP30P140LVT U1441 ( .A1(n1815), .A2(delay_matrix_N_1_next[8]), .B(
        n1807), .ZN(n1307) );
  OAI21D1BWP30P140LVT U1442 ( .A1(n1565), .A2(n1815), .B(n1307), .ZN(n1039) );
  OAI21D1BWP30P140LVT U1443 ( .A1(n1310), .A2(n1309), .B(n1308), .ZN(n1315) );
  INVD1BWP30P140LVT U1444 ( .I(n1311), .ZN(n1313) );
  AOI21D1BWP30P140LVT U1445 ( .A1(n561), .A2(delay_matrix_N_1_next[21]), .B(
        n1807), .ZN(n1316) );
  OAI211D1BWP30P140LVT U1446 ( .A1(n1933), .A2(n1318), .B(n1317), .C(n1316), 
        .ZN(n998) );
  INVD1BWP30P140LVT U1447 ( .I(delay_matrix_N_1[35]), .ZN(n1321) );
  AOI21D1BWP30P140LVT U1448 ( .A1(n561), .A2(delay_matrix_N_1_next[35]), .B(
        n1807), .ZN(n1319) );
  OAI211D1BWP30P140LVT U1449 ( .A1(n1957), .A2(n1321), .B(n1320), .C(n1319), 
        .ZN(n984) );
  MUX2NUD1BWP30P140LVT U1450 ( .I0(n1631), .I1(delay_matrix_N_1_next[24]), .S(
        n1819), .ZN(n1322) );
  MUX2NUD1BWP30P140LVT U1451 ( .I0(n1631), .I1(delay_matrix_N_1_next[38]), .S(
        n1817), .ZN(n1323) );
  ND2D1BWP30P140LVT U1452 ( .A1(n1324), .A2(copy_ptr_next[6]), .ZN(n1326) );
  INVD1BWP30P140LVT U1453 ( .I(copy_ptr_next[7]), .ZN(n1325) );
  XOR2UD1BWP30P140LVT U1454 ( .A1(n1326), .A2(n1325), .Z(n1327) );
  MOAI22D1BWP30P140LVT U1455 ( .A1(n1835), .A2(n1325), .B1(n6), .B2(n1327), 
        .ZN(n948) );
  INVD1BWP30P140LVT U1456 ( .I(copy_ptr_next[4]), .ZN(n1898) );
  NR2D1BWP30P140LVT U1457 ( .A1(n1899), .A2(n1898), .ZN(n1329) );
  INVD1BWP30P140LVT U1458 ( .I(copy_ptr_next[5]), .ZN(n1328) );
  XNR2UD1BWP30P140LVT U1459 ( .A1(n1329), .A2(n1328), .ZN(n1330) );
  MOAI22D1BWP30P140LVT U1460 ( .A1(n1835), .A2(n1328), .B1(n6), .B2(n1330), 
        .ZN(n950) );
  AOI21D1BWP30P140LVT U1461 ( .A1(n1817), .A2(delay_matrix_N_1_next[36]), .B(
        n1807), .ZN(n1331) );
  OAI21D1BWP30P140LVT U1462 ( .A1(n1565), .A2(n1817), .B(n1331), .ZN(n1061) );
  OAI211D1BWP30P140LVT U1463 ( .A1(n2203), .A2(n1333), .B(n1332), .C(n1821), 
        .ZN(n910) );
  OAI211D1BWP30P140LVT U1464 ( .A1(n2199), .A2(n1333), .B(n1334), .C(n1821), 
        .ZN(n911) );
  INVD1BWP30P140LVT U1465 ( .I(pointer[5]), .ZN(n1338) );
  NR2D1BWP30P140LVT U1466 ( .A1(n1340), .A2(n1335), .ZN(n1336) );
  XNR2UD1BWP30P140LVT U1467 ( .A1(n1336), .A2(n1338), .ZN(n1337) );
  MOAI22D1BWP30P140LVT U1468 ( .A1(n1338), .A2(n1616), .B1(n4), .B2(n1337), 
        .ZN(n1174) );
  INVD1BWP30P140LVT U1469 ( .I(pointer[6]), .ZN(n1342) );
  NR2D1BWP30P140LVT U1470 ( .A1(n1340), .A2(n1339), .ZN(n1373) );
  XNR2UD1BWP30P140LVT U1471 ( .A1(n1373), .A2(n1342), .ZN(n1341) );
  MOAI22D1BWP30P140LVT U1472 ( .A1(n1342), .A2(n1616), .B1(n4), .B2(n1341), 
        .ZN(n1173) );
  INVD1BWP30P140LVT U1473 ( .I(pointer[17]), .ZN(n1346) );
  INVD1BWP30P140LVT U1474 ( .I(pointer[16]), .ZN(n1367) );
  NR2D1BWP30P140LVT U1475 ( .A1(n1445), .A2(n1367), .ZN(n1344) );
  XNR2UD1BWP30P140LVT U1476 ( .A1(n1344), .A2(n1346), .ZN(n1345) );
  MOAI22D1BWP30P140LVT U1477 ( .A1(n1346), .A2(n1616), .B1(n4), .B2(n1345), 
        .ZN(n1162) );
  INVD1BWP30P140LVT U1478 ( .I(pointer[15]), .ZN(n1353) );
  INVD1BWP30P140LVT U1479 ( .I(n1377), .ZN(n1381) );
  INVD1BWP30P140LVT U1480 ( .I(n1349), .ZN(n1350) );
  INVD1BWP30P140LVT U1481 ( .I(pointer[14]), .ZN(n1356) );
  NR2D1BWP30P140LVT U1482 ( .A1(n1354), .A2(n1356), .ZN(n1351) );
  XNR2UD1BWP30P140LVT U1483 ( .A1(n1351), .A2(n1353), .ZN(n1352) );
  MOAI22D1BWP30P140LVT U1484 ( .A1(n1353), .A2(n1616), .B1(n4), .B2(n1352), 
        .ZN(n1164) );
  XOR2UD1BWP30P140LVT U1485 ( .A1(n1354), .A2(n1356), .Z(n1355) );
  MOAI22D1BWP30P140LVT U1486 ( .A1(n1356), .A2(n1616), .B1(n4), .B2(n1355), 
        .ZN(n1165) );
  INVD1BWP30P140LVT U1487 ( .I(pointer[9]), .ZN(n1359) );
  ND2D1BWP30P140LVT U1488 ( .A1(n1364), .A2(pointer[8]), .ZN(n1357) );
  XOR2UD1BWP30P140LVT U1489 ( .A1(n1357), .A2(n1359), .Z(n1358) );
  MOAI22D1BWP30P140LVT U1490 ( .A1(n1359), .A2(n1616), .B1(n4), .B2(n1358), 
        .ZN(n1170) );
  INVD1BWP30P140LVT U1491 ( .I(pointer[8]), .ZN(n1361) );
  XNR2UD1BWP30P140LVT U1492 ( .A1(n1364), .A2(n1361), .ZN(n1360) );
  MOAI22D1BWP30P140LVT U1493 ( .A1(n1361), .A2(n1616), .B1(n4), .B2(n1360), 
        .ZN(n1171) );
  INVD1BWP30P140LVT U1494 ( .I(pointer[10]), .ZN(n1368) );
  INVD1BWP30P140LVT U1495 ( .I(n1362), .ZN(n1363) );
  ND2D1BWP30P140LVT U1496 ( .A1(n1364), .A2(n1363), .ZN(n1369) );
  XOR2UD1BWP30P140LVT U1497 ( .A1(n1369), .A2(n1368), .Z(n1365) );
  MOAI22D1BWP30P140LVT U1498 ( .A1(n1368), .A2(n1616), .B1(n4), .B2(n1365), 
        .ZN(n1169) );
  XOR2UD1BWP30P140LVT U1499 ( .A1(n1445), .A2(n1367), .Z(n1366) );
  MOAI22D1BWP30P140LVT U1500 ( .A1(n1367), .A2(n1616), .B1(n4), .B2(n1366), 
        .ZN(n1163) );
  INVD1BWP30P140LVT U1501 ( .I(pointer[11]), .ZN(n1372) );
  NR2D1BWP30P140LVT U1502 ( .A1(n1369), .A2(n1368), .ZN(n1370) );
  XNR2UD1BWP30P140LVT U1503 ( .A1(n1370), .A2(n1372), .ZN(n1371) );
  MOAI22D1BWP30P140LVT U1504 ( .A1(n1372), .A2(n1616), .B1(n4), .B2(n1371), 
        .ZN(n1168) );
  INVD1BWP30P140LVT U1505 ( .I(pointer[7]), .ZN(n1376) );
  ND2D1BWP30P140LVT U1506 ( .A1(n1373), .A2(pointer[6]), .ZN(n1374) );
  XOR2UD1BWP30P140LVT U1507 ( .A1(n1374), .A2(n1376), .Z(n1375) );
  MOAI22D1BWP30P140LVT U1508 ( .A1(n1376), .A2(n1616), .B1(n4), .B2(n1375), 
        .ZN(n1172) );
  INVD1BWP30P140LVT U1509 ( .I(pointer[13]), .ZN(n1380) );
  INVD1BWP30P140LVT U1510 ( .I(pointer[12]), .ZN(n1383) );
  NR2D1BWP30P140LVT U1511 ( .A1(n1377), .A2(n1383), .ZN(n1378) );
  XNR2UD1BWP30P140LVT U1512 ( .A1(n1378), .A2(n1380), .ZN(n1379) );
  MOAI22D1BWP30P140LVT U1513 ( .A1(n1380), .A2(n1616), .B1(n4), .B2(n1379), 
        .ZN(n1166) );
  XNR2UD1BWP30P140LVT U1514 ( .A1(n1381), .A2(n1383), .ZN(n1382) );
  MOAI22D1BWP30P140LVT U1515 ( .A1(n1383), .A2(n1616), .B1(n4), .B2(n1382), 
        .ZN(n1167) );
  INVD1BWP30P140LVT U1516 ( .I(pointer[30]), .ZN(n1386) );
  HA1D1BWP30P140LVT U1517 ( .A(pointer[30]), .B(n1384), .CO(n219), .S(n1385)
         );
  MOAI22D1BWP30P140LVT U1518 ( .A1(n1386), .A2(n1616), .B1(n4), .B2(n1385), 
        .ZN(n1149) );
  AOI21D1BWP30P140LVT U1519 ( .A1(n1392), .A2(
        delay_matrix_N_1_next_original[19]), .B(n1807), .ZN(n1387) );
  OAI21D1BWP30P140LVT U1520 ( .A1(n1798), .A2(n1392), .B(n1387), .ZN(n876) );
  AOI21D1BWP30P140LVT U1521 ( .A1(n1392), .A2(
        delay_matrix_N_1_next_original[21]), .B(n1807), .ZN(n1388) );
  OAI21D1BWP30P140LVT U1522 ( .A1(n1779), .A2(n1392), .B(n1388), .ZN(n874) );
  AOI21D1BWP30P140LVT U1523 ( .A1(n1392), .A2(
        delay_matrix_N_1_next_original[14]), .B(n1807), .ZN(n1389) );
  OAI21D1BWP30P140LVT U1524 ( .A1(n1793), .A2(n1392), .B(n1389), .ZN(n881) );
  INVD2BWP30P140LVT U1525 ( .I(delay_matrix_element[6]), .ZN(n1805) );
  AOI21D1BWP30P140LVT U1526 ( .A1(n1392), .A2(
        delay_matrix_N_1_next_original[20]), .B(n1807), .ZN(n1390) );
  OAI21D1BWP30P140LVT U1527 ( .A1(n1805), .A2(n1392), .B(n1390), .ZN(n875) );
  AOI21D1BWP30P140LVT U1528 ( .A1(n1392), .A2(
        delay_matrix_N_1_next_original[16]), .B(n1807), .ZN(n1391) );
  OAI21D1BWP30P140LVT U1529 ( .A1(n1810), .A2(n1392), .B(n1391), .ZN(n879) );
  AOI21D1BWP30P140LVT U1530 ( .A1(n1398), .A2(
        delay_matrix_N_1_next_original[33]), .B(n1807), .ZN(n1393) );
  OAI21D1BWP30P140LVT U1531 ( .A1(n1798), .A2(n1398), .B(n1393), .ZN(n904) );
  AOI21D1BWP30P140LVT U1532 ( .A1(n1398), .A2(
        delay_matrix_N_1_next_original[36]), .B(n1807), .ZN(n1394) );
  OAI21D1BWP30P140LVT U1533 ( .A1(n1776), .A2(n1398), .B(n1394), .ZN(n901) );
  AOI21D1BWP30P140LVT U1534 ( .A1(n1398), .A2(
        delay_matrix_N_1_next_original[30]), .B(n1807), .ZN(n1395) );
  OAI21D1BWP30P140LVT U1535 ( .A1(n1810), .A2(n1398), .B(n1395), .ZN(n907) );
  AOI21D1BWP30P140LVT U1536 ( .A1(n1398), .A2(
        delay_matrix_N_1_next_original[34]), .B(n1807), .ZN(n1396) );
  OAI21D1BWP30P140LVT U1537 ( .A1(n1805), .A2(n1398), .B(n1396), .ZN(n903) );
  AOI21D1BWP30P140LVT U1538 ( .A1(n1398), .A2(
        delay_matrix_N_1_next_original[32]), .B(n1807), .ZN(n1397) );
  OAI21D1BWP30P140LVT U1539 ( .A1(n1790), .A2(n1398), .B(n1397), .ZN(n905) );
  AOI21D1BWP30P140LVT U1540 ( .A1(n1404), .A2(
        delay_matrix_N_1_next_original[2]), .B(n1807), .ZN(n1399) );
  OAI21D1BWP30P140LVT U1541 ( .A1(n1810), .A2(n1404), .B(n1399), .ZN(n893) );
  AOI21D1BWP30P140LVT U1542 ( .A1(n1404), .A2(
        delay_matrix_N_1_next_original[6]), .B(n1807), .ZN(n1400) );
  OAI21D1BWP30P140LVT U1543 ( .A1(n1805), .A2(n1404), .B(n1400), .ZN(n889) );
  AOI21D1BWP30P140LVT U1544 ( .A1(n1404), .A2(
        delay_matrix_N_1_next_original[0]), .B(n1807), .ZN(n1401) );
  OAI21D1BWP30P140LVT U1545 ( .A1(n1793), .A2(n1404), .B(n1401), .ZN(n895) );
  AOI21D1BWP30P140LVT U1546 ( .A1(n1404), .A2(
        delay_matrix_N_1_next_original[5]), .B(n1807), .ZN(n1402) );
  OAI21D1BWP30P140LVT U1547 ( .A1(n1798), .A2(n1404), .B(n1402), .ZN(n890) );
  AOI21D1BWP30P140LVT U1548 ( .A1(n1404), .A2(
        delay_matrix_N_1_next_original[7]), .B(n1807), .ZN(n1403) );
  OAI21D1BWP30P140LVT U1549 ( .A1(n1779), .A2(n1404), .B(n1403), .ZN(n888) );
  OAI21D1BWP30P140LVT U1550 ( .A1(n1407), .A2(n1406), .B(n1405), .ZN(n1412) );
  INVD1BWP30P140LVT U1551 ( .I(n1408), .ZN(n1410) );
  ND2OPTIBD1BWP30P140LVT U1552 ( .A1(n1820), .A2(n1929), .ZN(n1414) );
  AOI21D1BWP30P140LVT U1553 ( .A1(n561), .A2(delay_matrix_N_1_next[23]), .B(
        n1807), .ZN(n1413) );
  OAI211D1BWP30P140LVT U1554 ( .A1(n1933), .A2(n1415), .B(n1414), .C(n1413), 
        .ZN(n996) );
  ND2OPTIBD1BWP30P140LVT U1555 ( .A1(n1820), .A2(n1953), .ZN(n1417) );
  AOI21D1BWP30P140LVT U1556 ( .A1(n561), .A2(delay_matrix_N_1_next[37]), .B(
        n1807), .ZN(n1416) );
  OAI211D1BWP30P140LVT U1557 ( .A1(n1957), .A2(n1418), .B(n1417), .C(n1416), 
        .ZN(n982) );
  INVD1BWP30P140LVT U1558 ( .I(pointer[29]), .ZN(n1421) );
  HA1D1BWP30P140LVT U1559 ( .A(pointer[29]), .B(n1419), .CO(n1384), .S(n1420)
         );
  MOAI22D1BWP30P140LVT U1560 ( .A1(n1421), .A2(n1616), .B1(n4), .B2(n1420), 
        .ZN(n1150) );
  INVD1BWP30P140LVT U1561 ( .I(pointer[20]), .ZN(n1425) );
  INVD1BWP30P140LVT U1562 ( .I(n1422), .ZN(n1423) );
  NR2D1BWP30P140LVT U1563 ( .A1(n1445), .A2(n1423), .ZN(n1440) );
  INVD1BWP30P140LVT U1564 ( .I(n1440), .ZN(n1427) );
  XOR2UD1BWP30P140LVT U1565 ( .A1(n1427), .A2(n1425), .Z(n1424) );
  MOAI22D1BWP30P140LVT U1566 ( .A1(n1425), .A2(n1616), .B1(n4), .B2(n1424), 
        .ZN(n1159) );
  INVD1BWP30P140LVT U1567 ( .I(pointer[22]), .ZN(n1429) );
  NR2D1BWP30P140LVT U1568 ( .A1(n1427), .A2(n1426), .ZN(n1436) );
  XNR2UD1BWP30P140LVT U1569 ( .A1(n1436), .A2(n1429), .ZN(n1428) );
  MOAI22D1BWP30P140LVT U1570 ( .A1(n1429), .A2(n1616), .B1(n4), .B2(n1428), 
        .ZN(n1157) );
  INVD1BWP30P140LVT U1571 ( .I(pointer[18]), .ZN(n1432) );
  NR2D1BWP30P140LVT U1572 ( .A1(n1445), .A2(n1430), .ZN(n1454) );
  XNR2UD1BWP30P140LVT U1573 ( .A1(n1454), .A2(n1432), .ZN(n1431) );
  MOAI22D1BWP30P140LVT U1574 ( .A1(n1432), .A2(n1616), .B1(n4), .B2(n1431), 
        .ZN(n1161) );
  INVD1BWP30P140LVT U1575 ( .I(pointer[27]), .ZN(n1435) );
  HA1D1BWP30P140LVT U1576 ( .A(pointer[27]), .B(n1433), .CO(n1458), .S(n1434)
         );
  MOAI22D1BWP30P140LVT U1577 ( .A1(n1435), .A2(n1616), .B1(n4), .B2(n1434), 
        .ZN(n1152) );
  INVD1BWP30P140LVT U1578 ( .I(pointer[23]), .ZN(n1439) );
  XOR2UD1BWP30P140LVT U1579 ( .A1(n1437), .A2(n1439), .Z(n1438) );
  MOAI22D1BWP30P140LVT U1580 ( .A1(n1439), .A2(n1616), .B1(n4), .B2(n1438), 
        .ZN(n1156) );
  INVD1BWP30P140LVT U1581 ( .I(pointer[21]), .ZN(n1443) );
  XOR2UD1BWP30P140LVT U1582 ( .A1(n1441), .A2(n1443), .Z(n1442) );
  MOAI22D1BWP30P140LVT U1583 ( .A1(n1443), .A2(n1616), .B1(n4), .B2(n1442), 
        .ZN(n1158) );
  INVD1BWP30P140LVT U1584 ( .I(pointer[25]), .ZN(n1448) );
  NR2D1BWP30P140LVT U1585 ( .A1(n1445), .A2(n1444), .ZN(n1449) );
  XOR2UD1BWP30P140LVT U1586 ( .A1(n1446), .A2(n1448), .Z(n1447) );
  MOAI22D1BWP30P140LVT U1587 ( .A1(n1448), .A2(n1616), .B1(n4), .B2(n1447), 
        .ZN(n1154) );
  INVD1BWP30P140LVT U1588 ( .I(pointer[24]), .ZN(n1451) );
  XNR2UD1BWP30P140LVT U1589 ( .A1(n1449), .A2(n1451), .ZN(n1450) );
  MOAI22D1BWP30P140LVT U1590 ( .A1(n1451), .A2(n1616), .B1(n4), .B2(n1450), 
        .ZN(n1155) );
  INVD1BWP30P140LVT U1591 ( .I(pointer[26]), .ZN(n1453) );
  HA1D1BWP30P140LVT U1592 ( .A(pointer[26]), .B(n14), .CO(n1433), .S(n1452) );
  MOAI22D1BWP30P140LVT U1593 ( .A1(n1453), .A2(n1616), .B1(n4), .B2(n1452), 
        .ZN(n1153) );
  INVD1BWP30P140LVT U1594 ( .I(pointer[19]), .ZN(n1457) );
  XOR2UD1BWP30P140LVT U1595 ( .A1(n1455), .A2(n1457), .Z(n1456) );
  MOAI22D1BWP30P140LVT U1596 ( .A1(n1457), .A2(n1616), .B1(n4), .B2(n1456), 
        .ZN(n1160) );
  INVD1BWP30P140LVT U1597 ( .I(pointer[28]), .ZN(n1460) );
  HA1D1BWP30P140LVT U1598 ( .A(pointer[28]), .B(n1458), .CO(n1419), .S(n1459)
         );
  MOAI22D1BWP30P140LVT U1599 ( .A1(n1460), .A2(n1616), .B1(n4), .B2(n1459), 
        .ZN(n1151) );
  OAI222D1BWP30P140LVT U1600 ( .A1(n1463), .A2(n5), .B1(n1462), .B2(n1988), 
        .C1(n1461), .C2(n1751), .ZN(n964) );
  OAI211D1BWP30P140LVT U1601 ( .A1(n1465), .A2(n1333), .B(n1464), .C(n1821), 
        .ZN(n912) );
  AOI21D1BWP30P140LVT U1602 ( .A1(n1819), .A2(delay_matrix_N_1_next[20]), .B(
        n1807), .ZN(n1466) );
  OAI21D1BWP30P140LVT U1603 ( .A1(n1637), .A2(n1819), .B(n1466), .ZN(n1027) );
  AOI21D1BWP30P140LVT U1604 ( .A1(n1815), .A2(delay_matrix_N_1_next[6]), .B(
        n1807), .ZN(n1467) );
  OAI21D1BWP30P140LVT U1605 ( .A1(n1637), .A2(n1815), .B(n1467), .ZN(n1041) );
  AOI21D1BWP30P140LVT U1606 ( .A1(n1817), .A2(delay_matrix_N_1_next[34]), .B(
        n1807), .ZN(n1468) );
  OAI21D1BWP30P140LVT U1607 ( .A1(n1637), .A2(n1817), .B(n1468), .ZN(n1063) );
  AOI21D1BWP30P140LVT U1608 ( .A1(n1813), .A2(delay_matrix_N_1_next[48]), .B(
        n1807), .ZN(n1469) );
  OAI21D1BWP30P140LVT U1609 ( .A1(n1637), .A2(n1813), .B(n1469), .ZN(n1077) );
  INVD1BWP30P140LVT U1610 ( .I(n1470), .ZN(n1833) );
  INVD1BWP30P140LVT U1611 ( .I(ptr_next[4]), .ZN(n1832) );
  NR2D1BWP30P140LVT U1612 ( .A1(n1833), .A2(n1832), .ZN(n1472) );
  INVD1BWP30P140LVT U1613 ( .I(ptr_next[5]), .ZN(n1471) );
  XNR2UD1BWP30P140LVT U1614 ( .A1(n1472), .A2(n1471), .ZN(n1473) );
  MOAI22D1BWP30P140LVT U1615 ( .A1(n1471), .A2(n1835), .B1(n6), .B2(n1473), 
        .ZN(n1110) );
  NR2D1BWP30P140LVT U1616 ( .A1(n1833), .A2(n1474), .ZN(n1477) );
  INVD1BWP30P140LVT U1617 ( .I(ptr_next[6]), .ZN(n1475) );
  XNR2UD1BWP30P140LVT U1618 ( .A1(n1477), .A2(n1475), .ZN(n1476) );
  MOAI22D1BWP30P140LVT U1619 ( .A1(n1475), .A2(n1835), .B1(n6), .B2(n1476), 
        .ZN(n1109) );
  ND2D1BWP30P140LVT U1620 ( .A1(n1477), .A2(ptr_next[6]), .ZN(n1479) );
  INVD1BWP30P140LVT U1621 ( .I(ptr_next[7]), .ZN(n1478) );
  XOR2UD1BWP30P140LVT U1622 ( .A1(n1479), .A2(n1478), .Z(n1480) );
  MOAI22D1BWP30P140LVT U1623 ( .A1(n1478), .A2(n1835), .B1(n6), .B2(n1480), 
        .ZN(n1108) );
  INVD1BWP30P140LVT U1624 ( .I(copy_pointer[26]), .ZN(n1494) );
  ND2D1BWP30P140LVT U1625 ( .A1(copy_pointer[18]), .A2(copy_pointer[19]), .ZN(
        n1481) );
  NR2D1BWP30P140LVT U1626 ( .A1(n1501), .A2(n1481), .ZN(n1496) );
  ND2D1BWP30P140LVT U1627 ( .A1(copy_pointer[22]), .A2(copy_pointer[23]), .ZN(
        n1482) );
  NR2D1BWP30P140LVT U1628 ( .A1(n1530), .A2(n1482), .ZN(n1483) );
  NR2D1BWP30P140LVT U1629 ( .A1(n1520), .A2(n1484), .ZN(n1492) );
  NR2D1BWP30P140LVT U1630 ( .A1(n1524), .A2(n1485), .ZN(n1509) );
  ND2D1BWP30P140LVT U1631 ( .A1(copy_pointer[14]), .A2(copy_pointer[15]), .ZN(
        n1486) );
  NR2D1BWP30P140LVT U1632 ( .A1(n1510), .A2(n1486), .ZN(n1487) );
  NR2D1BWP30P140LVT U1633 ( .A1(n1535), .A2(n1488), .ZN(n1490) );
  MOAI22D1BWP30P140LVT U1634 ( .A1(n1616), .A2(n1494), .B1(n4), .B2(n1493), 
        .ZN(n1121) );
  INVD1BWP30P140LVT U1635 ( .I(n1496), .ZN(n1497) );
  NR2D1BWP30P140LVT U1636 ( .A1(n1540), .A2(n1497), .ZN(n1527) );
  INVD1BWP30P140LVT U1637 ( .I(copy_pointer[21]), .ZN(n1498) );
  XOR2UD1BWP30P140LVT U1638 ( .A1(n1499), .A2(n1498), .Z(n1500) );
  MOAI22D1BWP30P140LVT U1639 ( .A1(n1616), .A2(n1498), .B1(n4), .B2(n1500), 
        .ZN(n1126) );
  NR2D1BWP30P140LVT U1640 ( .A1(n1540), .A2(n1501), .ZN(n1548) );
  ND2D1BWP30P140LVT U1641 ( .A1(n1548), .A2(copy_pointer[18]), .ZN(n1503) );
  INVD1BWP30P140LVT U1642 ( .I(copy_pointer[19]), .ZN(n1502) );
  XOR2UD1BWP30P140LVT U1643 ( .A1(n1503), .A2(n1502), .Z(n1504) );
  MOAI22D1BWP30P140LVT U1644 ( .A1(n1616), .A2(n1502), .B1(n4), .B2(n1504), 
        .ZN(n1128) );
  INVD1BWP30P140LVT U1645 ( .I(copy_pointer[16]), .ZN(n1539) );
  XOR2UD1BWP30P140LVT U1646 ( .A1(n1540), .A2(n1539), .Z(n1505) );
  MOAI22D1BWP30P140LVT U1647 ( .A1(n1616), .A2(n1539), .B1(n4), .B2(n1505), 
        .ZN(n1131) );
  HA1D1BWP30P140LVT U1648 ( .A(copy_pointer[26]), .B(n15), .CO(n1517), .S(
        n1493) );
  MOAI22D1BWP30P140LVT U1649 ( .A1(n1616), .A2(n1507), .B1(n4), .B2(n1506), 
        .ZN(n1117) );
  INVD1BWP30P140LVT U1650 ( .I(n1513), .ZN(n1573) );
  INVD1BWP30P140LVT U1651 ( .I(n1510), .ZN(n1511) );
  ND2D1BWP30P140LVT U1652 ( .A1(n1573), .A2(n1511), .ZN(n1604) );
  INVD1BWP30P140LVT U1653 ( .I(copy_pointer[14]), .ZN(n1603) );
  XOR2UD1BWP30P140LVT U1654 ( .A1(n1604), .A2(n1603), .Z(n1512) );
  MOAI22D1BWP30P140LVT U1655 ( .A1(n1616), .A2(n1603), .B1(n4), .B2(n1512), 
        .ZN(n1133) );
  INVD1BWP30P140LVT U1656 ( .I(copy_pointer[12]), .ZN(n1572) );
  NR2D1BWP30P140LVT U1657 ( .A1(n1513), .A2(n1572), .ZN(n1515) );
  INVD1BWP30P140LVT U1658 ( .I(copy_pointer[13]), .ZN(n1514) );
  XNR2UD1BWP30P140LVT U1659 ( .A1(n1515), .A2(n1514), .ZN(n1516) );
  MOAI22D1BWP30P140LVT U1660 ( .A1(n1616), .A2(n1514), .B1(n4), .B2(n1516), 
        .ZN(n1134) );
  INVD1BWP30P140LVT U1661 ( .I(copy_pointer[27]), .ZN(n1519) );
  HA1D1BWP30P140LVT U1662 ( .A(copy_pointer[27]), .B(n1517), .CO(n1600), .S(
        n1518) );
  MOAI22D1BWP30P140LVT U1663 ( .A1(n1616), .A2(n1519), .B1(n4), .B2(n1518), 
        .ZN(n1120) );
  NR2D1BWP30P140LVT U1664 ( .A1(n1540), .A2(n1520), .ZN(n1545) );
  INVD1BWP30P140LVT U1665 ( .I(copy_pointer[25]), .ZN(n1521) );
  XOR2UD1BWP30P140LVT U1666 ( .A1(n1522), .A2(n1521), .Z(n1523) );
  MOAI22D1BWP30P140LVT U1667 ( .A1(n1616), .A2(n1521), .B1(n4), .B2(n1523), 
        .ZN(n1122) );
  INVD1BWP30P140LVT U1668 ( .I(n1524), .ZN(n1525) );
  ND2D1BWP30P140LVT U1669 ( .A1(n1614), .A2(n1525), .ZN(n1609) );
  INVD1BWP30P140LVT U1670 ( .I(copy_pointer[10]), .ZN(n1608) );
  XOR2UD1BWP30P140LVT U1671 ( .A1(n1609), .A2(n1608), .Z(n1526) );
  MOAI22D1BWP30P140LVT U1672 ( .A1(n1616), .A2(n1608), .B1(n4), .B2(n1526), 
        .ZN(n1137) );
  INVD1BWP30P140LVT U1673 ( .I(n1527), .ZN(n1531) );
  INVD1BWP30P140LVT U1674 ( .I(copy_pointer[20]), .ZN(n1528) );
  XOR2UD1BWP30P140LVT U1675 ( .A1(n1531), .A2(n1528), .Z(n1529) );
  MOAI22D1BWP30P140LVT U1676 ( .A1(n1616), .A2(n1528), .B1(n4), .B2(n1529), 
        .ZN(n1127) );
  NR2D1BWP30P140LVT U1677 ( .A1(n1531), .A2(n1530), .ZN(n1582) );
  INVD1BWP30P140LVT U1678 ( .I(copy_pointer[23]), .ZN(n1532) );
  XOR2UD1BWP30P140LVT U1679 ( .A1(n1533), .A2(n1532), .Z(n1534) );
  MOAI22D1BWP30P140LVT U1680 ( .A1(n1616), .A2(n1532), .B1(n4), .B2(n1534), 
        .ZN(n1124) );
  NR2D1BWP30P140LVT U1681 ( .A1(n1593), .A2(n1535), .ZN(n1579) );
  ND2D1BWP30P140LVT U1682 ( .A1(n1579), .A2(copy_pointer[6]), .ZN(n1537) );
  INVD1BWP30P140LVT U1683 ( .I(copy_pointer[7]), .ZN(n1536) );
  XOR2UD1BWP30P140LVT U1684 ( .A1(n1537), .A2(n1536), .Z(n1538) );
  MOAI22D1BWP30P140LVT U1685 ( .A1(n1616), .A2(n1536), .B1(n4), .B2(n1538), 
        .ZN(n1140) );
  NR2D1BWP30P140LVT U1686 ( .A1(n1540), .A2(n1539), .ZN(n1542) );
  INVD1BWP30P140LVT U1687 ( .I(copy_pointer[17]), .ZN(n1541) );
  XNR2UD1BWP30P140LVT U1688 ( .A1(n1542), .A2(n1541), .ZN(n1543) );
  MOAI22D1BWP30P140LVT U1689 ( .A1(n1616), .A2(n1541), .B1(n4), .B2(n1543), 
        .ZN(n1130) );
  INVD1BWP30P140LVT U1690 ( .I(copy_pointer[24]), .ZN(n1544) );
  XNR2UD1BWP30P140LVT U1691 ( .A1(n1545), .A2(n1544), .ZN(n1546) );
  MOAI22D1BWP30P140LVT U1692 ( .A1(n1616), .A2(n1544), .B1(n4), .B2(n1546), 
        .ZN(n1123) );
  INVD1BWP30P140LVT U1693 ( .I(copy_pointer[18]), .ZN(n1547) );
  XNR2UD1BWP30P140LVT U1694 ( .A1(n1548), .A2(n1547), .ZN(n1549) );
  MOAI22D1BWP30P140LVT U1695 ( .A1(n1616), .A2(n1547), .B1(n4), .B2(n1549), 
        .ZN(n1129) );
  INVD1BWP30P140LVT U1696 ( .I(n1550), .ZN(n1551) );
  AOI21D1BWP30P140LVT U1697 ( .A1(n1553), .A2(n1552), .B(n1551), .ZN(n1558) );
  INVD1BWP30P140LVT U1698 ( .I(n1554), .ZN(n1556) );
  XOR2UD1BWP30P140LVT U1699 ( .A1(n1558), .A2(n1557), .Z(n1958) );
  AOI21D1BWP30P140LVT U1700 ( .A1(n1813), .A2(delay_matrix_N_1_next[47]), .B(
        n1807), .ZN(n1559) );
  OAI21D1BWP30P140LVT U1701 ( .A1(n1692), .A2(n1813), .B(n1559), .ZN(n1078) );
  AOI21D1BWP30P140LVT U1702 ( .A1(n1817), .A2(delay_matrix_N_1_next[33]), .B(
        n1807), .ZN(n1560) );
  OAI21D1BWP30P140LVT U1703 ( .A1(n1692), .A2(n1817), .B(n1560), .ZN(n1064) );
  AOI21D1BWP30P140LVT U1704 ( .A1(n1815), .A2(delay_matrix_N_1_next[5]), .B(
        n1807), .ZN(n1561) );
  OAI21D1BWP30P140LVT U1705 ( .A1(n1692), .A2(n1815), .B(n1561), .ZN(n1042) );
  AOI21D1BWP30P140LVT U1706 ( .A1(n1819), .A2(delay_matrix_N_1_next[19]), .B(
        n1807), .ZN(n1562) );
  OAI21D1BWP30P140LVT U1707 ( .A1(n1692), .A2(n1819), .B(n1562), .ZN(n1028) );
  AOI21D1BWP30P140LVT U1708 ( .A1(n561), .A2(delay_matrix_N_1_next[8]), .B(
        n1807), .ZN(n1564) );
  OAI211D1BWP30P140LVT U1709 ( .A1(n1565), .A2(n2181), .B(n1564), .C(n1563), 
        .ZN(n1011) );
  AOI21D1BWP30P140LVT U1710 ( .A1(n1333), .A2(
        delay_matrix_N_1_next_original[46]), .B(n1807), .ZN(n1566) );
  OAI21D1BWP30P140LVT U1711 ( .A1(n1790), .A2(n1333), .B(n1566), .ZN(n919) );
  AOI21D1BWP30P140LVT U1712 ( .A1(n1333), .A2(
        delay_matrix_N_1_next_original[50]), .B(n1807), .ZN(n1567) );
  OAI21D1BWP30P140LVT U1713 ( .A1(n1776), .A2(n1333), .B(n1567), .ZN(n915) );
  AOI21D1BWP30P140LVT U1714 ( .A1(n1333), .A2(
        delay_matrix_N_1_next_original[42]), .B(n1807), .ZN(n1568) );
  OAI21D1BWP30P140LVT U1715 ( .A1(n1793), .A2(n1333), .B(n1568), .ZN(n923) );
  AOI21D1BWP30P140LVT U1716 ( .A1(n1333), .A2(
        delay_matrix_N_1_next_original[44]), .B(n1807), .ZN(n1569) );
  OAI21D1BWP30P140LVT U1717 ( .A1(n1810), .A2(n1333), .B(n1569), .ZN(n921) );
  AOI21D1BWP30P140LVT U1718 ( .A1(n1333), .A2(
        delay_matrix_N_1_next_original[47]), .B(n1807), .ZN(n1570) );
  OAI21D1BWP30P140LVT U1719 ( .A1(n1798), .A2(n1333), .B(n1570), .ZN(n918) );
  AOI21D1BWP30P140LVT U1720 ( .A1(n1333), .A2(
        delay_matrix_N_1_next_original[48]), .B(n1807), .ZN(n1571) );
  OAI21D1BWP30P140LVT U1721 ( .A1(n1805), .A2(n1333), .B(n1571), .ZN(n917) );
  XNR2UD1BWP30P140LVT U1722 ( .A1(n1573), .A2(n1572), .ZN(n1574) );
  MOAI22D1BWP30P140LVT U1723 ( .A1(n1616), .A2(n1572), .B1(n4), .B2(n1574), 
        .ZN(n1135) );
  ND2D1BWP30P140LVT U1724 ( .A1(n1614), .A2(copy_pointer[8]), .ZN(n1576) );
  INVD1BWP30P140LVT U1725 ( .I(copy_pointer[9]), .ZN(n1575) );
  XOR2UD1BWP30P140LVT U1726 ( .A1(n1576), .A2(n1575), .Z(n1577) );
  MOAI22D1BWP30P140LVT U1727 ( .A1(n1616), .A2(n1575), .B1(n4), .B2(n1577), 
        .ZN(n1138) );
  INVD1BWP30P140LVT U1728 ( .I(copy_pointer[6]), .ZN(n1578) );
  XNR2UD1BWP30P140LVT U1729 ( .A1(n1579), .A2(n1578), .ZN(n1580) );
  MOAI22D1BWP30P140LVT U1730 ( .A1(n1616), .A2(n1578), .B1(n4), .B2(n1580), 
        .ZN(n1141) );
  INVD1BWP30P140LVT U1731 ( .I(copy_pointer[22]), .ZN(n1581) );
  XNR2UD1BWP30P140LVT U1732 ( .A1(n1582), .A2(n1581), .ZN(n1583) );
  MOAI22D1BWP30P140LVT U1733 ( .A1(n1616), .A2(n1581), .B1(n4), .B2(n1583), 
        .ZN(n1125) );
  INVD1BWP30P140LVT U1734 ( .I(n1584), .ZN(n1749) );
  AOI21D1BWP30P140LVT U1735 ( .A1(n1749), .A2(n1748), .B(n1585), .ZN(n1589) );
  OAI22D1BWP30P140LVT U1736 ( .A1(n1587), .A2(n2191), .B1(n1586), .B2(n5), 
        .ZN(n1588) );
  AOI21D1BWP30P140LVT U1737 ( .A1(n1589), .A2(n1245), .B(n1588), .ZN(n1591) );
  NR2D1BWP30P140LVT U1738 ( .A1(n1593), .A2(n1592), .ZN(n1595) );
  INVD1BWP30P140LVT U1739 ( .I(copy_pointer[5]), .ZN(n1594) );
  XNR2UD1BWP30P140LVT U1740 ( .A1(n1595), .A2(n1594), .ZN(n1596) );
  MOAI22D1BWP30P140LVT U1741 ( .A1(n1616), .A2(n1594), .B1(n4), .B2(n1596), 
        .ZN(n1142) );
  INVD1BWP30P140LVT U1742 ( .I(copy_pointer[29]), .ZN(n1599) );
  HA1D1BWP30P140LVT U1743 ( .A(copy_pointer[29]), .B(n1597), .CO(n1836), .S(
        n1598) );
  MOAI22D1BWP30P140LVT U1744 ( .A1(n1616), .A2(n1599), .B1(n4), .B2(n1598), 
        .ZN(n1118) );
  INVD1BWP30P140LVT U1745 ( .I(copy_pointer[28]), .ZN(n1602) );
  HA1D1BWP30P140LVT U1746 ( .A(copy_pointer[28]), .B(n1600), .CO(n1597), .S(
        n1601) );
  MOAI22D1BWP30P140LVT U1747 ( .A1(n1616), .A2(n1602), .B1(n4), .B2(n1601), 
        .ZN(n1119) );
  NR2D1BWP30P140LVT U1748 ( .A1(n1604), .A2(n1603), .ZN(n1606) );
  INVD1BWP30P140LVT U1749 ( .I(copy_pointer[15]), .ZN(n1605) );
  XNR2UD1BWP30P140LVT U1750 ( .A1(n1606), .A2(n1605), .ZN(n1607) );
  MOAI22D1BWP30P140LVT U1751 ( .A1(n1616), .A2(n1605), .B1(n4), .B2(n1607), 
        .ZN(n1132) );
  NR2D1BWP30P140LVT U1752 ( .A1(n1609), .A2(n1608), .ZN(n1611) );
  INVD1BWP30P140LVT U1753 ( .I(copy_pointer[11]), .ZN(n1610) );
  XNR2UD1BWP30P140LVT U1754 ( .A1(n1611), .A2(n1610), .ZN(n1612) );
  MOAI22D1BWP30P140LVT U1755 ( .A1(n1616), .A2(n1610), .B1(n4), .B2(n1612), 
        .ZN(n1136) );
  INVD1BWP30P140LVT U1756 ( .I(copy_pointer[8]), .ZN(n1613) );
  XNR2UD1BWP30P140LVT U1757 ( .A1(n1614), .A2(n1613), .ZN(n1615) );
  MOAI22D1BWP30P140LVT U1758 ( .A1(n1616), .A2(n1613), .B1(n4), .B2(n1615), 
        .ZN(n1139) );
  MUX2NUD1BWP30P140LVT U1759 ( .I0(n1638), .I1(delay_matrix_N_1_next[53]), .S(
        n1813), .ZN(n1617) );
  MUX2NUD1BWP30P140LVT U1760 ( .I0(n1638), .I1(delay_matrix_N_1_next[25]), .S(
        n1819), .ZN(n1618) );
  INVD1BWP30P140LVT U1761 ( .I(copy_ptr_next[1]), .ZN(n1619) );
  XNR2UD1BWP30P140LVT U1762 ( .A1(n1619), .A2(copy_ptr_next[0]), .ZN(n1620) );
  MOAI22D1BWP30P140LVT U1763 ( .A1(n1835), .A2(n1619), .B1(n1620), .B2(n6), 
        .ZN(n954) );
  ND2OPTIBD1BWP30P140LVT U1764 ( .A1(n1820), .A2(n1982), .ZN(n1622) );
  AOI21D1BWP30P140LVT U1765 ( .A1(n561), .A2(delay_matrix_N_1_next[51]), .B(
        n1807), .ZN(n1621) );
  OAI211D1BWP30P140LVT U1766 ( .A1(n1988), .A2(n1623), .B(n1622), .C(n1621), 
        .ZN(n968) );
  MUX2NUD1BWP30P140LVT U1767 ( .I0(n1638), .I1(delay_matrix_N_1_next[11]), .S(
        n1815), .ZN(n1624) );
  AOI21D1BWP30P140LVT U1768 ( .A1(n561), .A2(delay_matrix_N_1_next[1]), .B(
        n1807), .ZN(n1626) );
  OAI211D1BWP30P140LVT U1769 ( .A1(n1627), .A2(n2181), .B(n1626), .C(n1625), 
        .ZN(n1018) );
  INVD1BWP30P140LVT U1770 ( .I(n1638), .ZN(n1630) );
  AOI21D1BWP30P140LVT U1771 ( .A1(n561), .A2(delay_matrix_N_1_next[11]), .B(
        n1807), .ZN(n1629) );
  OAI211D1BWP30P140LVT U1772 ( .A1(n1630), .A2(n2181), .B(n1629), .C(n1628), 
        .ZN(n1008) );
  INVD1BWP30P140LVT U1773 ( .I(n1631), .ZN(n1634) );
  AOI21D1BWP30P140LVT U1774 ( .A1(n561), .A2(delay_matrix_N_1_next[10]), .B(
        n1807), .ZN(n1633) );
  OAI211D1BWP30P140LVT U1775 ( .A1(n1634), .A2(n2181), .B(n1633), .C(n1632), 
        .ZN(n1009) );
  AOI21D1BWP30P140LVT U1776 ( .A1(n561), .A2(delay_matrix_N_1_next[6]), .B(
        n1807), .ZN(n1636) );
  OAI211D1BWP30P140LVT U1777 ( .A1(n1637), .A2(n2181), .B(n1636), .C(n1635), 
        .ZN(n1013) );
  MUX2NUD1BWP30P140LVT U1778 ( .I0(n1638), .I1(delay_matrix_N_1_next[39]), .S(
        n1817), .ZN(n1639) );
  AOI21D1BWP30P140LVT U1779 ( .A1(n561), .A2(
        delay_matrix_N_1_next_original[31]), .B(n1807), .ZN(n1640) );
  OAI211D1BWP30P140LVT U1780 ( .A1(n2207), .A2(n1678), .B(n1641), .C(n1640), 
        .ZN(n836) );
  AOI21D1BWP30P140LVT U1781 ( .A1(n561), .A2(
        delay_matrix_N_1_next_original[43]), .B(n1807), .ZN(n1642) );
  OAI211D1BWP30P140LVT U1782 ( .A1(n1806), .A2(n1665), .B(n1643), .C(n1642), 
        .ZN(n824) );
  AOI21D1BWP30P140LVT U1783 ( .A1(n561), .A2(delay_matrix_N_1_next[0]), .B(
        n1807), .ZN(n1644) );
  OAI211D1BWP30P140LVT U1784 ( .A1(n1646), .A2(n2181), .B(n1645), .C(n1644), 
        .ZN(n1019) );
  AOI21D1BWP30P140LVT U1785 ( .A1(scenario_update), .A2(
        delay_matrix_N_1_next_original[4]), .B(n1807), .ZN(n1647) );
  OAI211D1BWP30P140LVT U1786 ( .A1(n1790), .A2(n2196), .B(n1648), .C(n1647), 
        .ZN(n863) );
  AOI21D1BWP30P140LVT U1787 ( .A1(n1802), .A2(
        delay_matrix_N_1_next_original[7]), .B(n1807), .ZN(n1649) );
  OAI211D1BWP30P140LVT U1788 ( .A1(n1779), .A2(n2196), .B(n1650), .C(n1649), 
        .ZN(n860) );
  AOI21D1BWP30P140LVT U1789 ( .A1(n1802), .A2(
        delay_matrix_N_1_next_original[34]), .B(n1807), .ZN(n1651) );
  OAI211D1BWP30P140LVT U1790 ( .A1(n2207), .A2(n1805), .B(n1652), .C(n1651), 
        .ZN(n833) );
  AOI21D1BWP30P140LVT U1791 ( .A1(n561), .A2(
        delay_matrix_N_1_next_original[17]), .B(n1807), .ZN(n1653) );
  OAI211D1BWP30P140LVT U1792 ( .A1(n2202), .A2(n1678), .B(n1654), .C(n1653), 
        .ZN(n850) );
  AOI21D1BWP30P140LVT U1793 ( .A1(n561), .A2(delay_matrix_N_1_next_original[1]), .B(n1807), .ZN(n1655) );
  OAI211D1BWP30P140LVT U1794 ( .A1(n1665), .A2(n2196), .B(n1656), .C(n1655), 
        .ZN(n866) );
  AOI21D1BWP30P140LVT U1795 ( .A1(n1773), .A2(
        delay_matrix_N_1_next_original[35]), .B(n1807), .ZN(n1657) );
  OAI211D1BWP30P140LVT U1796 ( .A1(n2207), .A2(n1779), .B(n1658), .C(n1657), 
        .ZN(n832) );
  AOI21D1BWP30P140LVT U1797 ( .A1(n561), .A2(
        delay_matrix_N_1_next_original[45]), .B(n1807), .ZN(n1659) );
  OAI211D1BWP30P140LVT U1798 ( .A1(n1678), .A2(n1806), .B(n1660), .C(n1659), 
        .ZN(n822) );
  AOI21D1BWP30P140LVT U1799 ( .A1(n561), .A2(
        delay_matrix_N_1_next_original[29]), .B(n1807), .ZN(n1661) );
  OAI211D1BWP30P140LVT U1800 ( .A1(n2207), .A2(n1665), .B(n1662), .C(n1661), 
        .ZN(n838) );
  AOI21D1BWP30P140LVT U1801 ( .A1(n561), .A2(
        delay_matrix_N_1_next_original[15]), .B(n1807), .ZN(n1663) );
  OAI211D1BWP30P140LVT U1802 ( .A1(n2202), .A2(n1665), .B(n1664), .C(n1663), 
        .ZN(n852) );
  AOI21D1BWP30P140LVT U1803 ( .A1(n561), .A2(
        delay_matrix_N_1_next_original[28]), .B(n1807), .ZN(n1666) );
  OAI211D1BWP30P140LVT U1804 ( .A1(n2207), .A2(n1793), .B(n1667), .C(n1666), 
        .ZN(n839) );
  AOI21D1BWP30P140LVT U1805 ( .A1(n1773), .A2(
        delay_matrix_N_1_next_original[50]), .B(n1807), .ZN(n1668) );
  OAI211D1BWP30P140LVT U1806 ( .A1(n1806), .A2(n1776), .B(n1669), .C(n1668), 
        .ZN(n817) );
  AOI21D1BWP30P140LVT U1807 ( .A1(n1802), .A2(
        delay_matrix_N_1_next_original[20]), .B(n1807), .ZN(n1670) );
  OAI211D1BWP30P140LVT U1808 ( .A1(n2202), .A2(n1805), .B(n1671), .C(n1670), 
        .ZN(n847) );
  AOI21D1BWP30P140LVT U1809 ( .A1(n1802), .A2(
        delay_matrix_N_1_next_original[46]), .B(n1807), .ZN(n1672) );
  OAI211D1BWP30P140LVT U1810 ( .A1(n1806), .A2(n1790), .B(n1673), .C(n1672), 
        .ZN(n821) );
  AOI21D1BWP30P140LVT U1811 ( .A1(n1802), .A2(
        delay_matrix_N_1_next_original[21]), .B(n1807), .ZN(n1674) );
  OAI211D1BWP30P140LVT U1812 ( .A1(n2202), .A2(n1779), .B(n1675), .C(n1674), 
        .ZN(n846) );
  AOI21D1BWP30P140LVT U1813 ( .A1(scenario_update), .A2(
        delay_matrix_N_1_next_original[3]), .B(n1807), .ZN(n1676) );
  OAI211D1BWP30P140LVT U1814 ( .A1(n1678), .A2(n2196), .B(n1677), .C(n1676), 
        .ZN(n864) );
  INVD1BWP30P140LVT U1815 ( .I(ptr_next[26]), .ZN(n1680) );
  MOAI22D1BWP30P140LVT U1816 ( .A1(n1680), .A2(n1835), .B1(n6), .B2(n1679), 
        .ZN(n1089) );
  NR2D1BWP30P140LVT U1817 ( .A1(n1727), .A2(n1682), .ZN(n1904) );
  INVD1BWP30P140LVT U1818 ( .I(ptr_next[24]), .ZN(n1683) );
  XNR2UD1BWP30P140LVT U1819 ( .A1(n1904), .A2(n1683), .ZN(n1684) );
  MOAI22D1BWP30P140LVT U1820 ( .A1(n1683), .A2(n1835), .B1(n6), .B2(n1684), 
        .ZN(n1091) );
  INVD1BWP30P140LVT U1821 ( .I(n1685), .ZN(n1686) );
  NR2D1BWP30P140LVT U1822 ( .A1(n1727), .A2(n1686), .ZN(n1697) );
  INVD1BWP30P140LVT U1823 ( .I(n1697), .ZN(n1708) );
  NR2D1BWP30P140LVT U1824 ( .A1(n1708), .A2(n1687), .ZN(n1894) );
  INVD1BWP30P140LVT U1825 ( .I(ptr_next[22]), .ZN(n1688) );
  XNR2UD1BWP30P140LVT U1826 ( .A1(n1894), .A2(n1688), .ZN(n1689) );
  MOAI22D1BWP30P140LVT U1827 ( .A1(n1688), .A2(n1835), .B1(n6), .B2(n1689), 
        .ZN(n1093) );
  AOI21D1BWP30P140LVT U1828 ( .A1(n561), .A2(delay_matrix_N_1_next[5]), .B(
        n1807), .ZN(n1691) );
  OAI211D1BWP30P140LVT U1829 ( .A1(n1692), .A2(n2181), .B(n1691), .C(n1690), 
        .ZN(n1014) );
  NR2D1BWP30P140LVT U1830 ( .A1(n1727), .A2(n1693), .ZN(n1721) );
  INVD1BWP30P140LVT U1831 ( .I(ptr_next[19]), .ZN(n1694) );
  XOR2UD1BWP30P140LVT U1832 ( .A1(n1695), .A2(n1694), .Z(n1696) );
  MOAI22D1BWP30P140LVT U1833 ( .A1(n1694), .A2(n1835), .B1(n6), .B2(n1696), 
        .ZN(n1096) );
  INVD1BWP30P140LVT U1834 ( .I(ptr_next[21]), .ZN(n1698) );
  XOR2UD1BWP30P140LVT U1835 ( .A1(n1699), .A2(n1698), .Z(n1700) );
  MOAI22D1BWP30P140LVT U1836 ( .A1(n1698), .A2(n1835), .B1(n6), .B2(n1700), 
        .ZN(n1094) );
  INVD1BWP30P140LVT U1837 ( .I(ptr_next[8]), .ZN(n1702) );
  XNR2UD1BWP30P140LVT U1838 ( .A1(n1716), .A2(n1702), .ZN(n1703) );
  MOAI22D1BWP30P140LVT U1839 ( .A1(n1702), .A2(n1835), .B1(n6), .B2(n1703), 
        .ZN(n1107) );
  INVD1BWP30P140LVT U1840 ( .I(ptr_next[9]), .ZN(n1704) );
  XOR2UD1BWP30P140LVT U1841 ( .A1(n1705), .A2(n1704), .Z(n1706) );
  MOAI22D1BWP30P140LVT U1842 ( .A1(n1704), .A2(n1835), .B1(n6), .B2(n1706), 
        .ZN(n1106) );
  INVD1BWP30P140LVT U1843 ( .I(ptr_next[20]), .ZN(n1707) );
  XOR2UD1BWP30P140LVT U1844 ( .A1(n1708), .A2(n1707), .Z(n1709) );
  MOAI22D1BWP30P140LVT U1845 ( .A1(n1707), .A2(n1835), .B1(n6), .B2(n1709), 
        .ZN(n1095) );
  INVD1BWP30P140LVT U1846 ( .I(n1729), .ZN(n1737) );
  INVD1BWP30P140LVT U1847 ( .I(n1711), .ZN(n1712) );
  ND2D1BWP30P140LVT U1848 ( .A1(n1737), .A2(n1712), .ZN(n1740) );
  INVD1BWP30P140LVT U1849 ( .I(ptr_next[14]), .ZN(n1739) );
  XOR2UD1BWP30P140LVT U1850 ( .A1(n1740), .A2(n1739), .Z(n1713) );
  MOAI22D1BWP30P140LVT U1851 ( .A1(n1739), .A2(n1835), .B1(n6), .B2(n1713), 
        .ZN(n1101) );
  INVD1BWP30P140LVT U1852 ( .I(n1714), .ZN(n1715) );
  ND2D1BWP30P140LVT U1853 ( .A1(n1716), .A2(n1715), .ZN(n1734) );
  INVD1BWP30P140LVT U1854 ( .I(ptr_next[10]), .ZN(n1733) );
  NR2D1BWP30P140LVT U1855 ( .A1(n1734), .A2(n1733), .ZN(n1718) );
  INVD1BWP30P140LVT U1856 ( .I(ptr_next[11]), .ZN(n1717) );
  XNR2UD1BWP30P140LVT U1857 ( .A1(n1718), .A2(n1717), .ZN(n1719) );
  MOAI22D1BWP30P140LVT U1858 ( .A1(n1717), .A2(n1835), .B1(n6), .B2(n1719), 
        .ZN(n1104) );
  INVD1BWP30P140LVT U1859 ( .I(ptr_next[18]), .ZN(n1720) );
  XNR2UD1BWP30P140LVT U1860 ( .A1(n1721), .A2(n1720), .ZN(n1722) );
  MOAI22D1BWP30P140LVT U1861 ( .A1(n1720), .A2(n1835), .B1(n6), .B2(n1722), 
        .ZN(n1097) );
  INVD1BWP30P140LVT U1862 ( .I(ptr_next[16]), .ZN(n1726) );
  NR2D1BWP30P140LVT U1863 ( .A1(n1727), .A2(n1726), .ZN(n1724) );
  INVD1BWP30P140LVT U1864 ( .I(ptr_next[17]), .ZN(n1723) );
  XNR2UD1BWP30P140LVT U1865 ( .A1(n1724), .A2(n1723), .ZN(n1725) );
  MOAI22D1BWP30P140LVT U1866 ( .A1(n1723), .A2(n1835), .B1(n6), .B2(n1725), 
        .ZN(n1098) );
  XOR2UD1BWP30P140LVT U1867 ( .A1(n1727), .A2(n1726), .Z(n1728) );
  MOAI22D1BWP30P140LVT U1868 ( .A1(n1726), .A2(n1835), .B1(n6), .B2(n1728), 
        .ZN(n1099) );
  INVD1BWP30P140LVT U1869 ( .I(ptr_next[12]), .ZN(n1736) );
  NR2D1BWP30P140LVT U1870 ( .A1(n1729), .A2(n1736), .ZN(n1731) );
  INVD1BWP30P140LVT U1871 ( .I(ptr_next[13]), .ZN(n1730) );
  XNR2UD1BWP30P140LVT U1872 ( .A1(n1731), .A2(n1730), .ZN(n1732) );
  MOAI22D1BWP30P140LVT U1873 ( .A1(n1730), .A2(n1835), .B1(n6), .B2(n1732), 
        .ZN(n1102) );
  XOR2UD1BWP30P140LVT U1874 ( .A1(n1734), .A2(n1733), .Z(n1735) );
  MOAI22D1BWP30P140LVT U1875 ( .A1(n1733), .A2(n1835), .B1(n6), .B2(n1735), 
        .ZN(n1105) );
  XNR2UD1BWP30P140LVT U1876 ( .A1(n1737), .A2(n1736), .ZN(n1738) );
  MOAI22D1BWP30P140LVT U1877 ( .A1(n1736), .A2(n1835), .B1(n6), .B2(n1738), 
        .ZN(n1103) );
  NR2D1BWP30P140LVT U1878 ( .A1(n1740), .A2(n1739), .ZN(n1742) );
  INVD1BWP30P140LVT U1879 ( .I(ptr_next[15]), .ZN(n1741) );
  XNR2UD1BWP30P140LVT U1880 ( .A1(n1742), .A2(n1741), .ZN(n1743) );
  MOAI22D1BWP30P140LVT U1881 ( .A1(n1741), .A2(n1835), .B1(n6), .B2(n1743), 
        .ZN(n1100) );
  INVD1BWP30P140LVT U1882 ( .I(n1983), .ZN(n1746) );
  AOI21D1BWP30P140LVT U1883 ( .A1(n561), .A2(delay_matrix_N_1_next[7]), .B(
        n1807), .ZN(n1745) );
  OAI211D1BWP30P140LVT U1884 ( .A1(n1746), .A2(n2181), .B(n1745), .C(n1744), 
        .ZN(n1012) );
  AOI21D1BWP30P140LVT U1885 ( .A1(n1749), .A2(n1748), .B(n1747), .ZN(n1750) );
  OAI21D1BWP30P140LVT U1886 ( .A1(n4), .A2(n1245), .B(n1750), .ZN(n1755) );
  IAO21D1BWP30P140LVT U1887 ( .A1(n1753), .A2(n5), .B(n1752), .ZN(n1754) );
  MUX2NUD1BWP30P140LVT U1888 ( .I0(n1983), .I1(delay_matrix_N_1_next[49]), .S(
        n1813), .ZN(n1756) );
  INVD1BWP30P140LVT U1889 ( .I(n1820), .ZN(n1759) );
  AOI21D1BWP30P140LVT U1890 ( .A1(n561), .A2(delay_matrix_N_1_next[9]), .B(
        n1807), .ZN(n1758) );
  OAI211D1BWP30P140LVT U1891 ( .A1(n1759), .A2(n2181), .B(n1758), .C(n1757), 
        .ZN(n1010) );
  MUX2NUD1BWP30P140LVT U1892 ( .I0(n1983), .I1(delay_matrix_N_1_next[7]), .S(
        n1815), .ZN(n1761) );
  AOI21D1BWP30P140LVT U1893 ( .A1(scenario_update), .A2(
        delay_matrix_N_1_next_original[14]), .B(n1807), .ZN(n1764) );
  OAI211D1BWP30P140LVT U1894 ( .A1(n1766), .A2(n1765), .B(n1764), .C(n1763), 
        .ZN(n853) );
  AOI21D1BWP30P140LVT U1895 ( .A1(n1802), .A2(
        delay_matrix_N_1_next_original[32]), .B(n1807), .ZN(n1767) );
  OAI211D1BWP30P140LVT U1896 ( .A1(n2207), .A2(n1790), .B(n1768), .C(n1767), 
        .ZN(n835) );
  AOI21D1BWP30P140LVT U1897 ( .A1(n561), .A2(delay_matrix_N_1_next_original[0]), .B(n1807), .ZN(n1769) );
  OAI211D1BWP30P140LVT U1898 ( .A1(n1793), .A2(n2196), .B(n1770), .C(n1769), 
        .ZN(n867) );
  AOI21D1BWP30P140LVT U1899 ( .A1(scenario_update), .A2(
        delay_matrix_N_1_next_original[2]), .B(n1807), .ZN(n1771) );
  OAI211D1BWP30P140LVT U1900 ( .A1(n1810), .A2(n2196), .B(n1772), .C(n1771), 
        .ZN(n865) );
  AOI21D1BWP30P140LVT U1901 ( .A1(n1773), .A2(
        delay_matrix_N_1_next_original[36]), .B(n1807), .ZN(n1774) );
  OAI211D1BWP30P140LVT U1902 ( .A1(n2207), .A2(n1776), .B(n1775), .C(n1774), 
        .ZN(n831) );
  AOI21D1BWP30P140LVT U1903 ( .A1(n1802), .A2(
        delay_matrix_N_1_next_original[49]), .B(n1807), .ZN(n1777) );
  OAI211D1BWP30P140LVT U1904 ( .A1(n1806), .A2(n1779), .B(n1778), .C(n1777), 
        .ZN(n818) );
  AOI21D1BWP30P140LVT U1905 ( .A1(n561), .A2(
        delay_matrix_N_1_next_original[44]), .B(n1807), .ZN(n1780) );
  OAI211D1BWP30P140LVT U1906 ( .A1(n1806), .A2(n1810), .B(n1781), .C(n1780), 
        .ZN(n823) );
  AOI21D1BWP30P140LVT U1907 ( .A1(n1802), .A2(
        delay_matrix_N_1_next_original[5]), .B(n1807), .ZN(n1782) );
  OAI211D1BWP30P140LVT U1908 ( .A1(n1798), .A2(n2196), .B(n1783), .C(n1782), 
        .ZN(n862) );
  AOI21D1BWP30P140LVT U1909 ( .A1(n1802), .A2(
        delay_matrix_N_1_next_original[19]), .B(n1807), .ZN(n1784) );
  OAI211D1BWP30P140LVT U1910 ( .A1(n2202), .A2(n1798), .B(n1785), .C(n1784), 
        .ZN(n848) );
  AOI21D1BWP30P140LVT U1911 ( .A1(n1802), .A2(
        delay_matrix_N_1_next_original[33]), .B(n1807), .ZN(n1786) );
  OAI211D1BWP30P140LVT U1912 ( .A1(n2207), .A2(n1798), .B(n1787), .C(n1786), 
        .ZN(n834) );
  AOI21D1BWP30P140LVT U1913 ( .A1(n1802), .A2(
        delay_matrix_N_1_next_original[18]), .B(n1807), .ZN(n1788) );
  OAI211D1BWP30P140LVT U1914 ( .A1(n2202), .A2(n1790), .B(n1789), .C(n1788), 
        .ZN(n849) );
  AOI21D1BWP30P140LVT U1915 ( .A1(n561), .A2(
        delay_matrix_N_1_next_original[42]), .B(n1807), .ZN(n1791) );
  OAI211D1BWP30P140LVT U1916 ( .A1(n1806), .A2(n1793), .B(n1792), .C(n1791), 
        .ZN(n825) );
  AOI21D1BWP30P140LVT U1917 ( .A1(scenario_update), .A2(
        delay_matrix_N_1_next_original[6]), .B(n1807), .ZN(n1794) );
  OAI211D1BWP30P140LVT U1918 ( .A1(n1805), .A2(n2196), .B(n1795), .C(n1794), 
        .ZN(n861) );
  AOI21D1BWP30P140LVT U1919 ( .A1(n1802), .A2(
        delay_matrix_N_1_next_original[47]), .B(n1807), .ZN(n1796) );
  OAI211D1BWP30P140LVT U1920 ( .A1(n1806), .A2(n1798), .B(n1797), .C(n1796), 
        .ZN(n820) );
  AOI21D1BWP30P140LVT U1921 ( .A1(n561), .A2(
        delay_matrix_N_1_next_original[16]), .B(n1807), .ZN(n1799) );
  OAI211D1BWP30P140LVT U1922 ( .A1(n2202), .A2(n1810), .B(n1800), .C(n1799), 
        .ZN(n851) );
  AOI21D1BWP30P140LVT U1923 ( .A1(n1802), .A2(
        delay_matrix_N_1_next_original[48]), .B(n1807), .ZN(n1803) );
  OAI211D1BWP30P140LVT U1924 ( .A1(n1806), .A2(n1805), .B(n1804), .C(n1803), 
        .ZN(n819) );
  AOI21D1BWP30P140LVT U1925 ( .A1(n561), .A2(
        delay_matrix_N_1_next_original[30]), .B(n1807), .ZN(n1808) );
  OAI211D1BWP30P140LVT U1926 ( .A1(n2207), .A2(n1810), .B(n1809), .C(n1808), 
        .ZN(n837) );
  MUX2NUD1BWP30P140LVT U1927 ( .I0(n1983), .I1(delay_matrix_N_1_next[35]), .S(
        n1817), .ZN(n1811) );
  MUX2NUD1BWP30P140LVT U1928 ( .I0(n1983), .I1(delay_matrix_N_1_next[21]), .S(
        n1819), .ZN(n1812) );
  MUX2NUD1BWP30P140LVT U1929 ( .I0(n1820), .I1(delay_matrix_N_1_next[51]), .S(
        n1813), .ZN(n1814) );
  MUX2NUD1BWP30P140LVT U1930 ( .I0(n1820), .I1(delay_matrix_N_1_next[9]), .S(
        n1815), .ZN(n1816) );
  MUX2NUD1BWP30P140LVT U1931 ( .I0(n1820), .I1(delay_matrix_N_1_next[37]), .S(
        n1817), .ZN(n1818) );
  MUX2NUD1BWP30P140LVT U1932 ( .I0(n1820), .I1(delay_matrix_N_1_next[23]), .S(
        n1819), .ZN(n1822) );
  XNR2UD1BWP30P140LVT U1933 ( .A1(n1824), .A2(ptr_next[0]), .ZN(n1823) );
  MOAI22D1BWP30P140LVT U1934 ( .A1(n1824), .A2(n1835), .B1(n1823), .B2(n6), 
        .ZN(n1114) );
  INVD1BWP30P140LVT U1935 ( .I(n1825), .ZN(n1830) );
  ND2D1BWP30P140LVT U1936 ( .A1(n1830), .A2(ptr_next[2]), .ZN(n1827) );
  INVD1BWP30P140LVT U1937 ( .I(ptr_next[3]), .ZN(n1826) );
  XOR2UD1BWP30P140LVT U1938 ( .A1(n1827), .A2(n1826), .Z(n1828) );
  MOAI22D1BWP30P140LVT U1939 ( .A1(n1826), .A2(n1835), .B1(n6), .B2(n1828), 
        .ZN(n1112) );
  INVD1BWP30P140LVT U1940 ( .I(ptr_next[2]), .ZN(n1829) );
  XNR2UD1BWP30P140LVT U1941 ( .A1(n1830), .A2(n1829), .ZN(n1831) );
  MOAI22D1BWP30P140LVT U1942 ( .A1(n1829), .A2(n1835), .B1(n6), .B2(n1831), 
        .ZN(n1113) );
  XOR2UD1BWP30P140LVT U1943 ( .A1(n1833), .A2(n1832), .Z(n1834) );
  MOAI22D1BWP30P140LVT U1944 ( .A1(n1832), .A2(n1835), .B1(n6), .B2(n1834), 
        .ZN(n1111) );
  HA1D1BWP30P140LVT U1945 ( .A(copy_pointer[30]), .B(n1836), .CO(n1837), .S(
        n1506) );
  MOAI22D1BWP30P140LVT U1946 ( .A1(n1616), .A2(n1839), .B1(n4), .B2(n1838), 
        .ZN(n1116) );
  INVD1BWP30P140LVT U1947 ( .I(copy_ptr_next[30]), .ZN(n1842) );
  HA1D1BWP30P140LVT U1948 ( .A(copy_ptr_next[30]), .B(n1840), .CO(n236), .S(
        n1841) );
  MOAI22D1BWP30P140LVT U1949 ( .A1(n1835), .A2(n1842), .B1(n6), .B2(n1841), 
        .ZN(n925) );
  INVD1BWP30P140LVT U1950 ( .I(copy_ptr_next[27]), .ZN(n1845) );
  HA1D1BWP30P140LVT U1951 ( .A(copy_ptr_next[27]), .B(n1843), .CO(n1848), .S(
        n1844) );
  MOAI22D1BWP30P140LVT U1952 ( .A1(n1835), .A2(n1845), .B1(n6), .B2(n1844), 
        .ZN(n928) );
  INVD1BWP30P140LVT U1953 ( .I(copy_ptr_next[26]), .ZN(n1847) );
  HA1D1BWP30P140LVT U1954 ( .A(copy_ptr_next[26]), .B(n16), .CO(n1843), .S(
        n1846) );
  MOAI22D1BWP30P140LVT U1955 ( .A1(n1835), .A2(n1847), .B1(n6), .B2(n1846), 
        .ZN(n929) );
  INVD1BWP30P140LVT U1956 ( .I(copy_ptr_next[28]), .ZN(n1850) );
  HA1D1BWP30P140LVT U1957 ( .A(copy_ptr_next[28]), .B(n1848), .CO(n1855), .S(
        n1849) );
  MOAI22D1BWP30P140LVT U1958 ( .A1(n1835), .A2(n1850), .B1(n6), .B2(n1849), 
        .ZN(n927) );
  NR2D1BWP30P140LVT U1959 ( .A1(n1890), .A2(n1851), .ZN(n1859) );
  INVD1BWP30P140LVT U1960 ( .I(copy_ptr_next[25]), .ZN(n1852) );
  XOR2UD1BWP30P140LVT U1961 ( .A1(n1853), .A2(n1852), .Z(n1854) );
  MOAI22D1BWP30P140LVT U1962 ( .A1(n1835), .A2(n1852), .B1(n6), .B2(n1854), 
        .ZN(n930) );
  INVD1BWP30P140LVT U1963 ( .I(copy_ptr_next[29]), .ZN(n1857) );
  HA1D1BWP30P140LVT U1964 ( .A(copy_ptr_next[29]), .B(n1855), .CO(n1840), .S(
        n1856) );
  MOAI22D1BWP30P140LVT U1965 ( .A1(n1835), .A2(n1857), .B1(n6), .B2(n1856), 
        .ZN(n926) );
  INVD1BWP30P140LVT U1966 ( .I(copy_ptr_next[24]), .ZN(n1858) );
  XNR2UD1BWP30P140LVT U1967 ( .A1(n1859), .A2(n1858), .ZN(n1860) );
  MOAI22D1BWP30P140LVT U1968 ( .A1(n1835), .A2(n1858), .B1(n6), .B2(n1860), 
        .ZN(n931) );
  INVD1BWP30P140LVT U1969 ( .I(n1861), .ZN(n1862) );
  NR2D1BWP30P140LVT U1970 ( .A1(n1890), .A2(n1862), .ZN(n1873) );
  INVD1BWP30P140LVT U1971 ( .I(n1873), .ZN(n1866) );
  INVD1BWP30P140LVT U1972 ( .I(copy_ptr_next[20]), .ZN(n1863) );
  XOR2UD1BWP30P140LVT U1973 ( .A1(n1866), .A2(n1863), .Z(n1864) );
  MOAI22D1BWP30P140LVT U1974 ( .A1(n1835), .A2(n1863), .B1(n6), .B2(n1864), 
        .ZN(n935) );
  NR2D1BWP30P140LVT U1975 ( .A1(n1866), .A2(n1865), .ZN(n1871) );
  INVD1BWP30P140LVT U1976 ( .I(copy_ptr_next[23]), .ZN(n1867) );
  XOR2UD1BWP30P140LVT U1977 ( .A1(n1868), .A2(n1867), .Z(n1869) );
  MOAI22D1BWP30P140LVT U1978 ( .A1(n1835), .A2(n1867), .B1(n6), .B2(n1869), 
        .ZN(n932) );
  INVD1BWP30P140LVT U1979 ( .I(copy_ptr_next[22]), .ZN(n1870) );
  XNR2UD1BWP30P140LVT U1980 ( .A1(n1871), .A2(n1870), .ZN(n1872) );
  MOAI22D1BWP30P140LVT U1981 ( .A1(n1835), .A2(n1870), .B1(n6), .B2(n1872), 
        .ZN(n933) );
  INVD1BWP30P140LVT U1982 ( .I(copy_ptr_next[21]), .ZN(n1874) );
  XOR2UD1BWP30P140LVT U1983 ( .A1(n1875), .A2(n1874), .Z(n1876) );
  MOAI22D1BWP30P140LVT U1984 ( .A1(n1835), .A2(n1874), .B1(n6), .B2(n1876), 
        .ZN(n934) );
  NR2D1BWP30P140LVT U1985 ( .A1(n1890), .A2(n1877), .ZN(n1880) );
  INVD1BWP30P140LVT U1986 ( .I(copy_ptr_next[18]), .ZN(n1878) );
  XNR2UD1BWP30P140LVT U1987 ( .A1(n1880), .A2(n1878), .ZN(n1879) );
  MOAI22D1BWP30P140LVT U1988 ( .A1(n1835), .A2(n1878), .B1(n6), .B2(n1879), 
        .ZN(n937) );
  INVD1BWP30P140LVT U1989 ( .I(copy_ptr_next[19]), .ZN(n1881) );
  XOR2UD1BWP30P140LVT U1990 ( .A1(n1882), .A2(n1881), .Z(n1883) );
  MOAI22D1BWP30P140LVT U1991 ( .A1(n1835), .A2(n1881), .B1(n6), .B2(n1883), 
        .ZN(n936) );
  NR2D1BWP30P140LVT U1992 ( .A1(n1885), .A2(n1884), .ZN(n1887) );
  INVD1BWP30P140LVT U1993 ( .I(copy_ptr_next[15]), .ZN(n1886) );
  XNR2UD1BWP30P140LVT U1994 ( .A1(n1887), .A2(n1886), .ZN(n1888) );
  MOAI22D1BWP30P140LVT U1995 ( .A1(n1835), .A2(n1886), .B1(n6), .B2(n1888), 
        .ZN(n940) );
  NR2D1BWP30P140LVT U1996 ( .A1(n1890), .A2(n1889), .ZN(n1892) );
  INVD1BWP30P140LVT U1997 ( .I(copy_ptr_next[17]), .ZN(n1891) );
  XNR2UD1BWP30P140LVT U1998 ( .A1(n1892), .A2(n1891), .ZN(n1893) );
  MOAI22D1BWP30P140LVT U1999 ( .A1(n1835), .A2(n1891), .B1(n6), .B2(n1893), 
        .ZN(n938) );
  INVD1BWP30P140LVT U2000 ( .I(ptr_next[23]), .ZN(n1895) );
  XOR2UD1BWP30P140LVT U2001 ( .A1(n1896), .A2(n1895), .Z(n1897) );
  MOAI22D1BWP30P140LVT U2002 ( .A1(n1895), .A2(n1835), .B1(n6), .B2(n1897), 
        .ZN(n1092) );
  XOR2UD1BWP30P140LVT U2003 ( .A1(n1899), .A2(n1898), .Z(n1900) );
  MOAI22D1BWP30P140LVT U2004 ( .A1(n1835), .A2(n1898), .B1(n6), .B2(n1900), 
        .ZN(n951) );
  INVD1BWP30P140LVT U2005 ( .I(ptr_next[30]), .ZN(n1903) );
  MOAI22D1BWP30P140LVT U2006 ( .A1(n1903), .A2(n1835), .B1(n6), .B2(n1902), 
        .ZN(n1085) );
  INVD1BWP30P140LVT U2007 ( .I(ptr_next[25]), .ZN(n1905) );
  XOR2UD1BWP30P140LVT U2008 ( .A1(n1906), .A2(n1905), .Z(n1907) );
  MOAI22D1BWP30P140LVT U2009 ( .A1(n1905), .A2(n1835), .B1(n6), .B2(n1907), 
        .ZN(n1090) );
  INVD1BWP30P140LVT U2010 ( .I(ptr_next[27]), .ZN(n1910) );
  MOAI22D1BWP30P140LVT U2011 ( .A1(n1910), .A2(n1835), .B1(n6), .B2(n1909), 
        .ZN(n1088) );
  INVD1BWP30P140LVT U2012 ( .I(ptr_next[28]), .ZN(n1913) );
  HA1D1BWP30P140LVT U2013 ( .A(ptr_next[28]), .B(n1911), .CO(n1914), .S(n1912)
         );
  MOAI22D1BWP30P140LVT U2014 ( .A1(n1913), .A2(n1835), .B1(n6), .B2(n1912), 
        .ZN(n1087) );
  INVD1BWP30P140LVT U2015 ( .I(ptr_next[29]), .ZN(n1916) );
  MOAI22D1BWP30P140LVT U2016 ( .A1(n1916), .A2(n1835), .B1(n6), .B2(n1915), 
        .ZN(n1086) );
  AOI21D1BWP30P140LVT U2017 ( .A1(n1984), .A2(delay_matrix_N_1_next[17]), .B(
        n1807), .ZN(n1917) );
  OAI211D1BWP30P140LVT U2018 ( .A1(n1933), .A2(n1919), .B(n1918), .C(n1917), 
        .ZN(n1002) );
  AOI21D1BWP30P140LVT U2019 ( .A1(n1984), .A2(delay_matrix_N_1_next[18]), .B(
        n1807), .ZN(n1920) );
  OAI211D1BWP30P140LVT U2020 ( .A1(n1933), .A2(n1922), .B(n1921), .C(n1920), 
        .ZN(n1001) );
  AOI21D1BWP30P140LVT U2021 ( .A1(n1984), .A2(delay_matrix_N_1_next[16]), .B(
        n1807), .ZN(n1923) );
  OAI211D1BWP30P140LVT U2022 ( .A1(n1933), .A2(n1925), .B(n1924), .C(n1923), 
        .ZN(n1003) );
  AOI21D1BWP30P140LVT U2023 ( .A1(n1984), .A2(delay_matrix_N_1_next[15]), .B(
        n1807), .ZN(n1926) );
  OAI211D1BWP30P140LVT U2024 ( .A1(n1933), .A2(n1928), .B(n1927), .C(n1926), 
        .ZN(n1004) );
  AOI21D1BWP30P140LVT U2025 ( .A1(n1984), .A2(delay_matrix_N_1_next[19]), .B(
        n1807), .ZN(n1930) );
  OAI211D1BWP30P140LVT U2026 ( .A1(n1933), .A2(n1932), .B(n1931), .C(n1930), 
        .ZN(n1000) );
  INVD1BWP30P140LVT U2027 ( .I(delay_matrix_N_1[34]), .ZN(n1936) );
  AOI21D1BWP30P140LVT U2028 ( .A1(n1984), .A2(delay_matrix_N_1_next[34]), .B(
        n1807), .ZN(n1934) );
  OAI211D1BWP30P140LVT U2029 ( .A1(n1957), .A2(n1936), .B(n1935), .C(n1934), 
        .ZN(n985) );
  INVD1BWP30P140LVT U2030 ( .I(delay_matrix_N_1[29]), .ZN(n1939) );
  AOI21D1BWP30P140LVT U2031 ( .A1(n1984), .A2(delay_matrix_N_1_next[29]), .B(
        n1807), .ZN(n1937) );
  OAI211D1BWP30P140LVT U2032 ( .A1(n1957), .A2(n1939), .B(n1938), .C(n1937), 
        .ZN(n990) );
  INVD1BWP30P140LVT U2033 ( .I(delay_matrix_N_1[31]), .ZN(n1942) );
  AOI21D1BWP30P140LVT U2034 ( .A1(n1984), .A2(delay_matrix_N_1_next[31]), .B(
        n1807), .ZN(n1940) );
  OAI211D1BWP30P140LVT U2035 ( .A1(n1957), .A2(n1942), .B(n1941), .C(n1940), 
        .ZN(n988) );
  INVD1BWP30P140LVT U2036 ( .I(delay_matrix_N_1[30]), .ZN(n1945) );
  AOI21D1BWP30P140LVT U2037 ( .A1(n1984), .A2(delay_matrix_N_1_next[30]), .B(
        n1807), .ZN(n1943) );
  OAI211D1BWP30P140LVT U2038 ( .A1(n1957), .A2(n1945), .B(n1944), .C(n1943), 
        .ZN(n989) );
  INVD1BWP30P140LVT U2039 ( .I(delay_matrix_N_1[33]), .ZN(n1948) );
  AOI21D1BWP30P140LVT U2040 ( .A1(n1984), .A2(delay_matrix_N_1_next[33]), .B(
        n1807), .ZN(n1946) );
  OAI211D1BWP30P140LVT U2041 ( .A1(n1957), .A2(n1948), .B(n1947), .C(n1946), 
        .ZN(n986) );
  INVD1BWP30P140LVT U2042 ( .I(delay_matrix_N_1[36]), .ZN(n1952) );
  AOI21D1BWP30P140LVT U2043 ( .A1(n1984), .A2(delay_matrix_N_1_next[36]), .B(
        n1807), .ZN(n1950) );
  OAI211D1BWP30P140LVT U2044 ( .A1(n1957), .A2(n1952), .B(n1951), .C(n1950), 
        .ZN(n983) );
  INVD1BWP30P140LVT U2045 ( .I(delay_matrix_N_1[32]), .ZN(n1956) );
  AOI21D1BWP30P140LVT U2046 ( .A1(n1984), .A2(delay_matrix_N_1_next[32]), .B(
        n1807), .ZN(n1954) );
  OAI211D1BWP30P140LVT U2047 ( .A1(n1957), .A2(n1956), .B(n1955), .C(n1954), 
        .ZN(n987) );
  AOI21D1BWP30P140LVT U2048 ( .A1(n1984), .A2(delay_matrix_N_1_next[47]), .B(
        n1807), .ZN(n1959) );
  OAI211D1BWP30P140LVT U2049 ( .A1(n1988), .A2(n1961), .B(n1960), .C(n1959), 
        .ZN(n972) );
  AOI21D1BWP30P140LVT U2050 ( .A1(n1984), .A2(delay_matrix_N_1_next[48]), .B(
        n1807), .ZN(n1963) );
  OAI211D1BWP30P140LVT U2051 ( .A1(n1988), .A2(n1965), .B(n1964), .C(n1963), 
        .ZN(n971) );
  AOI21D1BWP30P140LVT U2052 ( .A1(n1984), .A2(delay_matrix_N_1_next[45]), .B(
        n1807), .ZN(n1967) );
  OAI211D1BWP30P140LVT U2053 ( .A1(n1988), .A2(n1969), .B(n1968), .C(n1967), 
        .ZN(n974) );
  AOI21D1BWP30P140LVT U2054 ( .A1(n1984), .A2(delay_matrix_N_1_next[43]), .B(
        n1807), .ZN(n1971) );
  OAI211D1BWP30P140LVT U2055 ( .A1(n1988), .A2(n1973), .B(n1972), .C(n1971), 
        .ZN(n976) );
  AOI21D1BWP30P140LVT U2056 ( .A1(n1984), .A2(delay_matrix_N_1_next[46]), .B(
        n1807), .ZN(n1975) );
  OAI211D1BWP30P140LVT U2057 ( .A1(n1988), .A2(n1977), .B(n1976), .C(n1975), 
        .ZN(n973) );
  AOI21D1BWP30P140LVT U2058 ( .A1(n1984), .A2(delay_matrix_N_1_next[44]), .B(
        n1807), .ZN(n1979) );
  OAI211D1BWP30P140LVT U2059 ( .A1(n1988), .A2(n1981), .B(n1980), .C(n1979), 
        .ZN(n975) );
  AOI21D1BWP30P140LVT U2060 ( .A1(n1984), .A2(delay_matrix_N_1_next[49]), .B(
        n1807), .ZN(n1985) );
  OAI211D1BWP30P140LVT U2061 ( .A1(n1988), .A2(n1987), .B(n1986), .C(n1985), 
        .ZN(n970) );
  INVD1BWP30P140LVT U2062 ( .I(calc_glob_controller_prefetch_start_int[0]), 
        .ZN(n2059) );
  OR2D1BWP30P140LVT U2063 ( .A1(n1990), .A2(n1989), .Z(n1993) );
  OAI22D1BWP30P140LVT U2064 ( .A1(n2023), .A2(n2059), .B1(n2079), .B2(n2014), 
        .ZN(N4201) );
  INVD1BWP30P140LVT U2065 ( .I(calc_glob_controller_prefetch_start_int[1]), 
        .ZN(n2066) );
  OAI22D1BWP30P140LVT U2066 ( .A1(n2023), .A2(n2066), .B1(n2079), .B2(n2086), 
        .ZN(N4202) );
  INVD1BWP30P140LVT U2067 ( .I(calc_glob_controller_prefetch_start_int[7]), 
        .ZN(n2064) );
  OAI22D1BWP30P140LVT U2068 ( .A1(n2023), .A2(n2064), .B1(n2079), .B2(n2103), 
        .ZN(N4208) );
  INVD1BWP30P140LVT U2069 ( .I(calc_glob_controller_prefetch_start_int[2]), 
        .ZN(n2063) );
  OAI22D1BWP30P140LVT U2070 ( .A1(n2023), .A2(n2063), .B1(n2079), .B2(n12), 
        .ZN(N4203) );
  INVD1BWP30P140LVT U2071 ( .I(calc_glob_controller_prefetch_start_int[6]), 
        .ZN(n2065) );
  OAI22D1BWP30P140LVT U2072 ( .A1(n2023), .A2(n2065), .B1(n2079), .B2(n2121), 
        .ZN(N4207) );
  INVD2BWP30P140LVT U2073 ( .I(n1995), .ZN(n1997) );
  INVD1BWP30P140LVT U2074 ( .I(local_controller_id_int[5]), .ZN(n2060) );
  OAI22D1BWP30P140LVT U2075 ( .A1(n1997), .A2(n2060), .B1(n2079), .B2(n1996), 
        .ZN(N4214) );
  INVD1BWP30P140LVT U2076 ( .I(local_controller_id_int[1]), .ZN(n2056) );
  OAI22D1BWP30P140LVT U2077 ( .A1(n1997), .A2(n2056), .B1(n2079), .B2(n2115), 
        .ZN(N4210) );
  INVD1BWP30P140LVT U2078 ( .I(local_controller_id_int[4]), .ZN(n2061) );
  OAI22D1BWP30P140LVT U2079 ( .A1(n1997), .A2(n2061), .B1(n2079), .B2(n2009), 
        .ZN(N4213) );
  INVD1BWP30P140LVT U2080 ( .I(local_controller_id_int[3]), .ZN(n2062) );
  OAI22D1BWP30P140LVT U2081 ( .A1(n1997), .A2(n2062), .B1(n2079), .B2(n2006), 
        .ZN(N4212) );
  INVD1BWP30P140LVT U2082 ( .I(local_controller_id_int[0]), .ZN(n2057) );
  OAI22D1BWP30P140LVT U2083 ( .A1(n1997), .A2(n2057), .B1(n2079), .B2(n2021), 
        .ZN(N4209) );
  INVD1BWP30P140LVT U2084 ( .I(local_controller_id_int[2]), .ZN(n2058) );
  OAI22D1BWP30P140LVT U2085 ( .A1(n1997), .A2(n2058), .B1(n2079), .B2(n2118), 
        .ZN(N4211) );
  INR2D1BWP30P140LVT U2086 ( .A1(prefetch_bypass_start_addr[1]), .B1(n2172), 
        .ZN(n1998) );
  OAI21D1BWP30P140LVT U2087 ( .A1(n2124), .A2(n2086), .B(n1999), .ZN(n795) );
  MOAI22D1BWP30P140LVT U2088 ( .A1(n2003), .A2(n2002), .B1(table_ptr[1]), .B2(
        n2001), .ZN(n811) );
  INR2D1BWP30P140LVT U2089 ( .A1(prefetch_bypass_start_addr[11]), .B1(n2172), 
        .ZN(n2004) );
  OAI21D1BWP30P140LVT U2090 ( .A1(n2124), .A2(n2006), .B(n2005), .ZN(n785) );
  INR2D1BWP30P140LVT U2091 ( .A1(prefetch_bypass_start_addr[12]), .B1(n2172), 
        .ZN(n2007) );
  OAI21D1BWP30P140LVT U2092 ( .A1(n2124), .A2(n2009), .B(n2008), .ZN(n784) );
  INR2D1BWP30P140LVT U2093 ( .A1(prefetch_bypass_start_addr[3]), .B1(n2172), 
        .ZN(n2010) );
  OAI21D1BWP30P140LVT U2094 ( .A1(n2124), .A2(n2091), .B(n2011), .ZN(n793) );
  INR2D1BWP30P140LVT U2095 ( .A1(prefetch_bypass_start_addr[0]), .B1(n2172), 
        .ZN(n2012) );
  OAI21D1BWP30P140LVT U2096 ( .A1(n2124), .A2(n2014), .B(n2013), .ZN(n796) );
  INR2D1BWP30P140LVT U2097 ( .A1(prefetch_bypass_start_addr[5]), .B1(n2172), 
        .ZN(n2015) );
  OAI21D1BWP30P140LVT U2098 ( .A1(n2124), .A2(n2097), .B(n2016), .ZN(n791) );
  INR2D1BWP30P140LVT U2099 ( .A1(prefetch_bypass_start_addr[2]), .B1(n2172), 
        .ZN(n2017) );
  OAI21D1BWP30P140LVT U2100 ( .A1(n2124), .A2(n12), .B(n2018), .ZN(n794) );
  INR2D1BWP30P140LVT U2101 ( .A1(prefetch_bypass_start_addr[8]), .B1(n2172), 
        .ZN(n2019) );
  OAI21D1BWP30P140LVT U2102 ( .A1(n2124), .A2(n2021), .B(n2020), .ZN(n788) );
  NR2D1BWP30P140LVT U2103 ( .A1(n2087), .A2(n2086), .ZN(n2049) );
  NR2D1BWP30P140LVT U2104 ( .A1(n2156), .A2(n2014), .ZN(n2051) );
  ND2OPTIBD1BWP30P140LVT U2105 ( .A1(n2087), .A2(n2086), .ZN(n2050) );
  OAI21D1BWP30P140LVT U2106 ( .A1(n2049), .A2(n2051), .B(n2050), .ZN(n2028) );
  OR2D1BWP30P140LVT U2107 ( .A1(n2088), .A2(n12), .Z(n2027) );
  XNR2UD1BWP30P140LVT U2108 ( .A1(n2028), .A2(n2022), .ZN(n2024) );
  BUFFD4BWP30P140LVT U2109 ( .I(n2023), .Z(n2081) );
  INR2D1BWP30P140LVT U2110 ( .A1(n2024), .B1(n2081), .ZN(N4192) );
  XNR2UD1BWP30P140LVT U2111 ( .A1(n2156), .A2(n2155), .ZN(n2025) );
  INR2D1BWP30P140LVT U2112 ( .A1(n2025), .B1(n2081), .ZN(N4190) );
  AOI21D1BWP30P140LVT U2113 ( .A1(n2028), .A2(n2027), .B(n2089), .ZN(n2034) );
  NR2D1BWP30P140LVT U2114 ( .A1(n2092), .A2(n2091), .ZN(n2031) );
  ND2OPTIBD1BWP30P140LVT U2115 ( .A1(n2092), .A2(n2091), .ZN(n2032) );
  OR2D1BWP30P140LVT U2116 ( .A1(n2094), .A2(n2), .Z(n2037) );
  XNR2UD1BWP30P140LVT U2117 ( .A1(n2038), .A2(n2029), .ZN(n2030) );
  INR2D1BWP30P140LVT U2118 ( .A1(n2030), .B1(n2081), .ZN(N4194) );
  XOR2UD1BWP30P140LVT U2119 ( .A1(n2034), .A2(n2033), .Z(n2035) );
  INR2D1BWP30P140LVT U2120 ( .A1(n2035), .B1(n2081), .ZN(N4193) );
  NR2D1BWP30P140LVT U2121 ( .A1(n2098), .A2(n2097), .ZN(n2044) );
  OAI21D1BWP30P140LVT U2122 ( .A1(n2047), .A2(n2044), .B(n2045), .ZN(n2042) );
  OR2D1BWP30P140LVT U2123 ( .A1(n2100), .A2(n2121), .Z(n2040) );
  XNR2UD1BWP30P140LVT U2124 ( .A1(n2042), .A2(n2041), .ZN(n2043) );
  INR2D1BWP30P140LVT U2125 ( .A1(n2043), .B1(n2081), .ZN(N4196) );
  XOR2UD1BWP30P140LVT U2126 ( .A1(n2047), .A2(n2046), .Z(n2048) );
  INR2D1BWP30P140LVT U2127 ( .A1(n2048), .B1(n2081), .ZN(N4195) );
  XOR2UD1BWP30P140LVT U2128 ( .A1(n2052), .A2(n2051), .Z(n2053) );
  INR2D1BWP30P140LVT U2129 ( .A1(n2053), .B1(n2081), .ZN(N4191) );
  NR3D0P7BWP30P140LVT U2130 ( .A1(n2068), .A2(n2067), .A3(n2056), .ZN(N4232)
         );
  NR3D0P7BWP30P140LVT U2131 ( .A1(n2068), .A2(n2067), .A3(n2057), .ZN(N4231)
         );
  NR3D0P7BWP30P140LVT U2132 ( .A1(n2068), .A2(n2067), .A3(n2058), .ZN(N4233)
         );
  INVD1BWP30P140LVT U2133 ( .I(calc_glob_dest_addr_int[1]), .ZN(n2076) );
  NR3D0P7BWP30P140LVT U2134 ( .A1(n2068), .A2(n2067), .A3(n2076), .ZN(N4238)
         );
  NR3D0P7BWP30P140LVT U2135 ( .A1(n2068), .A2(n2067), .A3(n2059), .ZN(N4223)
         );
  NR3D0P7BWP30P140LVT U2136 ( .A1(n2068), .A2(n2067), .A3(n2060), .ZN(N4236)
         );
  NR3D0P7BWP30P140LVT U2137 ( .A1(n2068), .A2(n2067), .A3(n2061), .ZN(N4235)
         );
  NR3D0P7BWP30P140LVT U2138 ( .A1(n2068), .A2(n2067), .A3(n2062), .ZN(N4234)
         );
  INVD1BWP30P140LVT U2139 ( .I(calc_glob_dest_addr_int[2]), .ZN(n2073) );
  NR3D0P7BWP30P140LVT U2140 ( .A1(n2068), .A2(n2067), .A3(n2073), .ZN(N4239)
         );
  NR3D0P7BWP30P140LVT U2141 ( .A1(n2068), .A2(n2067), .A3(n2063), .ZN(N4225)
         );
  NR3D0P7BWP30P140LVT U2142 ( .A1(n2068), .A2(n2067), .A3(n2064), .ZN(N4230)
         );
  NR3D0P7BWP30P140LVT U2143 ( .A1(n2068), .A2(n2067), .A3(n2065), .ZN(N4229)
         );
  INVD1BWP30P140LVT U2144 ( .I(calc_glob_dest_addr_int[3]), .ZN(n2070) );
  NR3D0P7BWP30P140LVT U2145 ( .A1(n2068), .A2(n2067), .A3(n2070), .ZN(N4240)
         );
  INVD1BWP30P140LVT U2146 ( .I(calc_glob_controller_prefetch_start_int[4]), 
        .ZN(n2080) );
  NR3D0P7BWP30P140LVT U2147 ( .A1(n2068), .A2(n2067), .A3(n2080), .ZN(N4227)
         );
  INVD1BWP30P140LVT U2148 ( .I(calc_glob_controller_prefetch_start_int[3]), 
        .ZN(n2078) );
  NR3D0P7BWP30P140LVT U2149 ( .A1(n2068), .A2(n2067), .A3(n2078), .ZN(N4226)
         );
  NR3D0P7BWP30P140LVT U2150 ( .A1(n2068), .A2(n2067), .A3(n2066), .ZN(N4224)
         );
  INVD1BWP30P140LVT U2151 ( .I(calc_glob_controller_prefetch_start_int[5]), 
        .ZN(n2077) );
  NR3D0P7BWP30P140LVT U2152 ( .A1(n2068), .A2(n2067), .A3(n2077), .ZN(N4228)
         );
  INVD1BWP30P140LVT U2153 ( .I(n2225), .ZN(n2071) );
  OAI22D1BWP30P140LVT U2154 ( .A1(n2081), .A2(n2070), .B1(n2069), .B2(n2071), 
        .ZN(N4200) );
  OAI22D1BWP30P140LVT U2155 ( .A1(n2081), .A2(n2073), .B1(n2072), .B2(n2071), 
        .ZN(N4199) );
  INVD1BWP30P140LVT U2156 ( .I(n2226), .ZN(n2074) );
  OAI22D1BWP30P140LVT U2157 ( .A1(n2081), .A2(n2076), .B1(n2075), .B2(n2074), 
        .ZN(N4198) );
  OAI22D1BWP30P140LVT U2158 ( .A1(n2081), .A2(n2077), .B1(n2079), .B2(n2097), 
        .ZN(N4206) );
  OAI22D1BWP30P140LVT U2159 ( .A1(n2081), .A2(n2078), .B1(n2079), .B2(n2091), 
        .ZN(N4204) );
  OAI22D1BWP30P140LVT U2160 ( .A1(n2081), .A2(n2080), .B1(n2079), .B2(n2), 
        .ZN(N4205) );
  INR2D1BWP30P140LVT U2161 ( .A1(prefetch_bypass_start_addr[4]), .B1(n2172), 
        .ZN(n2082) );
  OAI21D1BWP30P140LVT U2162 ( .A1(n2124), .A2(n2), .B(n2083), .ZN(n792) );
  NR2D1BWP30P140LVT U2163 ( .A1(n2087), .A2(n2086), .ZN(n2147) );
  NR2D1BWP30P140LVT U2164 ( .A1(n2156), .A2(n2155), .ZN(n2150) );
  ND2OPTIBD1BWP30P140LVT U2165 ( .A1(n2087), .A2(n2086), .ZN(n2148) );
  OR2D1BWP30P140LVT U2166 ( .A1(n2088), .A2(n12), .Z(n2141) );
  ND2OPTIBD1BWP30P140LVT U2167 ( .A1(n2088), .A2(n12), .ZN(n2140) );
  INVD1BWP30P140LVT U2168 ( .I(n2140), .ZN(n2089) );
  INVD1BWP30P140LVT U2169 ( .I(n2090), .ZN(n2091) );
  NR2D1BWP30P140LVT U2170 ( .A1(n2092), .A2(n2091), .ZN(n2132) );
  ND2OPTIBD1BWP30P140LVT U2171 ( .A1(n2092), .A2(n2091), .ZN(n2133) );
  OR2D1BWP30P140LVT U2172 ( .A1(n2094), .A2(n2), .Z(n2161) );
  INVD1BWP30P140LVT U2173 ( .I(n2160), .ZN(n2095) );
  AOI21D2BWP30P140LVT U2174 ( .A1(n2163), .A2(n2161), .B(n2095), .ZN(n2171) );
  INVD1BWP30P140LVT U2175 ( .I(n2096), .ZN(n2097) );
  NR2D1BWP30P140LVT U2176 ( .A1(n2098), .A2(n2097), .ZN(n2167) );
  OR2D1BWP30P140LVT U2177 ( .A1(n2100), .A2(n2121), .Z(n2126) );
  INVD1BWP30P140LVT U2178 ( .I(n2125), .ZN(n2101) );
  INVD1BWP30P140LVT U2179 ( .I(n2102), .ZN(n2103) );
  OR2D1BWP30P140LVT U2180 ( .A1(n2104), .A2(n2103), .Z(n2106) );
  ND2D1BWP30P140LVT U2181 ( .A1(n2106), .A2(n2105), .ZN(n2107) );
  XOR2UD1BWP30P140LVT U2182 ( .A1(n2108), .A2(n2107), .Z(n2109) );
  INR2D1BWP30P140LVT U2183 ( .A1(prefetch_bypass_cycles[7]), .B1(n2172), .ZN(
        n2110) );
  INR2D1BWP30P140LVT U2184 ( .A1(prefetch_bypass_start_addr[9]), .B1(n2172), 
        .ZN(n2113) );
  OAI21D1BWP30P140LVT U2185 ( .A1(n2124), .A2(n2115), .B(n2114), .ZN(n787) );
  INR2D1BWP30P140LVT U2186 ( .A1(prefetch_bypass_start_addr[10]), .B1(n2172), 
        .ZN(n2116) );
  OAI21D1BWP30P140LVT U2187 ( .A1(n2124), .A2(n2118), .B(n2117), .ZN(n786) );
  INR2D1BWP30P140LVT U2188 ( .A1(prefetch_bypass_start_addr[6]), .B1(n2172), 
        .ZN(n2119) );
  ND2OPTIBD1BWP30P140LVT U2189 ( .A1(n2174), .A2(n2119), .ZN(n2120) );
  OAI21D1BWP30P140LVT U2190 ( .A1(n2124), .A2(n2121), .B(n2120), .ZN(n790) );
  INR2D1BWP30P140LVT U2191 ( .A1(prefetch_bypass_start_addr[7]), .B1(n2172), 
        .ZN(n2122) );
  OAI21D1BWP30P140LVT U2192 ( .A1(n2124), .A2(n2103), .B(n2123), .ZN(n789) );
  ND2D1BWP30P140LVT U2193 ( .A1(n2126), .A2(n2125), .ZN(n2127) );
  XNR2UD1BWP30P140LVT U2194 ( .A1(n2128), .A2(n2127), .ZN(n2131) );
  INR2D1BWP30P140LVT U2195 ( .A1(prefetch_bypass_cycles[6]), .B1(n2172), .ZN(
        n2129) );
  IOA21D1BWP30P140LVT U2196 ( .A1(n2131), .A2(n2176), .B(n2130), .ZN(n798) );
  INVD1BWP30P140LVT U2197 ( .I(n2132), .ZN(n2134) );
  ND2D1BWP30P140LVT U2198 ( .A1(n2134), .A2(n2133), .ZN(n2135) );
  XOR2UD1BWP30P140LVT U2199 ( .A1(n2136), .A2(n2135), .Z(n2139) );
  INR2D1BWP30P140LVT U2200 ( .A1(prefetch_bypass_cycles[3]), .B1(n2172), .ZN(
        n2137) );
  IOA21D1BWP30P140LVT U2201 ( .A1(n2176), .A2(n2139), .B(n2138), .ZN(n801) );
  ND2D1BWP30P140LVT U2202 ( .A1(n2141), .A2(n2140), .ZN(n2142) );
  XNR2UD1BWP30P140LVT U2203 ( .A1(n2143), .A2(n2142), .ZN(n2146) );
  INR2D1BWP30P140LVT U2204 ( .A1(prefetch_bypass_cycles[2]), .B1(n2172), .ZN(
        n2144) );
  IOA21D1BWP30P140LVT U2205 ( .A1(n2176), .A2(n2146), .B(n2145), .ZN(n802) );
  INVD1BWP30P140LVT U2206 ( .I(n2147), .ZN(n2149) );
  ND2D1BWP30P140LVT U2207 ( .A1(n2149), .A2(n2148), .ZN(n2151) );
  XOR2UD1BWP30P140LVT U2208 ( .A1(n2151), .A2(n2150), .Z(n2154) );
  INR2D1BWP30P140LVT U2209 ( .A1(prefetch_bypass_cycles[1]), .B1(n2172), .ZN(
        n2152) );
  IOA21D1BWP30P140LVT U2210 ( .A1(n2176), .A2(n2154), .B(n2153), .ZN(n803) );
  XNR2UD1BWP30P140LVT U2211 ( .A1(n2156), .A2(n2155), .ZN(n2159) );
  INR2D1BWP30P140LVT U2212 ( .A1(prefetch_bypass_cycles[0]), .B1(n2172), .ZN(
        n2157) );
  IOA21D1BWP30P140LVT U2213 ( .A1(n2176), .A2(n2159), .B(n2158), .ZN(n804) );
  ND2D1BWP30P140LVT U2214 ( .A1(n2161), .A2(n2160), .ZN(n2162) );
  XNR2UD1BWP30P140LVT U2215 ( .A1(n2163), .A2(n2162), .ZN(n2166) );
  INR2D1BWP30P140LVT U2216 ( .A1(prefetch_bypass_cycles[4]), .B1(n2172), .ZN(
        n2164) );
  IOA21D1BWP30P140LVT U2217 ( .A1(n2166), .A2(n2176), .B(n2165), .ZN(n800) );
  INVD1BWP30P140LVT U2218 ( .I(n2167), .ZN(n2169) );
  ND2D1BWP30P140LVT U2219 ( .A1(n2169), .A2(n2168), .ZN(n2170) );
  XOR2UD1BWP30P140LVT U2220 ( .A1(n2171), .A2(n2170), .Z(n2177) );
  INR2D1BWP30P140LVT U2221 ( .A1(prefetch_bypass_cycles[5]), .B1(n2172), .ZN(
        n2173) );
  IOA21D1BWP30P140LVT U2222 ( .A1(n2177), .A2(n2176), .B(n2175), .ZN(n799) );
  AOI22D1BWP30P140LVT U2223 ( .A1(obj_id[0]), .A2(n2179), .B1(n1802), .B2(
        obj_id_next[0]), .ZN(n2178) );
  OAI21D1BWP30P140LVT U2224 ( .A1(n2187), .A2(n2181), .B(n2178), .ZN(n963) );
  AOI22D1BWP30P140LVT U2225 ( .A1(obj_id[1]), .A2(n2179), .B1(n1773), .B2(
        obj_id_next[1]), .ZN(n2180) );
  OAI21D1BWP30P140LVT U2226 ( .A1(n2190), .A2(n2181), .B(n2180), .ZN(n962) );
  AOI22D1BWP30P140LVT U2227 ( .A1(obj_id[2]), .A2(n2183), .B1(n1773), .B2(
        obj_id_next[2]), .ZN(n2182) );
  OAI21D1BWP30P140LVT U2228 ( .A1(n2187), .A2(n2185), .B(n2182), .ZN(n961) );
  AOI22D1BWP30P140LVT U2229 ( .A1(obj_id[3]), .A2(n2183), .B1(n1802), .B2(
        obj_id_next[3]), .ZN(n2184) );
  OAI21D1BWP30P140LVT U2230 ( .A1(n2190), .A2(n2185), .B(n2184), .ZN(n960) );
  AOI22D1BWP30P140LVT U2231 ( .A1(obj_id[4]), .A2(n2188), .B1(n1773), .B2(
        obj_id_next[4]), .ZN(n2186) );
  OAI21D1BWP30P140LVT U2232 ( .A1(n2191), .A2(n2187), .B(n2186), .ZN(n959) );
  AOI22D1BWP30P140LVT U2233 ( .A1(obj_id[5]), .A2(n2188), .B1(n1802), .B2(
        obj_id_next[5]), .ZN(n2189) );
  OAI21D1BWP30P140LVT U2234 ( .A1(n2191), .A2(n2190), .B(n2189), .ZN(n958) );
  AOI22D1BWP30P140LVT U2235 ( .A1(delay_matrix_N_1_original[10]), .A2(n2194), 
        .B1(scenario_update), .B2(delay_matrix_N_1_next_original[10]), .ZN(
        n2192) );
  OAI211D1BWP30P140LVT U2236 ( .A1(n2206), .A2(n2196), .B(n2192), .C(n1821), 
        .ZN(n857) );
  AOI22D1BWP30P140LVT U2237 ( .A1(delay_matrix_N_1_original[12]), .A2(n2194), 
        .B1(n561), .B2(delay_matrix_N_1_next_original[12]), .ZN(n2193) );
  OAI21D1BWP30P140LVT U2238 ( .A1(n2199), .A2(n2196), .B(n2193), .ZN(n855) );
  AOI22D1BWP30P140LVT U2239 ( .A1(delay_matrix_N_1_original[13]), .A2(n2194), 
        .B1(n561), .B2(delay_matrix_N_1_next_original[13]), .ZN(n2195) );
  OAI21D1BWP30P140LVT U2240 ( .A1(n2203), .A2(n2196), .B(n2195), .ZN(n854) );
  AOI22D1BWP30P140LVT U2241 ( .A1(delay_matrix_N_1_original[24]), .A2(n2200), 
        .B1(n561), .B2(delay_matrix_N_1_next_original[24]), .ZN(n2197) );
  OAI211D1BWP30P140LVT U2242 ( .A1(n2206), .A2(n2202), .B(n2197), .C(n1821), 
        .ZN(n843) );
  AOI22D1BWP30P140LVT U2243 ( .A1(delay_matrix_N_1_original[26]), .A2(n2200), 
        .B1(n1802), .B2(delay_matrix_N_1_next_original[26]), .ZN(n2198) );
  OAI21D1BWP30P140LVT U2244 ( .A1(n2199), .A2(n2202), .B(n2198), .ZN(n841) );
  AOI22D1BWP30P140LVT U2245 ( .A1(delay_matrix_N_1_original[27]), .A2(n2200), 
        .B1(n561), .B2(delay_matrix_N_1_next_original[27]), .ZN(n2201) );
  OAI21D1BWP30P140LVT U2246 ( .A1(n2203), .A2(n2202), .B(n2201), .ZN(n840) );
  AOI22D1BWP30P140LVT U2247 ( .A1(n2204), .A2(delay_matrix_N_1_original[38]), 
        .B1(n1773), .B2(delay_matrix_N_1_next_original[38]), .ZN(n2205) );
  OAI211D1BWP30P140LVT U2248 ( .A1(n2207), .A2(n2206), .B(n2205), .C(n1821), 
        .ZN(n829) );
endmodule


module addrGen ( CLK, rst, start, addr, counter_up );
  output [5:0] addr;
  output [7:0] counter_up;
  input CLK, rst, start;
  wire   n37, n38, N28, N29, N30, N31, N32, N33, N34, N35, n12, n13, n14, n15,
         n16, n17, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34;

  DFQD1BWP30P140LVT counter_up_reg_0_ ( .D(N28), .CP(CLK), .Q(counter_up[0])
         );
  DFQD1BWP30P140LVT counter_up_reg_1_ ( .D(N29), .CP(CLK), .Q(counter_up[1])
         );
  DFQD1BWP30P140LVT counter_up_reg_2_ ( .D(N30), .CP(CLK), .Q(counter_up[2])
         );
  DFQD1BWP30P140LVT counter_up_reg_3_ ( .D(N31), .CP(CLK), .Q(counter_up[3])
         );
  DFQD1BWP30P140LVT counter_up_reg_4_ ( .D(N32), .CP(CLK), .Q(counter_up[4])
         );
  DFQD1BWP30P140LVT counter_up_reg_5_ ( .D(N33), .CP(CLK), .Q(counter_up[5])
         );
  DFQD1BWP30P140LVT counter_up_reg_6_ ( .D(N34), .CP(CLK), .Q(counter_up[6])
         );
  DFQD1BWP30P140LVT counter_up_reg_7_ ( .D(N35), .CP(CLK), .Q(counter_up[7])
         );
  DFQD1BWP30P140LVT addr_reg_4_ ( .D(n16), .CP(CLK), .Q(addr[4]) );
  DFQD1BWP30P140LVT addr_reg_0_ ( .D(n12), .CP(CLK), .Q(addr[0]) );
  DFQD1BWP30P140LVT addr_reg_2_ ( .D(n14), .CP(CLK), .Q(n38) );
  DFQD1BWP30P140LVT addr_reg_3_ ( .D(n15), .CP(CLK), .Q(n37) );
  DFQD4BWP30P140LVT addr_reg_5_ ( .D(n17), .CP(CLK), .Q(addr[5]) );
  DFQD4BWP30P140LVT addr_reg_1_ ( .D(n13), .CP(CLK), .Q(addr[1]) );
  INVD8BWP30P140LVT U3 ( .I(n26), .ZN(addr[3]) );
  INVD2BWP30P140LVT U4 ( .I(n37), .ZN(n26) );
  ND2D1BWP30P140LVT U5 ( .A1(n20), .A2(counter_up[7]), .ZN(n2) );
  ND2D1BWP30P140LVT U6 ( .A1(n29), .A2(n33), .ZN(n31) );
  INVD1BWP30P140LVT U7 ( .I(addr[1]), .ZN(n33) );
  AN4D0BWP30P140LVT U8 ( .A1(addr[5]), .A2(addr[3]), .A3(addr[2]), .A4(addr[1]), .Z(n3) );
  ND2D1BWP30P140LVT U9 ( .A1(n29), .A2(n26), .ZN(n25) );
  INVD1BWP30P140LVT U10 ( .I(counter_up[6]), .ZN(n11) );
  NR2D1BWP30P140LVT U11 ( .A1(n18), .A2(n11), .ZN(n20) );
  ND2D1BWP30P140LVT U12 ( .A1(n9), .A2(counter_up[5]), .ZN(n18) );
  INVD1BWP30P140LVT U13 ( .I(counter_up[4]), .ZN(n7) );
  NR2D1BWP30P140LVT U14 ( .A1(n8), .A2(n7), .ZN(n9) );
  ND2D1BWP30P140LVT U15 ( .A1(n6), .A2(counter_up[3]), .ZN(n8) );
  NR2D1BWP30P140LVT U16 ( .A1(n5), .A2(n4), .ZN(n6) );
  ND2D1BWP30P140LVT U17 ( .A1(counter_up[1]), .A2(counter_up[0]), .ZN(n5) );
  INVD1BWP30P140LVT U18 ( .I(n19), .ZN(n28) );
  IND2D1BWP30P140LVT U19 ( .A1(n10), .B1(n2), .ZN(n19) );
  INVD1BWP30P140LVT U20 ( .I(addr[4]), .ZN(n22) );
  INVD1BWP30P140LVT U21 ( .I(addr[0]), .ZN(n32) );
  INVD4BWP30P140LVT U22 ( .I(n1), .ZN(addr[2]) );
  INVD1BWP30P140LVT U23 ( .I(n38), .ZN(n1) );
  IND2D1BWP30P140LVT U24 ( .A1(rst), .B1(start), .ZN(n10) );
  INVD1BWP30P140LVT U25 ( .I(counter_up[2]), .ZN(n4) );
  NR2D1BWP30P140LVT U26 ( .A1(counter_up[0]), .A2(n19), .ZN(N28) );
  AOI211D1BWP30P140LVT U27 ( .A1(addr[4]), .A2(n3), .B(n2), .C(n10), .ZN(n29)
         );
  MAOI22D1BWP30P140LVT U28 ( .A1(addr[0]), .A2(n19), .B1(n29), .B2(addr[0]), 
        .ZN(n12) );
  OA211D1BWP30P140LVT U29 ( .A1(counter_up[1]), .A2(counter_up[0]), .B(n28), 
        .C(n5), .Z(N29) );
  AOI211D1BWP30P140LVT U30 ( .A1(n5), .A2(n4), .B(n6), .C(n19), .ZN(N30) );
  OA211D1BWP30P140LVT U31 ( .A1(n6), .A2(counter_up[3]), .B(n28), .C(n8), .Z(
        N31) );
  AOI211D1BWP30P140LVT U32 ( .A1(n8), .A2(n7), .B(n9), .C(n19), .ZN(N32) );
  OA211D1BWP30P140LVT U33 ( .A1(n9), .A2(counter_up[5]), .B(n28), .C(n18), .Z(
        N33) );
  AOI211D1BWP30P140LVT U34 ( .A1(n18), .A2(n11), .B(n20), .C(n10), .ZN(N34) );
  IAO21D1BWP30P140LVT U35 ( .A1(n20), .A2(counter_up[7]), .B(n19), .ZN(N35) );
  ND3D1BWP30P140LVT U36 ( .A1(addr[2]), .A2(addr[1]), .A3(addr[0]), .ZN(n24)
         );
  IND3D1BWP30P140LVT U37 ( .A1(n24), .B1(addr[3]), .B2(n29), .ZN(n23) );
  OAI21D1BWP30P140LVT U38 ( .A1(n29), .A2(n28), .B(addr[5]), .ZN(n21) );
  OAI21D1BWP30P140LVT U39 ( .A1(n23), .A2(n22), .B(n21), .ZN(n17) );
  AOI21D1BWP30P140LVT U40 ( .A1(n29), .A2(n24), .B(n28), .ZN(n27) );
  AOI32D1BWP30P140LVT U41 ( .A1(n27), .A2(addr[4]), .A3(n25), .B1(n23), .B2(
        n22), .ZN(n16) );
  OAI22D1BWP30P140LVT U42 ( .A1(n27), .A2(n26), .B1(n25), .B2(n24), .ZN(n15)
         );
  AOI21D1BWP30P140LVT U43 ( .A1(n29), .A2(n32), .B(n28), .ZN(n34) );
  ND3D1BWP30P140LVT U44 ( .A1(addr[1]), .A2(n29), .A3(addr[0]), .ZN(n30) );
  AOI32D1BWP30P140LVT U45 ( .A1(n34), .A2(addr[2]), .A3(n31), .B1(n30), .B2(n1), .ZN(n14) );
  OAI22D1BWP30P140LVT U46 ( .A1(n34), .A2(n33), .B1(n32), .B2(n31), .ZN(n13)
         );
endmodule


module prefetch_bypass_module ( CLK, reset, start, 
        prefetch_bypass_dest_addr_int, prefetch_bypass_cycles, 
        prefetch_bypass_start_addr, local_controller_id, sample_address, 
        data_in, prefetch_bypass_path_input_data, 
        prefetch_bypass_path_input_addr, prefetch_bypass_valid );
  input [3:0] prefetch_bypass_dest_addr_int;
  input [7:0] prefetch_bypass_cycles;
  input [13:0] prefetch_bypass_start_addr;
  input [5:0] local_controller_id;
  input [7:0] sample_address;
  input [31:0] data_in;
  output [31:0] prefetch_bypass_path_input_data;
  output [3:0] prefetch_bypass_path_input_addr;
  input CLK, reset, start;
  output prefetch_bypass_valid;
  wire   n62, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N79, N80, N82,
         N85, N88, N91, N94, N97, N100, N103, N106, N109, N112, N115, N118,
         N121, N124, N127, N130, N133, N136, N139, N142, N145, N148, N151,
         N154, N157, N160, N163, N166, N169, N172, N175, N178, N181, N184, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n61;
  wire   [7:0] prefetch_bypass_counter;
  tri   [31:0] prefetch_bypass_path_input_data;
  tri   [3:0] prefetch_bypass_path_input_addr;

  DFQD1BWP30P140LVT prefetch_bypass_path_input_addr_reg_3_ ( .D(
        prefetch_bypass_dest_addr_int[3]), .CP(CLK), .Q(N79) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_addr_reg_2_ ( .D(
        prefetch_bypass_dest_addr_int[2]), .CP(CLK), .Q(N82) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_addr_reg_1_ ( .D(
        prefetch_bypass_dest_addr_int[1]), .CP(CLK), .Q(N85) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_addr_reg_0_ ( .D(
        prefetch_bypass_dest_addr_int[0]), .CP(CLK), .Q(N88) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_31_ ( .D(data_in[31]), 
        .CP(CLK), .Q(N91) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_30_ ( .D(data_in[30]), 
        .CP(CLK), .Q(N94) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_29_ ( .D(data_in[29]), 
        .CP(CLK), .Q(N97) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_28_ ( .D(data_in[28]), 
        .CP(CLK), .Q(N100) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_27_ ( .D(data_in[27]), 
        .CP(CLK), .Q(N103) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_26_ ( .D(data_in[26]), 
        .CP(CLK), .Q(N106) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_25_ ( .D(data_in[25]), 
        .CP(CLK), .Q(N109) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_24_ ( .D(data_in[24]), 
        .CP(CLK), .Q(N112) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_23_ ( .D(data_in[23]), 
        .CP(CLK), .Q(N115) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_22_ ( .D(data_in[22]), 
        .CP(CLK), .Q(N118) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_21_ ( .D(data_in[21]), 
        .CP(CLK), .Q(N121) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_20_ ( .D(data_in[20]), 
        .CP(CLK), .Q(N124) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_19_ ( .D(data_in[19]), 
        .CP(CLK), .Q(N127) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_18_ ( .D(data_in[18]), 
        .CP(CLK), .Q(N130) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_17_ ( .D(data_in[17]), 
        .CP(CLK), .Q(N133) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_16_ ( .D(data_in[16]), 
        .CP(CLK), .Q(N136) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_15_ ( .D(data_in[15]), 
        .CP(CLK), .Q(N139) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_14_ ( .D(data_in[14]), 
        .CP(CLK), .Q(N142) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_13_ ( .D(data_in[13]), 
        .CP(CLK), .Q(N145) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_12_ ( .D(data_in[12]), 
        .CP(CLK), .Q(N148) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_11_ ( .D(data_in[11]), 
        .CP(CLK), .Q(N151) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_10_ ( .D(data_in[10]), 
        .CP(CLK), .Q(N154) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_9_ ( .D(data_in[9]), 
        .CP(CLK), .Q(N157) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_8_ ( .D(data_in[8]), 
        .CP(CLK), .Q(N160) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_7_ ( .D(data_in[7]), 
        .CP(CLK), .Q(N163) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_6_ ( .D(data_in[6]), 
        .CP(CLK), .Q(N166) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_5_ ( .D(data_in[5]), 
        .CP(CLK), .Q(N169) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_4_ ( .D(data_in[4]), 
        .CP(CLK), .Q(N172) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_3_ ( .D(data_in[3]), 
        .CP(CLK), .Q(N175) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_2_ ( .D(data_in[2]), 
        .CP(CLK), .Q(N178) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_1_ ( .D(data_in[1]), 
        .CP(CLK), .Q(N181) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_data_reg_0_ ( .D(data_in[0]), 
        .CP(CLK), .Q(N184) );
  DFQD1BWP30P140LVT prefetch_bypass_counter_reg_0_ ( .D(N65), .CP(CLK), .Q(
        prefetch_bypass_counter[0]) );
  DFQD1BWP30P140LVT prefetch_bypass_counter_reg_1_ ( .D(N66), .CP(CLK), .Q(
        prefetch_bypass_counter[1]) );
  DFQD1BWP30P140LVT prefetch_bypass_counter_reg_2_ ( .D(N67), .CP(CLK), .Q(
        prefetch_bypass_counter[2]) );
  DFQD1BWP30P140LVT prefetch_bypass_counter_reg_3_ ( .D(N68), .CP(CLK), .Q(
        prefetch_bypass_counter[3]) );
  DFQD1BWP30P140LVT prefetch_bypass_counter_reg_4_ ( .D(N69), .CP(CLK), .Q(
        prefetch_bypass_counter[4]) );
  DFQD1BWP30P140LVT prefetch_bypass_counter_reg_5_ ( .D(N70), .CP(CLK), .Q(
        prefetch_bypass_counter[5]) );
  DFQD1BWP30P140LVT prefetch_bypass_counter_reg_6_ ( .D(N71), .CP(CLK), .Q(
        prefetch_bypass_counter[6]) );
  DFQD1BWP30P140LVT prefetch_bypass_counter_reg_7_ ( .D(N72), .CP(CLK), .Q(
        prefetch_bypass_counter[7]) );
  DFQD1BWP30P140LVT prefetch_bypass_path_input_addr_tri_enable_reg_3_ ( .D(N64), .CP(CLK), .Q(N80) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_0_ ( .I(N184), .OE(
        n61), .Z(prefetch_bypass_path_input_data[0]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_1_ ( .I(N181), .OE(
        n61), .Z(prefetch_bypass_path_input_data[1]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_2_ ( .I(N178), .OE(
        n61), .Z(prefetch_bypass_path_input_data[2]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_3_ ( .I(N175), .OE(
        n61), .Z(prefetch_bypass_path_input_data[3]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_4_ ( .I(N172), .OE(
        n61), .Z(prefetch_bypass_path_input_data[4]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_5_ ( .I(N169), .OE(
        n61), .Z(prefetch_bypass_path_input_data[5]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_6_ ( .I(N166), .OE(
        n61), .Z(prefetch_bypass_path_input_data[6]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_7_ ( .I(N163), .OE(
        n61), .Z(prefetch_bypass_path_input_data[7]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_8_ ( .I(N160), .OE(
        n61), .Z(prefetch_bypass_path_input_data[8]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_9_ ( .I(N157), .OE(
        n61), .Z(prefetch_bypass_path_input_data[9]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_10_ ( .I(N154), .OE(
        n61), .Z(prefetch_bypass_path_input_data[10]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_11_ ( .I(N151), .OE(
        n61), .Z(prefetch_bypass_path_input_data[11]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_12_ ( .I(N148), .OE(
        n61), .Z(prefetch_bypass_path_input_data[12]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_13_ ( .I(N145), .OE(
        n61), .Z(prefetch_bypass_path_input_data[13]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_14_ ( .I(N142), .OE(
        n61), .Z(prefetch_bypass_path_input_data[14]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_15_ ( .I(N139), .OE(
        n61), .Z(prefetch_bypass_path_input_data[15]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_16_ ( .I(N136), .OE(
        n61), .Z(prefetch_bypass_path_input_data[16]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_17_ ( .I(N133), .OE(
        n61), .Z(prefetch_bypass_path_input_data[17]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_18_ ( .I(N130), .OE(
        n61), .Z(prefetch_bypass_path_input_data[18]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_19_ ( .I(N127), .OE(
        n61), .Z(prefetch_bypass_path_input_data[19]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_20_ ( .I(N124), .OE(
        n61), .Z(prefetch_bypass_path_input_data[20]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_21_ ( .I(N121), .OE(
        n61), .Z(prefetch_bypass_path_input_data[21]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_22_ ( .I(N118), .OE(
        n61), .Z(prefetch_bypass_path_input_data[22]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_23_ ( .I(N115), .OE(
        n61), .Z(prefetch_bypass_path_input_data[23]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_24_ ( .I(N112), .OE(
        n61), .Z(prefetch_bypass_path_input_data[24]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_25_ ( .I(N109), .OE(
        n61), .Z(prefetch_bypass_path_input_data[25]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_26_ ( .I(N106), .OE(
        n61), .Z(prefetch_bypass_path_input_data[26]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_27_ ( .I(N103), .OE(
        n61), .Z(prefetch_bypass_path_input_data[27]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_28_ ( .I(N100), .OE(
        n61), .Z(prefetch_bypass_path_input_data[28]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_29_ ( .I(N97), .OE(
        n61), .Z(prefetch_bypass_path_input_data[29]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_30_ ( .I(N94), .OE(
        n61), .Z(prefetch_bypass_path_input_data[30]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_data_tri_31_ ( .I(N91), .OE(
        n61), .Z(prefetch_bypass_path_input_data[31]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_addr_tri_0_ ( .I(N88), .OE(n61), .Z(prefetch_bypass_path_input_addr[0]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_addr_tri_1_ ( .I(N85), .OE(n61), .Z(prefetch_bypass_path_input_addr[1]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_addr_tri_2_ ( .I(N82), .OE(n61), .Z(prefetch_bypass_path_input_addr[2]) );
  BUFTD4BWP30P140LVT prefetch_bypass_path_input_addr_tri_3_ ( .I(N79), .OE(n61), .Z(prefetch_bypass_path_input_addr[3]) );
  DFQD1BWP30P140LVT prefetch_bypass_valid_reg ( .D(N73), .CP(CLK), .Q(n62) );
  INVD2BWP30P140LVT U3 ( .I(N80), .ZN(n61) );
  XOR2UD1BWP30P140LVT U4 ( .A1(prefetch_bypass_start_addr[9]), .A2(
        local_controller_id[1]), .Z(n44) );
  NR3D0P7BWP30P140LVT U5 ( .A1(n33), .A2(n32), .A3(n31), .ZN(n38) );
  AOI221D1BWP30P140LVT U6 ( .A1(n36), .A2(prefetch_bypass_start_addr[1]), .B1(
        prefetch_bypass_start_addr[8]), .B2(n35), .C(n34), .ZN(n37) );
  IND4D1BWP30P140LVT U7 ( .A1(n40), .B1(n39), .B2(n38), .B3(n37), .ZN(n41) );
  ND3OPTPAD1BWP30P140LVT U8 ( .A1(n20), .A2(n19), .A3(n18), .ZN(n42) );
  OAI22D2BWP30P140LVT U9 ( .A1(n36), .A2(prefetch_bypass_start_addr[1]), .B1(
        n35), .B2(prefetch_bypass_start_addr[8]), .ZN(n34) );
  XOR2UD1BWP30P140LVT U10 ( .A1(local_controller_id[2]), .A2(
        prefetch_bypass_start_addr[10]), .Z(n43) );
  INVD4BWP30P140LVT U11 ( .I(N73), .ZN(N64) );
  INVD1BWP30P140LVT U12 ( .I(local_controller_id[0]), .ZN(n35) );
  XNR2UD1BWP30P140LVT U13 ( .A1(prefetch_bypass_start_addr[4]), .A2(
        sample_address[4]), .ZN(n18) );
  NR2D1BWP30P140LVT U14 ( .A1(n56), .A2(n55), .ZN(n59) );
  ND2D1BWP30P140LVT U15 ( .A1(prefetch_bypass_counter[5]), .A2(n54), .ZN(n55)
         );
  INVD1BWP30P140LVT U16 ( .I(prefetch_bypass_counter[4]), .ZN(n53) );
  NR2D1BWP30P140LVT U17 ( .A1(n53), .A2(n52), .ZN(n54) );
  ND2D1BWP30P140LVT U18 ( .A1(prefetch_bypass_counter[3]), .A2(n51), .ZN(n52)
         );
  NR2D1BWP30P140LVT U19 ( .A1(n50), .A2(n49), .ZN(n51) );
  ND2D1BWP30P140LVT U20 ( .A1(prefetch_bypass_counter[1]), .A2(
        prefetch_bypass_counter[0]), .ZN(n49) );
  INVD3BWP30P140LVT U21 ( .I(n1), .ZN(prefetch_bypass_valid) );
  INVD1BWP30P140LVT U22 ( .I(n62), .ZN(n1) );
  NR2D1BWP30P140LVT U23 ( .A1(prefetch_bypass_counter[0]), .A2(N64), .ZN(N65)
         );
  INVD1BWP30P140LVT U24 ( .I(prefetch_bypass_counter[3]), .ZN(n3) );
  INVD1BWP30P140LVT U25 ( .I(prefetch_bypass_counter[2]), .ZN(n50) );
  OAI22D1BWP30P140LVT U26 ( .A1(prefetch_bypass_cycles[2]), .A2(n50), .B1(
        prefetch_bypass_cycles[3]), .B2(n3), .ZN(n2) );
  AOI221D1BWP30P140LVT U27 ( .A1(n3), .A2(prefetch_bypass_cycles[3]), .B1(n50), 
        .B2(prefetch_bypass_cycles[2]), .C(n2), .ZN(n10) );
  INVD1BWP30P140LVT U28 ( .I(prefetch_bypass_counter[1]), .ZN(n6) );
  INVD1BWP30P140LVT U29 ( .I(prefetch_bypass_counter[0]), .ZN(n5) );
  OAI22D1BWP30P140LVT U30 ( .A1(prefetch_bypass_cycles[0]), .A2(n5), .B1(
        prefetch_bypass_cycles[1]), .B2(n6), .ZN(n4) );
  AOI221D1BWP30P140LVT U31 ( .A1(n6), .A2(prefetch_bypass_cycles[1]), .B1(n5), 
        .B2(prefetch_bypass_cycles[0]), .C(n4), .ZN(n9) );
  INVD1BWP30P140LVT U32 ( .I(prefetch_bypass_counter[6]), .ZN(n56) );
  INVD1BWP30P140LVT U33 ( .I(prefetch_bypass_counter[7]), .ZN(n58) );
  OAI22D1BWP30P140LVT U34 ( .A1(prefetch_bypass_cycles[7]), .A2(n58), .B1(
        prefetch_bypass_cycles[6]), .B2(n56), .ZN(n7) );
  AOI221D1BWP30P140LVT U35 ( .A1(n56), .A2(prefetch_bypass_cycles[6]), .B1(n58), .B2(prefetch_bypass_cycles[7]), .C(n7), .ZN(n8) );
  AN4D1BWP30P140LVT U36 ( .A1(n10), .A2(n9), .A3(prefetch_bypass_valid), .A4(
        n8), .Z(n48) );
  INVD1BWP30P140LVT U37 ( .I(prefetch_bypass_counter[5]), .ZN(n12) );
  OAI22D1BWP30P140LVT U38 ( .A1(prefetch_bypass_cycles[4]), .A2(n53), .B1(
        prefetch_bypass_cycles[5]), .B2(n12), .ZN(n11) );
  AOI221D1BWP30P140LVT U39 ( .A1(n12), .A2(prefetch_bypass_cycles[5]), .B1(n53), .B2(prefetch_bypass_cycles[4]), .C(n11), .ZN(n47) );
  INVD2BWP30P140LVT U40 ( .I(prefetch_bypass_start_addr[13]), .ZN(n14) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n14), .A2(local_controller_id[5]), .Z(n17) );
  INVD1BWP30P140LVT U42 ( .I(sample_address[6]), .ZN(n13) );
  CKAN2D1BWP30P140LVT U43 ( .A1(prefetch_bypass_start_addr[6]), .A2(n13), .Z(
        n16) );
  OAI22D1BWP30P140LVT U44 ( .A1(n14), .A2(local_controller_id[5]), .B1(n13), 
        .B2(prefetch_bypass_start_addr[6]), .ZN(n15) );
  NR3D0P7BWP30P140LVT U45 ( .A1(n17), .A2(n16), .A3(n15), .ZN(n20) );
  XNR2UD1BWP30P140LVT U46 ( .A1(sample_address[7]), .A2(
        prefetch_bypass_start_addr[7]), .ZN(n19) );
  INVD1BWP30P140LVT U47 ( .I(sample_address[3]), .ZN(n22) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n22), .A2(prefetch_bypass_start_addr[3]), .Z(
        n25) );
  INVD1BWP30P140LVT U49 ( .I(sample_address[5]), .ZN(n21) );
  CKAN2D1BWP30P140LVT U50 ( .A1(prefetch_bypass_start_addr[5]), .A2(n21), .Z(
        n24) );
  OAI22D1BWP30P140LVT U51 ( .A1(n22), .A2(prefetch_bypass_start_addr[3]), .B1(
        n21), .B2(prefetch_bypass_start_addr[5]), .ZN(n23) );
  OR3D1BWP30P140LVT U52 ( .A1(n25), .A2(n24), .A3(n23), .Z(n40) );
  INVD1BWP30P140LVT U53 ( .I(sample_address[2]), .ZN(n28) );
  INVD1BWP30P140LVT U54 ( .I(sample_address[0]), .ZN(n27) );
  OAI22D1BWP30P140LVT U55 ( .A1(n28), .A2(prefetch_bypass_start_addr[2]), .B1(
        n27), .B2(prefetch_bypass_start_addr[0]), .ZN(n26) );
  AOI221D1BWP30P140LVT U56 ( .A1(n28), .A2(prefetch_bypass_start_addr[2]), 
        .B1(prefetch_bypass_start_addr[0]), .B2(n27), .C(n26), .ZN(n39) );
  INVD1BWP30P140LVT U57 ( .I(prefetch_bypass_start_addr[12]), .ZN(n30) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n30), .A2(local_controller_id[4]), .Z(n33) );
  INVD1BWP30P140LVT U59 ( .I(prefetch_bypass_start_addr[11]), .ZN(n29) );
  CKAN2D1BWP30P140LVT U60 ( .A1(local_controller_id[3]), .A2(n29), .Z(n32) );
  OAI22D1BWP30P140LVT U61 ( .A1(n30), .A2(local_controller_id[4]), .B1(n29), 
        .B2(local_controller_id[3]), .ZN(n31) );
  INVD1BWP30P140LVT U62 ( .I(sample_address[1]), .ZN(n36) );
  NR4D1BWP30P140LVT U63 ( .A1(n44), .A2(n43), .A3(n42), .A4(n41), .ZN(n45) );
  OAI21D2BWP30P140LVT U64 ( .A1(prefetch_bypass_valid), .A2(n45), .B(start), 
        .ZN(n46) );
  AOI211OPTREPBD2BWP30P140LVT U65 ( .A1(n48), .A2(n47), .B(n46), .C(reset), 
        .ZN(N73) );
  OA211D1BWP30P140LVT U66 ( .A1(prefetch_bypass_counter[1]), .A2(
        prefetch_bypass_counter[0]), .B(n49), .C(N73), .Z(N66) );
  AOI211D1BWP30P140LVT U67 ( .A1(n50), .A2(n49), .B(n51), .C(N64), .ZN(N67) );
  OA211D1BWP30P140LVT U68 ( .A1(prefetch_bypass_counter[3]), .A2(n51), .B(N73), 
        .C(n52), .Z(N68) );
  AOI211D1BWP30P140LVT U69 ( .A1(n53), .A2(n52), .B(n54), .C(N64), .ZN(N69) );
  OA211D1BWP30P140LVT U70 ( .A1(prefetch_bypass_counter[5]), .A2(n54), .B(N73), 
        .C(n55), .Z(N70) );
  AOI211D1BWP30P140LVT U71 ( .A1(n56), .A2(n55), .B(n59), .C(N64), .ZN(N71) );
  INVD1BWP30P140LVT U72 ( .I(n59), .ZN(n57) );
  AOI221D1BWP30P140LVT U73 ( .A1(prefetch_bypass_counter[7]), .A2(n59), .B1(
        n58), .B2(n57), .C(N64), .ZN(N72) );
endmodule


module global_controller ( CLK, reset, boot_up, start, table_parse, 
        input_valid, glob_scen_noc_input_valid, delay_matrix_element, 
        obj_id_element, from_glob_prefetch_start, from_glob_prefetch_dest, 
        scenario_update, local_controller_id, tapping_loc_packet, 
        from_glob_prefetch_stop, hardware_latency1, hardware_latency2, 
        scenario_len, prefetch_bypass_dest_addr_int, prefetch_bypass_cycles, 
        prefetch_bypass_start_addr, addr, data_in, h_tree_input_data, 
        h_tree_input_addr, prefetch_bypass_path_input_data, 
        prefetch_bypass_path_input_addr, prefetch_bypass_valid );
  input [13:0] delay_matrix_element;
  input [1:0] obj_id_element;
  output [7:0] from_glob_prefetch_start;
  output [3:0] from_glob_prefetch_dest;
  output [5:0] local_controller_id;
  output [9:0] tapping_loc_packet;
  output [7:0] from_glob_prefetch_stop;
  input [13:0] hardware_latency1;
  input [13:0] hardware_latency2;
  input [10:0] scenario_len;
  output [3:0] prefetch_bypass_dest_addr_int;
  output [7:0] prefetch_bypass_cycles;
  output [13:0] prefetch_bypass_start_addr;
  output [5:0] addr;
  input [31:0] data_in;
  output [31:0] h_tree_input_data;
  output [5:0] h_tree_input_addr;
  output [31:0] prefetch_bypass_path_input_data;
  output [3:0] prefetch_bypass_path_input_addr;
  input CLK, reset, boot_up, start, table_parse, input_valid,
         glob_scen_noc_input_valid, scenario_update;
  output prefetch_bypass_valid;
  wire   n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, N38, N39,
         N42, N45, N48, N51, N54, N57, N60, N63, N66, N69, N72, N75, N78, N81,
         N84, N87, N90, N93, N96, N99, N102, N105, N108, N111, N114, N117,
         N120, N123, N126, N129, N132, N135, N138, N141, N144, N147, N150,
         N151, n79, n80, n82, n123;
  wire   [7:0] counter_up;
  tri   [31:0] h_tree_input_data;
  tri   [5:0] h_tree_input_addr;
  tri   [31:0] prefetch_bypass_path_input_data;
  tri   [3:0] prefetch_bypass_path_input_addr;

  table_parse_engine dut_parse_engine ( .CLK(CLK), .reset(reset), .boot_up(
        boot_up), .table_parse(table_parse), .input_valid(input_valid), 
        .glob_scen_noc_input_valid(glob_scen_noc_input_valid), 
        .delay_matrix_element(delay_matrix_element), .obj_id_element(
        obj_id_element), .local_controller_id({n136, n137, n138, n139, n140, 
        n141}), .calc_global_controller_prefetch_start({n124, n125, n126, n127, 
        n128, n129, n130, n131}), .calc_glob_dest_addr({n132, n133, n134, n135}), .tapping_loc_packet({n142, n143, n144, n145, n146, n147, n148, n149, n150, 
        n151}), .calc_glob_prefetch_stop({n152, n153, n154, n155, n156, n157, 
        n158, n159}), .scenario_update(scenario_update), .hardware_latency1(
        hardware_latency1), .hardware_latency2(hardware_latency2), 
        .scenario_len(scenario_len), .prefetch_bypass_dest_addr_int(
        prefetch_bypass_dest_addr_int), .prefetch_bypass_cycles(
        prefetch_bypass_cycles), .prefetch_bypass_start_addr({
        prefetch_bypass_start_addr[13], n160, prefetch_bypass_start_addr[11:6], 
        n161, prefetch_bypass_start_addr[4], n162, n163, n164, 
        prefetch_bypass_start_addr[0]}) );
  addrGen dut_addr_gen ( .CLK(CLK), .rst(reset), .start(start), .addr({addr[5], 
        n165, addr[3:1], n166}), .counter_up(counter_up) );
  prefetch_bypass_module dut_prefetch_bypass ( .CLK(CLK), .reset(reset), 
        .start(start), .prefetch_bypass_dest_addr_int(
        prefetch_bypass_dest_addr_int), .prefetch_bypass_cycles(
        prefetch_bypass_cycles), .prefetch_bypass_start_addr({
        prefetch_bypass_start_addr[13], n160, prefetch_bypass_start_addr[11:6], 
        n161, prefetch_bypass_start_addr[4], n162, n163, 
        prefetch_bypass_start_addr[1:0]}), .local_controller_id({addr[5], n165, 
        addr[3:1], n166}), .sample_address(counter_up), .data_in(data_in), 
        .prefetch_bypass_path_input_data(prefetch_bypass_path_input_data), 
        .prefetch_bypass_path_input_addr(prefetch_bypass_path_input_addr), 
        .prefetch_bypass_valid(prefetch_bypass_valid) );
  DFQD1BWP30P140LVT h_tree_input_addr_reg_5_ ( .D(addr[5]), .CP(CLK), .Q(N39)
         );
  DFQD1BWP30P140LVT h_tree_input_addr_reg_2_ ( .D(addr[2]), .CP(CLK), .Q(N48)
         );
  DFQD1BWP30P140LVT h_tree_input_addr_reg_1_ ( .D(addr[1]), .CP(CLK), .Q(N51)
         );
  DFQD1BWP30P140LVT h_tree_input_data_reg_31_ ( .D(data_in[31]), .CP(CLK), .Q(
        N57) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_30_ ( .D(data_in[30]), .CP(CLK), .Q(
        N60) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_29_ ( .D(data_in[29]), .CP(CLK), .Q(
        N63) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_28_ ( .D(data_in[28]), .CP(CLK), .Q(
        N66) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_27_ ( .D(data_in[27]), .CP(CLK), .Q(
        N69) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_26_ ( .D(data_in[26]), .CP(CLK), .Q(
        N72) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_25_ ( .D(data_in[25]), .CP(CLK), .Q(
        N75) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_24_ ( .D(data_in[24]), .CP(CLK), .Q(
        N78) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_23_ ( .D(data_in[23]), .CP(CLK), .Q(
        N81) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_22_ ( .D(data_in[22]), .CP(CLK), .Q(
        N84) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_21_ ( .D(data_in[21]), .CP(CLK), .Q(
        N87) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_20_ ( .D(data_in[20]), .CP(CLK), .Q(
        N90) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_19_ ( .D(data_in[19]), .CP(CLK), .Q(
        N93) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_18_ ( .D(data_in[18]), .CP(CLK), .Q(
        N96) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_17_ ( .D(data_in[17]), .CP(CLK), .Q(
        N99) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_16_ ( .D(data_in[16]), .CP(CLK), .Q(
        N102) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_15_ ( .D(data_in[15]), .CP(CLK), .Q(
        N105) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_14_ ( .D(data_in[14]), .CP(CLK), .Q(
        N108) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_13_ ( .D(data_in[13]), .CP(CLK), .Q(
        N111) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_12_ ( .D(data_in[12]), .CP(CLK), .Q(
        N114) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_11_ ( .D(data_in[11]), .CP(CLK), .Q(
        N117) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_10_ ( .D(data_in[10]), .CP(CLK), .Q(
        N120) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_9_ ( .D(data_in[9]), .CP(CLK), .Q(
        N123) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_8_ ( .D(data_in[8]), .CP(CLK), .Q(
        N126) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_7_ ( .D(data_in[7]), .CP(CLK), .Q(
        N129) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_6_ ( .D(data_in[6]), .CP(CLK), .Q(
        N132) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_5_ ( .D(data_in[5]), .CP(CLK), .Q(
        N135) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_4_ ( .D(data_in[4]), .CP(CLK), .Q(
        N138) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_3_ ( .D(data_in[3]), .CP(CLK), .Q(
        N141) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_2_ ( .D(data_in[2]), .CP(CLK), .Q(
        N144) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_1_ ( .D(data_in[1]), .CP(CLK), .Q(
        N147) );
  DFQD1BWP30P140LVT h_tree_input_data_reg_0_ ( .D(data_in[0]), .CP(CLK), .Q(
        N150) );
  DFQD1BWP30P140LVT h_tree_input_data_tri_enable_reg_0_ ( .D(N38), .CP(CLK), 
        .Q(N151) );
  DFQD1BWP30P140LVT h_tree_input_addr_reg_0_ ( .D(addr[0]), .CP(CLK), .Q(N54)
         );
  DFQD1BWP30P140LVT h_tree_input_addr_reg_4_ ( .D(addr[4]), .CP(CLK), .Q(N42)
         );
  DFQD1BWP30P140LVT h_tree_input_addr_reg_3_ ( .D(addr[3]), .CP(CLK), .Q(N45)
         );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_1_ ( .I(N147), .OE(n82), .Z(
        h_tree_input_data[1]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_14_ ( .I(N108), .OE(n82), .Z(
        h_tree_input_data[14]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_15_ ( .I(N105), .OE(n82), .Z(
        h_tree_input_data[15]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_16_ ( .I(N102), .OE(n82), .Z(
        h_tree_input_data[16]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_17_ ( .I(N99), .OE(n82), .Z(
        h_tree_input_data[17]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_18_ ( .I(N96), .OE(n82), .Z(
        h_tree_input_data[18]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_19_ ( .I(N93), .OE(n82), .Z(
        h_tree_input_data[19]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_20_ ( .I(N90), .OE(n82), .Z(
        h_tree_input_data[20]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_21_ ( .I(N87), .OE(n82), .Z(
        h_tree_input_data[21]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_22_ ( .I(N84), .OE(n82), .Z(
        h_tree_input_data[22]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_23_ ( .I(N81), .OE(n82), .Z(
        h_tree_input_data[23]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_24_ ( .I(N78), .OE(n82), .Z(
        h_tree_input_data[24]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_25_ ( .I(N75), .OE(n82), .Z(
        h_tree_input_data[25]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_0_ ( .I(N150), .OE(n123), .Z(
        h_tree_input_data[0]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_2_ ( .I(N144), .OE(n123), .Z(
        h_tree_input_data[2]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_3_ ( .I(N141), .OE(n123), .Z(
        h_tree_input_data[3]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_4_ ( .I(N138), .OE(n123), .Z(
        h_tree_input_data[4]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_5_ ( .I(N135), .OE(n123), .Z(
        h_tree_input_data[5]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_6_ ( .I(N132), .OE(n123), .Z(
        h_tree_input_data[6]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_7_ ( .I(N129), .OE(n123), .Z(
        h_tree_input_data[7]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_8_ ( .I(N126), .OE(n123), .Z(
        h_tree_input_data[8]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_9_ ( .I(N123), .OE(n123), .Z(
        h_tree_input_data[9]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_10_ ( .I(N120), .OE(n123), .Z(
        h_tree_input_data[10]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_11_ ( .I(N117), .OE(n123), .Z(
        h_tree_input_data[11]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_12_ ( .I(N114), .OE(n123), .Z(
        h_tree_input_data[12]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_13_ ( .I(N111), .OE(n123), .Z(
        h_tree_input_data[13]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_26_ ( .I(N72), .OE(n82), .Z(
        h_tree_input_data[26]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_27_ ( .I(N69), .OE(n123), .Z(
        h_tree_input_data[27]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_28_ ( .I(N66), .OE(n82), .Z(
        h_tree_input_data[28]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_29_ ( .I(N63), .OE(n123), .Z(
        h_tree_input_data[29]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_30_ ( .I(N60), .OE(n82), .Z(
        h_tree_input_data[30]) );
  BUFTD4BWP30P140LVT h_tree_input_data_tri_31_ ( .I(N57), .OE(n123), .Z(
        h_tree_input_data[31]) );
  BUFTD4BWP30P140LVT h_tree_input_addr_tri_0_ ( .I(N54), .OE(n82), .Z(
        h_tree_input_addr[0]) );
  BUFTD4BWP30P140LVT h_tree_input_addr_tri_1_ ( .I(N51), .OE(n123), .Z(
        h_tree_input_addr[1]) );
  BUFTD4BWP30P140LVT h_tree_input_addr_tri_2_ ( .I(N48), .OE(n82), .Z(
        h_tree_input_addr[2]) );
  BUFTD4BWP30P140LVT h_tree_input_addr_tri_3_ ( .I(N45), .OE(n123), .Z(
        h_tree_input_addr[3]) );
  BUFTD4BWP30P140LVT h_tree_input_addr_tri_4_ ( .I(N42), .OE(n82), .Z(
        h_tree_input_addr[4]) );
  BUFTD4BWP30P140LVT h_tree_input_addr_tri_5_ ( .I(N39), .OE(n123), .Z(
        h_tree_input_addr[5]) );
  BUFFD4BWP30P140LVT U5 ( .I(n165), .Z(addr[4]) );
  BUFFD2BWP30P140LVT U6 ( .I(n166), .Z(addr[0]) );
  INVD1BWP30P140LVT U7 ( .I(n164), .ZN(n79) );
  INVD1BWP30P140LVT U8 ( .I(n160), .ZN(n80) );
  INVD8BWP30P140LVT U9 ( .I(n79), .ZN(prefetch_bypass_start_addr[1]) );
  INVD2BWP30P140LVT U10 ( .I(n80), .ZN(prefetch_bypass_start_addr[12]) );
  BUFFD2BWP30P140LVT U11 ( .I(n124), .Z(from_glob_prefetch_start[7]) );
  BUFFD2BWP30P140LVT U12 ( .I(n158), .Z(from_glob_prefetch_stop[1]) );
  BUFFD2BWP30P140LVT U13 ( .I(n157), .Z(from_glob_prefetch_stop[2]) );
  BUFFD2BWP30P140LVT U14 ( .I(n156), .Z(from_glob_prefetch_stop[3]) );
  BUFFD2BWP30P140LVT U15 ( .I(n155), .Z(from_glob_prefetch_stop[4]) );
  BUFFD2BWP30P140LVT U16 ( .I(n154), .Z(from_glob_prefetch_stop[5]) );
  BUFFD2BWP30P140LVT U17 ( .I(n153), .Z(from_glob_prefetch_stop[6]) );
  BUFFD2BWP30P140LVT U18 ( .I(n152), .Z(from_glob_prefetch_stop[7]) );
  BUFFD2BWP30P140LVT U19 ( .I(n151), .Z(tapping_loc_packet[0]) );
  BUFFD2BWP30P140LVT U20 ( .I(n150), .Z(tapping_loc_packet[1]) );
  BUFFD2BWP30P140LVT U21 ( .I(n149), .Z(tapping_loc_packet[2]) );
  BUFFD2BWP30P140LVT U22 ( .I(n148), .Z(tapping_loc_packet[3]) );
  BUFFD2BWP30P140LVT U23 ( .I(n147), .Z(tapping_loc_packet[4]) );
  BUFFD2BWP30P140LVT U24 ( .I(n146), .Z(tapping_loc_packet[5]) );
  BUFFD2BWP30P140LVT U25 ( .I(n145), .Z(tapping_loc_packet[6]) );
  BUFFD2BWP30P140LVT U26 ( .I(n144), .Z(tapping_loc_packet[7]) );
  BUFFD2BWP30P140LVT U27 ( .I(n143), .Z(tapping_loc_packet[8]) );
  BUFFD2BWP30P140LVT U28 ( .I(n142), .Z(tapping_loc_packet[9]) );
  BUFFD2BWP30P140LVT U29 ( .I(n141), .Z(local_controller_id[0]) );
  BUFFD2BWP30P140LVT U30 ( .I(n159), .Z(from_glob_prefetch_stop[0]) );
  BUFFD2BWP30P140LVT U31 ( .I(n140), .Z(local_controller_id[1]) );
  BUFFD2BWP30P140LVT U32 ( .I(n139), .Z(local_controller_id[2]) );
  BUFFD2BWP30P140LVT U33 ( .I(n138), .Z(local_controller_id[3]) );
  BUFFD2BWP30P140LVT U34 ( .I(n137), .Z(local_controller_id[4]) );
  BUFFD2BWP30P140LVT U35 ( .I(n136), .Z(local_controller_id[5]) );
  BUFFD2BWP30P140LVT U36 ( .I(n135), .Z(from_glob_prefetch_dest[0]) );
  BUFFD2BWP30P140LVT U37 ( .I(n134), .Z(from_glob_prefetch_dest[1]) );
  BUFFD2BWP30P140LVT U38 ( .I(n133), .Z(from_glob_prefetch_dest[2]) );
  BUFFD2BWP30P140LVT U39 ( .I(n125), .Z(from_glob_prefetch_start[6]) );
  BUFFD2BWP30P140LVT U40 ( .I(n132), .Z(from_glob_prefetch_dest[3]) );
  BUFFD2BWP30P140LVT U41 ( .I(n131), .Z(from_glob_prefetch_start[0]) );
  BUFFD2BWP30P140LVT U42 ( .I(n130), .Z(from_glob_prefetch_start[1]) );
  BUFFD2BWP30P140LVT U43 ( .I(n129), .Z(from_glob_prefetch_start[2]) );
  BUFFD2BWP30P140LVT U44 ( .I(n128), .Z(from_glob_prefetch_start[3]) );
  BUFFD2BWP30P140LVT U45 ( .I(n127), .Z(from_glob_prefetch_start[4]) );
  BUFFD2BWP30P140LVT U46 ( .I(n126), .Z(from_glob_prefetch_start[5]) );
  BUFFD2BWP30P140LVT U47 ( .I(n161), .Z(prefetch_bypass_start_addr[5]) );
  BUFFD2BWP30P140LVT U48 ( .I(n162), .Z(prefetch_bypass_start_addr[3]) );
  BUFFD2BWP30P140LVT U49 ( .I(n163), .Z(prefetch_bypass_start_addr[2]) );
  INVD2BWP30P140LVT U50 ( .I(N151), .ZN(n123) );
  INVD2BWP30P140LVT U51 ( .I(N151), .ZN(n82) );
  IND2D1BWP30P140LVT U52 ( .A1(reset), .B1(start), .ZN(N38) );
endmodule

