`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////////////////////
// Company: Gatech	
// Engineer: Mandovi Mukherjee
// 
// Create Date: 01/08/2021 
// System Name: accelerator
// Module Name: local controller
// Project Name: ARION DRBE
// Description: fetch and push data out to network; assuming the output from
// global controller comes in the form of a packet
// Dependencies:
// Additional Comments: 
/////////////////////////////////////////////////////////////////////////////////////////////////////

module only_controller_prefetch_full(CLK, reset,  from_glob_controller_delay,  input_boundary_flag, prev_dest_address, from_glob_dest_addr, packet_out, boundary_next, dest_address, from_glob_controller_valid, D, write_flag, from_glob_prefetch_valid, from_glob_prefetch_start, from_glob_prefetch_stop, from_glob_prefetch_dest, prefetch_packet_out, write_boundary_next, input_write_boundary, prefetch_next_dest_addr, prefetch_next_stop_address, prefetch_boundary_prev, input_prefetch_boundary_flag, prefetch_stop_address, prefetch_dest_addr, scenario_update, data_from_sram,  A, sram_CEB, sram_WEB, sram_D, sram_BWEB);

    // parameter
    	parameter N_sample = 256;
	parameter datawidth = 16;
	parameter address_vector_width = 8; //can be 200 or 8: 8 for small tapeout
	parameter id_width = 4; // 16 local controllers in subscaled system
	parameter sample_address_width = 8; /// assuming 1024 rows and 64 columns: needs to change if arrangement is different
	parameter packet_width = 2*datawidth + address_vector_width;
	

//=== IO Ports ===//

     // Normal Mode Input
        input [31:0] D;

     // BIST Mode Input



    // input
    	input CLK; // system clock, generated by VCO
	input reset;	
	input from_glob_controller_valid;
	input input_boundary_flag;
	input input_prefetch_boundary_flag;
	input input_write_boundary;
	input [address_vector_width - 1:0] prev_dest_address;
	input [address_vector_width - 1:0] prefetch_next_dest_addr;
        input [address_vector_width - 1:0] prefetch_next_stop_address;
	input [address_vector_width - 1:0] from_glob_dest_addr;
	input [address_vector_width - 1:0] from_glob_prefetch_dest;
	input [sample_address_width - 1:0] from_glob_controller_delay;
	
        //input [sample_address_width-1:0] ext_sample_address_M;
	input write_flag;

	input from_glob_prefetch_valid;
	input [sample_address_width - 1:0] from_glob_prefetch_start;
	input [sample_address_width - 1:0] from_glob_prefetch_stop;
	input scenario_update;
    	input [2*datawidth - 1:0] data_from_sram;

    // output
        output reg [packet_width-1:0] packet_out;  
        output reg [packet_width-1:0] prefetch_packet_out;  
        output reg boundary_next;
        output reg write_boundary_next;
        output reg [address_vector_width - 1:0] dest_address;
        output reg prefetch_boundary_prev;
	output reg [address_vector_width - 1:0] prefetch_dest_addr;
    	output reg [sample_address_width - 1:0] prefetch_stop_address;
    	//output reg BIST;
    	//output reg AWT;
    	//output reg SLP;
    	//output reg SD;
	output reg [sample_address_width-1:0] A;
   	output reg sram_CEB;
    	output reg sram_WEB;
    	//output reg CEBM;
	output reg [2*datawidth - 1:0] sram_BWEB;
	output reg [2*datawidth - 1:0] sram_D;
	//output [sample_address_width-1:0] AM;


//////////// internal status regs/signals //////////////////////////////////
    //reg [packet_width-1:0] packet_out_internal;
    reg coeff_num;

    reg [2*datawidth - 1:0] packet_out_data;
    reg [sample_address_width:0] sample_address;	
    reg [sample_address_width-1:0] sample_address_M;
    reg [sample_address_width:0] prefetch_sample_address;
    reg prefetch_reqd;



    reg CEB;
    reg WEB;
    reg [2*datawidth - 1:0] BWEB;
    reg prefetch_CEB;
    reg write_CEB;

    reg [sample_address_width-1:0] final_sample_address;	
    reg [sample_address_width-1:0] write_sample_address;	



    wire CLK_n;
    reg int_write_flag;
    reg internal_boundary_next;
    reg ready0;
    reg ready1;
    reg ready2;
    reg prefetch_ready1;
    reg [1:0] prefetch_ready_counter;
    reg coeff_num_next;
    reg [sample_address_width - 1:0] next_scen_start_addr;
    reg scen_ready0;
    reg scen_ready1;
    reg scen_ready2;
    reg scen_ready3;
    reg scen_change;
    reg [address_vector_width - 1:0] next_scen_prefetch_dest;


///////////////////////////////////////////////////////////////////////////////    

////////// logic part ///////////////////////////////////////////////////////  


    //assign packet_out = packet_out_internal;
    //assign CLK_n = ~CLK;
    //assign A = int_write_flag ? write_sample_address :  final_sample_address;
    //assign AM = write_flag ? ext_sample_address_M : sample_address_M;
    //assign prefetch_ready1 = 0; 
    //assign sram_CEB = int_write_flag ? write_CEB : (CEB & prefetch_CEB);


////////////sequential logic
//
//

   always @(posedge CLK_n) begin
	if (int_write_flag) sram_CEB <= write_CEB;
	else if (prefetch_ready_counter[0] | prefetch_ready_counter[1] | prefetch_ready1) sram_CEB <= prefetch_CEB;
	else sram_CEB <= CEB;

   end

   always @(posedge CLK_n) begin
	if (int_write_flag) sram_WEB <= WEB;
	else sram_WEB <= 1;
   end
   always @(posedge CLK_n) begin
	if (int_write_flag) sram_BWEB <= BWEB;
	else sram_BWEB <= 32'hffffffff;

   end



   always @(posedge CLK_n) begin
	if (int_write_flag) A <= write_sample_address;
	else A <= final_sample_address;


   end
   always @(posedge CLK_n) begin
	if (reset == 1 || scen_ready3 == 1) begin
		coeff_num_next <= 0;
		next_scen_start_addr <= 0;
		next_scen_prefetch_dest <= 0;
	end
	else if (from_glob_prefetch_valid == 1) begin
		coeff_num_next <= 1;
		next_scen_start_addr <= from_glob_prefetch_start;
		next_scen_prefetch_dest <= from_glob_prefetch_dest;
	end
	else begin
		coeff_num_next <= coeff_num_next;
		next_scen_start_addr <= next_scen_start_addr;
		next_scen_prefetch_dest <= next_scen_prefetch_dest;
	end

   end

   always @(posedge CLK_n) begin
	if (scenario_update) begin
     		scen_ready0 <= 1;
     		scen_ready1 <= 0;
     		scen_ready2 <= 0;
     		scen_ready3 <= 0;
		scen_change <= 1;

	end
	else if (scen_ready0) begin
     		scen_ready0 <= 0;
     		scen_ready1 <= 1;
     		scen_ready2 <= 0;
     		scen_ready3 <= 0;
		scen_change <= 1;

	end
	else if (scen_ready1) begin
     		scen_ready0 <= 0;
     		scen_ready1 <= 0;
     		scen_ready2 <= 1;
     		scen_ready3 <= 0;
		scen_change <= 1;

	end
	else if (scen_ready2) begin
     		scen_ready0 <= 0;
     		scen_ready1 <= 0;
     		scen_ready2 <= 0;
     		scen_ready3 <= 1;
		scen_change <= 1;

	end
	else if (scen_ready3) begin
     		scen_ready0 <= 0;
     		scen_ready1 <= 0;
     		scen_ready2 <= 0;
     		scen_ready3 <= 0;
		scen_change <= 1;

	end
	else    begin
     		scen_ready0 <= 0;
     		scen_ready1 <= 0;
     		scen_ready2 <= 0;
     		scen_ready3 <= 0;
		scen_change <= 0;

	end

   end


    always @(posedge CLK_n) begin
	if (reset == 1 || write_boundary_next == 1)  begin
		int_write_flag <= 0;
		if (write_boundary_next == 1) begin
			sram_D <= D;
		end
		else begin
			sram_D <= 0;
		end

		WEB <= 1;
		BWEB <= 32'hffffffff;
		write_CEB <= 1;
		write_sample_address <= 8'h0;
		write_boundary_next <= 0;


	end


	else begin
		if (write_flag == 1 || input_write_boundary == 1) begin
			int_write_flag <= 1;
			sram_D <= D;
			WEB <= 0;
			BWEB <= 0;
			write_CEB <= 0;
			if (write_sample_address == 8'hfe) begin
				write_boundary_next <= 1;

			end
			else begin
				write_boundary_next <= 0;

			end
			write_sample_address <= write_sample_address;
		end
		else if (int_write_flag == 1) begin
			int_write_flag <= 1;
			sram_D <= D;
			WEB <= 0;
			BWEB <= 0;
			write_CEB <= 0;
			if (write_sample_address == 8'hfe) begin
				write_boundary_next <= 1;

			end
			else if (write_sample_address == 8'hff) begin
				write_boundary_next <= 0;

			end
			else begin
				write_boundary_next <= 0;

			end
			write_sample_address <= write_sample_address + 1;
		end

		else begin
			int_write_flag <= 0;
			sram_D <= 0;
			WEB <= 1;
			BWEB <= 32'hffffffff;
			write_CEB <= 1;
			write_sample_address <= 8'h0;
			write_boundary_next <= 0;

		end
	end

    end




    always @ (posedge CLK_n) begin
        if (reset==1) begin

			sample_address <= 9'b0;
			sample_address_M <= 0;
			packet_out <= 40'bz;
			dest_address <= 0;
			coeff_num <= 0;
			boundary_next <= 0;
			internal_boundary_next <= 0;
			//BIST <= 0;
			//AWT <= 0;
			//SLP <= 0;
			//SD <= 0;
			CEB <= 1;
			//CEBM <= 1;
			ready0 <= 0;
			ready1 <= 0;
			ready2 <= 0;
			
        end

        else if (from_glob_controller_valid == 1 || input_boundary_flag == 1) begin
			packet_out <= 40'bz;
			boundary_next <=0;
			internal_boundary_next <=0;
			if (from_glob_controller_valid == 1) begin
				sample_address <= {1'b0,from_glob_controller_delay};
				dest_address <= from_glob_dest_addr;
			end
			else begin
				sample_address <= sample_address + 1;
				dest_address <= prev_dest_address;
			end
			coeff_num <= 0;	
			sample_address_M <= 0;
                        //BIST <= 0;
			//AWT <= 0;
			//SLP <= 0;
			//SD <= 0;
			CEB <= 0;
			//CEBM <= 1;
			ready0 <= 0;
			ready1 <= 1;
			ready2 <= 0;


	end
        else if (ready0 == 1 || ready1 == 1 || ready2 == 1) begin
			packet_out <= 40'bz;
			boundary_next <=0;
			internal_boundary_next <=0;
			sample_address <= sample_address + 1;
			dest_address <= dest_address;

			sample_address_M <= 0;
                        //BIST <= 0;
			//AWT <= 0;
			//SLP <= 0;
			//SD <= 0;
			CEB <= 0;
			//CEBM <= 1;
			if (ready0 == 1) begin
				ready0 <= 0;
				ready1 <= 1;
				ready2 <= 0;
				coeff_num <= 0;	
			end

			else if (ready1 == 1) begin
				ready0 <= 0;
				ready1 <= 0;
				ready2 <= 1;
				coeff_num <= 0;	
			end
			else begin
				ready0 <= 0;
				ready1 <= 0;
				ready2 <= 0;
				coeff_num <= 1;
			end


	end


			

	else begin
			ready0 <= 0;
			ready1 <= 0;
			ready2 <= 0;
			if (coeff_num == 1 && scen_ready3 == 1) begin		// && write_flag == 0) begin
				packet_out <= {packet_out_data, dest_address};
				boundary_next <= 0;
				internal_boundary_next <= 0;
				if (coeff_num_next == 1) begin
					sample_address <= sample_address + 1;
					CEB <= 0;
					//CEBM <= 1;
					dest_address <= next_scen_prefetch_dest;
					coeff_num <= 1;
				end
				else begin
					sample_address <= 0;
					CEB <= 1;
					//CEBM <= 1;
					dest_address <= 0;
					coeff_num <= 0;
				end

			end
			else if (coeff_num == 1 && scen_ready0 == 1) begin		// && write_flag == 0) begin
				packet_out <= {packet_out_data, dest_address};
				boundary_next <= 0;
				internal_boundary_next <= 0;
				if (coeff_num_next == 1) begin
					sample_address <= {1'b0,next_scen_start_addr};
					CEB <= 0;
					//CEBM <= 1;
					dest_address <= dest_address;
					coeff_num <= 1;
				end
				else begin
					sample_address <= 0;
					CEB <= 0;
					//CEBM <= 1;
					dest_address <= dest_address;
					coeff_num <= 1;
				end

			end
			else if (coeff_num == 1 && (scen_ready1 == 1 || scen_ready2 == 1)) begin		// && write_flag == 0) begin
				packet_out <= {packet_out_data, dest_address};
				boundary_next <= 0;
				internal_boundary_next <= 0;
				if (coeff_num_next == 1) begin
					sample_address <= sample_address + 1;
					CEB <= 0;
					//CEBM <= 1;
					dest_address <= dest_address;
					coeff_num <= 1;
				end
				else begin
					sample_address <= 0;
					CEB <= 0;
					//CEBM <= 1;
					dest_address <= dest_address;
					coeff_num <= 1;
				end

			end


			else if (coeff_num == 1 && internal_boundary_next == 0) begin		// && write_flag == 0) begin
				packet_out <= {packet_out_data, dest_address};
				sample_address <= sample_address + 1;
				CEB <= 0;
				//CEBM <= 1;
				dest_address <= dest_address;
				coeff_num <= coeff_num;
				if (sample_address == 9'h0ff) begin
					boundary_next <= 1;
					internal_boundary_next <= internal_boundary_next;
				end
				else if (sample_address == 9'h100) begin
					boundary_next <= 0;
					internal_boundary_next <= internal_boundary_next;
				end

				else if (sample_address == 9'h101) begin
					boundary_next <= boundary_next;
					internal_boundary_next <= 1;
				end

				else begin
					boundary_next <= boundary_next;
					internal_boundary_next <= internal_boundary_next;
				end

			end
			else if (coeff_num == 1 && internal_boundary_next == 1) begin		// && write_flag == 0) begin
				packet_out <= {packet_out_data, dest_address};
				sample_address <= 9'h0;   /// should automatically go to 0th address
				CEB <= 1;
				//CEBM <= 1;
				dest_address <= dest_address;
				coeff_num <= 0;
				boundary_next <= boundary_next;
				internal_boundary_next <= 0;

			end
			else if (coeff_num == 0 && scen_ready0 == 1) begin		// && write_flag == 0) begin
				packet_out <= 40'bz;
				boundary_next <= 0;
				internal_boundary_next <= 0;
				if (coeff_num_next == 1) begin
					sample_address <= {1'b0,next_scen_start_addr};
					CEB <= 0;
					//CEBM <= 1;
					dest_address <= next_scen_prefetch_dest;
					coeff_num <= 0;
				end
				else begin
					sample_address <= 0;
					CEB <= 1;
					//CEBM <= 1;
					dest_address <= 0;
					coeff_num <= 0;
				end

			end
			else if (coeff_num == 0 && scen_ready1 == 1) begin		// && write_flag == 0) begin
				packet_out <= 40'bz;
				boundary_next <= 0;
				internal_boundary_next <= 0;
				if (coeff_num_next == 1) begin
					sample_address <= sample_address + 1;
					CEB <= 0;
					//CEBM <= 1;
					dest_address <= dest_address;
					coeff_num <= 0;
				end
				else begin
					sample_address <= 0;
					CEB <= 1;
					//CEBM <= 1;
					dest_address <= 0;
					coeff_num <= 0;
				end

			end
			else if (coeff_num == 0 && scen_ready2 == 1) begin		// && write_flag == 0) begin
				packet_out <= 40'bz;
				boundary_next <= 0;
				internal_boundary_next <= 0;
				if (coeff_num_next == 1) begin
					sample_address <= sample_address + 1;
					CEB <= 0;
					//CEBM <= 1;
					dest_address <= dest_address;
					coeff_num <= 0;
				end
				else begin
					sample_address <= 0;
					CEB <= 1;
					//CEBM <= 1;
					dest_address <= 0;
					coeff_num <= 0;
				end

			end
			else if (coeff_num == 0 && scen_ready3 == 1) begin		// && write_flag == 0) begin
				packet_out <= 40'bz;
				boundary_next <= 0;
				internal_boundary_next <= 0;
				if (coeff_num_next == 1) begin
					sample_address <= sample_address + 1;
					CEB <= 0;
					//CEBM <= 1;
					dest_address <= dest_address;
					coeff_num <= 1;  ///difference from previous states
				end
				else begin
					sample_address <= 0;
					CEB <= 1;
					//CEBM <= 1;
					dest_address <= 0;
					coeff_num <= 0;
				end

			end





			else begin
				packet_out <= 40'bz;
				sample_address <= sample_address;
				dest_address <= dest_address;
				coeff_num <= coeff_num;
				boundary_next <= boundary_next;
				CEB <= 1;
				//CEBM <= 1;
				internal_boundary_next <= internal_boundary_next;

			end


			sample_address_M <= 0;
                        //BIST <= 0;
			//AWT <= 0;
			//SLP <= 0;
			//SD <= 0;

	end  
     end

     always @(posedge CLK_n) begin   //// merge with prev always block: prefetch sample address is assigned in both
        if (reset == 1 || scenario_update == 1) begin
		prefetch_sample_address <= 9'h0ff;
		prefetch_packet_out <= 40'bz;
		prefetch_reqd <= 0;
		prefetch_dest_addr <= 0;
		prefetch_stop_address <= 0;
		prefetch_CEB <= 1;
		prefetch_boundary_prev <= 0;
		prefetch_ready1 <= 0;
		prefetch_ready_counter <= 2'b0;

        end

	else if (from_glob_prefetch_valid == 1 || input_prefetch_boundary_flag == 1) begin
		prefetch_reqd <= 1;
		prefetch_CEB <= 1;
		prefetch_boundary_prev <= 0;
		prefetch_ready1 <= 0;
		prefetch_ready_counter <= 2'b0;
		prefetch_packet_out <= 40'bz;
		if (from_glob_prefetch_valid == 1) begin
			prefetch_dest_addr <= from_glob_prefetch_dest;
			prefetch_sample_address <= {1'b0,from_glob_prefetch_start};
			prefetch_stop_address <= from_glob_prefetch_stop;
		end
		else begin
			prefetch_dest_addr <= prefetch_next_dest_addr;
			prefetch_stop_address <= prefetch_next_stop_address;
			prefetch_sample_address <= 9'h0ff;
		end
	end

	else if (prefetch_boundary_prev == 1)  begin
		prefetch_dest_addr <= prefetch_dest_addr;
		prefetch_stop_address <= prefetch_stop_address;
		prefetch_packet_out <= 40'bz;
		prefetch_sample_address <= 9'h0ff;
		prefetch_reqd <= 0;
		prefetch_CEB <= 1;
		prefetch_boundary_prev <= 0;   ////check condition
		prefetch_ready1 <= 0;
		prefetch_ready_counter <= 2'b0;
	end
	else if (coeff_num == 0 && input_boundary_flag == 0 && ready1 == 0 & ready2 == 0 && int_write_flag==0 && input_write_boundary == 0 && prefetch_reqd == 1 ) begin
		prefetch_dest_addr <= prefetch_dest_addr;
		prefetch_stop_address <= prefetch_stop_address;
		if (prefetch_ready1 == 1) begin
			prefetch_reqd <= 1;
			prefetch_packet_out <= 40'bz;
			prefetch_sample_address <= prefetch_sample_address - 1; //might need to stop after 1 prefetch
			prefetch_CEB <= 0;
			prefetch_boundary_prev <= prefetch_boundary_prev;   ////check condition
			if (prefetch_ready_counter == 2'b10) begin
				prefetch_ready1 <= 0;
			end
			else begin
				prefetch_ready1 <= 1;
			end 
			prefetch_ready_counter <= prefetch_ready_counter + 1;
		end
		else if (prefetch_ready_counter == 2'b11) begin
			prefetch_packet_out <= {packet_out_data,prefetch_dest_addr};
			prefetch_sample_address <= prefetch_sample_address - 1; //might need to stop after 1 prefetch
			prefetch_ready1 <= prefetch_ready1;
			if (prefetch_sample_address[7:0] == prefetch_stop_address || prefetch_sample_address == 9'h1fd ) begin
				prefetch_reqd <= 0;
				prefetch_CEB <= 1;
				prefetch_ready_counter <= 2'b0;	
				if (prefetch_sample_address == 9'h1fd) begin  //add condition for stop address at boundary of SRAM
					prefetch_boundary_prev <= 1;
				end
				else begin	
					prefetch_boundary_prev <= 0;
				end

			end	
			else begin
				prefetch_reqd <= prefetch_reqd;
				prefetch_CEB <= 0;
				prefetch_boundary_prev <= 0;
				prefetch_ready_counter <= prefetch_ready_counter;
			end

		end
		else begin  ///check this branch
			prefetch_reqd <= prefetch_reqd;
			prefetch_packet_out <= 40'bz;
			prefetch_sample_address <= prefetch_sample_address; 
			prefetch_CEB <= 0;
			prefetch_boundary_prev <= prefetch_boundary_prev;   ////check condition
			prefetch_ready1 <= 1;
			prefetch_ready_counter <= 2'b0;

		end
	

	end
	else begin
		prefetch_dest_addr <= prefetch_dest_addr;
		prefetch_reqd <= prefetch_reqd;
		prefetch_stop_address <= prefetch_stop_address;
		prefetch_sample_address <= prefetch_sample_address;
		prefetch_packet_out <= 40'bz;
		prefetch_CEB <= prefetch_CEB;
		prefetch_boundary_prev <= prefetch_boundary_prev;
		prefetch_ready1 <= 0;
		prefetch_ready_counter <= 2'b0;
	end


     end


     always @(posedge CLK_n) begin
	if (prefetch_ready_counter[0] | prefetch_ready_counter[1] | prefetch_ready1) begin
		final_sample_address <= prefetch_sample_address[7:0];
	end
	else begin
		final_sample_address <= sample_address[7:0];
	end

     end


     always @(posedge CLK) begin
	packet_out_data <= data_from_sram;

     end


    INVD6BWP30P140LVT UI_342 ( .I(CLK), .ZN(CLK_n) );

//    TS1N28HPCPLVTB256X32M4SWBASO UI_dut_mem (.SLP(SLP), .SD(SD), .CLK(CLK), .CEB(sram_CEB), .WEB(sram_WEB), .CEBM(CEBM), .WEBM(WEBM), .AWT(AWT), .A(A), .D(sram_D), .BWEB(sram_BWEB), .AM(AM), .DM(DM), .BWEBM(BWEBM), .BIST(BIST), .Q(data_from_sram));

	 
	 


   
endmodule
    
