
module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_0 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n8, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(o_data_bus[2]) );
  DFD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(o_data_bus[8]) );
  DFD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(o_data_bus[9]) );
  DFD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  INVD3BWP30P140 U3 ( .I(n35), .ZN(n124) );
  NR2D4BWP30P140 U4 ( .A1(n31), .A2(n30), .ZN(n35) );
  NR2D1BWP30P140 U5 ( .A1(i_cmd[1]), .A2(n109), .ZN(n42) );
  INVD6BWP30P140 U6 ( .I(n45), .ZN(n1) );
  ND2OPTPAD1BWP30P140 U7 ( .A1(i_cmd[0]), .A2(n29), .ZN(n30) );
  MUX2NOPTD2BWP30P140 U8 ( .I0(i_valid[0]), .I1(i_valid[1]), .S(i_cmd[1]), 
        .ZN(n31) );
  MUX2NOPTD2BWP30P140 U9 ( .I0(i_valid[0]), .I1(i_valid[1]), .S(i_cmd[0]), 
        .ZN(n41) );
  OR2D8BWP30P140 U10 ( .A1(n32), .A2(i_cmd[0]), .Z(n126) );
  CKND2D4BWP30P140 U11 ( .A1(i_valid[0]), .A2(n29), .ZN(n32) );
  INVD1BWP30P140 U12 ( .I(n126), .ZN(n8) );
  INVD8BWP30P140 U13 ( .I(n126), .ZN(n145) );
  INVD1BWP30P140 U14 ( .I(n32), .ZN(n114) );
  INVD1BWP30P140 U15 ( .I(i_cmd[0]), .ZN(n112) );
  ND3OPTPAD2BWP30P140 U16 ( .A1(i_cmd[1]), .A2(i_valid[1]), .A3(n29), .ZN(n115) );
  ND2D1BWP30P140 U17 ( .A1(n28), .A2(i_en), .ZN(n109) );
  ND2D1BWP30P140 U18 ( .A1(n126), .A2(n113), .ZN(N353) );
  IND2D1BWP30P140 U19 ( .A1(n112), .B1(n111), .ZN(n113) );
  NR2D1BWP30P140 U20 ( .A1(n110), .A2(n109), .ZN(n111) );
  INVD1BWP30P140 U21 ( .I(i_valid[1]), .ZN(n110) );
  OAI21D1BWP30P140 U22 ( .A1(n124), .A2(n108), .B(n107), .ZN(N287) );
  OAI21D1BWP30P140 U23 ( .A1(n124), .A2(n106), .B(n105), .ZN(N288) );
  ND2D1BWP30P140 U24 ( .A1(n8), .A2(i_data_bus[1]), .ZN(n105) );
  OAI22D1BWP30P140 U25 ( .A1(n126), .A2(n77), .B1(n124), .B2(n36), .ZN(N292)
         );
  OAI22D1BWP30P140 U26 ( .A1(n147), .A2(n37), .B1(n126), .B2(n99), .ZN(N304)
         );
  OAI22D1BWP30P140 U27 ( .A1(n147), .A2(n38), .B1(n126), .B2(n101), .ZN(N305)
         );
  OAI22D1BWP30P140 U28 ( .A1(n147), .A2(n39), .B1(n126), .B2(n49), .ZN(N317)
         );
  OAI22D1BWP30P140 U29 ( .A1(n147), .A2(n40), .B1(n126), .B2(n104), .ZN(N318)
         );
  ND2D1BWP30P140 U30 ( .A1(n102), .A2(i_data_bus[47]), .ZN(n94) );
  ND2D1BWP30P140 U31 ( .A1(n102), .A2(i_data_bus[51]), .ZN(n54) );
  ND2D1BWP30P140 U32 ( .A1(n102), .A2(i_data_bus[52]), .ZN(n82) );
  ND2D1BWP30P140 U33 ( .A1(n102), .A2(i_data_bus[53]), .ZN(n80) );
  ND2D1BWP30P140 U34 ( .A1(n102), .A2(i_data_bus[54]), .ZN(n74) );
  ND2D1BWP30P140 U35 ( .A1(n102), .A2(i_data_bus[55]), .ZN(n72) );
  ND2D1BWP30P140 U36 ( .A1(n102), .A2(i_data_bus[56]), .ZN(n70) );
  ND2D1BWP30P140 U37 ( .A1(n102), .A2(i_data_bus[57]), .ZN(n68) );
  ND2D1BWP30P140 U38 ( .A1(n102), .A2(i_data_bus[58]), .ZN(n66) );
  ND2D1BWP30P140 U39 ( .A1(n102), .A2(i_data_bus[59]), .ZN(n58) );
  ND2D1BWP30P140 U40 ( .A1(n102), .A2(i_data_bus[60]), .ZN(n56) );
  ND2D1BWP30P140 U41 ( .A1(n102), .A2(i_data_bus[61]), .ZN(n46) );
  ND2D1BWP30P140 U42 ( .A1(n102), .A2(i_data_bus[62]), .ZN(n48) );
  ND2D1BWP30P140 U43 ( .A1(n102), .A2(i_data_bus[63]), .ZN(n103) );
  INR2D4BWP30P140 U44 ( .A1(n42), .B1(n41), .ZN(n45) );
  INVD1BWP30P140 U45 ( .I(n109), .ZN(n29) );
  INVD1BWP30P140 U46 ( .I(rst), .ZN(n28) );
  INVD6BWP30P140 U47 ( .I(n35), .ZN(n147) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[51]), .ZN(n33) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[19]), .ZN(n55) );
  OAI22D1BWP30P140 U50 ( .A1(n147), .A2(n33), .B1(n126), .B2(n55), .ZN(N306)
         );
  INVD1BWP30P140 U51 ( .I(i_data_bus[61]), .ZN(n34) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[29]), .ZN(n47) );
  OAI22D1BWP30P140 U53 ( .A1(n147), .A2(n34), .B1(n126), .B2(n47), .ZN(N316)
         );
  INVD1BWP30P140 U54 ( .I(i_data_bus[5]), .ZN(n77) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[37]), .ZN(n36) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[49]), .ZN(n37) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[17]), .ZN(n99) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[50]), .ZN(n38) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[18]), .ZN(n101) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[62]), .ZN(n39) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[30]), .ZN(n49) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[63]), .ZN(n40) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[31]), .ZN(n104) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[3]), .ZN(n125) );
  INVD6BWP30P140 U65 ( .I(n115), .ZN(n102) );
  ND2OPTIBD1BWP30P140 U66 ( .A1(n102), .A2(i_data_bus[35]), .ZN(n43) );
  OAI21D1BWP30P140 U67 ( .A1(n1), .A2(n125), .B(n43), .ZN(N322) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[4]), .ZN(n122) );
  ND2OPTIBD1BWP30P140 U69 ( .A1(n102), .A2(i_data_bus[36]), .ZN(n44) );
  OAI21D1BWP30P140 U70 ( .A1(n1), .A2(n122), .B(n44), .ZN(N323) );
  OAI21D1BWP30P140 U71 ( .A1(n1), .A2(n47), .B(n46), .ZN(N348) );
  OAI21D1BWP30P140 U72 ( .A1(n1), .A2(n49), .B(n48), .ZN(N349) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[9]), .ZN(n51) );
  ND2OPTIBD1BWP30P140 U74 ( .A1(n102), .A2(i_data_bus[41]), .ZN(n50) );
  OAI21D1BWP30P140 U75 ( .A1(n1), .A2(n51), .B(n50), .ZN(N328) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U77 ( .A1(n102), .A2(i_data_bus[32]), .ZN(n52) );
  OAI21D1BWP30P140 U78 ( .A1(n1), .A2(n53), .B(n52), .ZN(N319) );
  OAI21D1BWP30P140 U79 ( .A1(n1), .A2(n55), .B(n54), .ZN(N338) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[28]), .ZN(n57) );
  OAI21D1BWP30P140 U81 ( .A1(n1), .A2(n57), .B(n56), .ZN(N347) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[27]), .ZN(n59) );
  OAI21D1BWP30P140 U83 ( .A1(n1), .A2(n59), .B(n58), .ZN(N346) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[8]), .ZN(n61) );
  ND2OPTIBD1BWP30P140 U85 ( .A1(n102), .A2(i_data_bus[40]), .ZN(n60) );
  OAI21D1BWP30P140 U86 ( .A1(n1), .A2(n61), .B(n60), .ZN(N327) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[1]), .ZN(n63) );
  ND2OPTIBD1BWP30P140 U88 ( .A1(n102), .A2(i_data_bus[33]), .ZN(n62) );
  OAI21D1BWP30P140 U89 ( .A1(n1), .A2(n63), .B(n62), .ZN(N320) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[2]), .ZN(n65) );
  ND2OPTIBD1BWP30P140 U91 ( .A1(n102), .A2(i_data_bus[34]), .ZN(n64) );
  OAI21D1BWP30P140 U92 ( .A1(n1), .A2(n65), .B(n64), .ZN(N321) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[26]), .ZN(n67) );
  OAI21D1BWP30P140 U94 ( .A1(n1), .A2(n67), .B(n66), .ZN(N345) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[25]), .ZN(n69) );
  OAI21D1BWP30P140 U96 ( .A1(n1), .A2(n69), .B(n68), .ZN(N344) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[24]), .ZN(n71) );
  OAI21D1BWP30P140 U98 ( .A1(n1), .A2(n71), .B(n70), .ZN(N343) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[23]), .ZN(n73) );
  OAI21D1BWP30P140 U100 ( .A1(n1), .A2(n73), .B(n72), .ZN(N342) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[22]), .ZN(n75) );
  OAI21D1BWP30P140 U102 ( .A1(n1), .A2(n75), .B(n74), .ZN(N341) );
  ND2OPTIBD1BWP30P140 U103 ( .A1(n102), .A2(i_data_bus[37]), .ZN(n76) );
  OAI21D1BWP30P140 U104 ( .A1(n1), .A2(n77), .B(n76), .ZN(N324) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[6]), .ZN(n120) );
  ND2OPTIBD1BWP30P140 U106 ( .A1(n102), .A2(i_data_bus[38]), .ZN(n78) );
  OAI21D1BWP30P140 U107 ( .A1(n1), .A2(n120), .B(n78), .ZN(N325) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[7]), .ZN(n118) );
  ND2OPTIBD1BWP30P140 U109 ( .A1(n102), .A2(i_data_bus[39]), .ZN(n79) );
  OAI21D1BWP30P140 U110 ( .A1(n1), .A2(n118), .B(n79), .ZN(N326) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[21]), .ZN(n81) );
  OAI21D1BWP30P140 U112 ( .A1(n1), .A2(n81), .B(n80), .ZN(N340) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[20]), .ZN(n83) );
  OAI21D1BWP30P140 U114 ( .A1(n1), .A2(n83), .B(n82), .ZN(N339) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[10]), .ZN(n85) );
  ND2OPTIBD1BWP30P140 U116 ( .A1(n102), .A2(i_data_bus[42]), .ZN(n84) );
  OAI21D1BWP30P140 U117 ( .A1(n1), .A2(n85), .B(n84), .ZN(N329) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[11]), .ZN(n87) );
  ND2OPTIBD1BWP30P140 U119 ( .A1(n102), .A2(i_data_bus[43]), .ZN(n86) );
  OAI21D1BWP30P140 U120 ( .A1(n1), .A2(n87), .B(n86), .ZN(N330) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[12]), .ZN(n89) );
  ND2OPTIBD1BWP30P140 U122 ( .A1(n102), .A2(i_data_bus[44]), .ZN(n88) );
  OAI21D1BWP30P140 U123 ( .A1(n1), .A2(n89), .B(n88), .ZN(N331) );
  INVD1BWP30P140 U124 ( .I(i_data_bus[13]), .ZN(n91) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n102), .A2(i_data_bus[45]), .ZN(n90) );
  OAI21D1BWP30P140 U126 ( .A1(n1), .A2(n91), .B(n90), .ZN(N332) );
  INVD1BWP30P140 U127 ( .I(i_data_bus[14]), .ZN(n93) );
  ND2OPTIBD1BWP30P140 U128 ( .A1(n102), .A2(i_data_bus[46]), .ZN(n92) );
  OAI21D1BWP30P140 U129 ( .A1(n1), .A2(n93), .B(n92), .ZN(N333) );
  INVD1BWP30P140 U130 ( .I(i_data_bus[15]), .ZN(n95) );
  OAI21D1BWP30P140 U131 ( .A1(n1), .A2(n95), .B(n94), .ZN(N334) );
  INVD1BWP30P140 U132 ( .I(i_data_bus[16]), .ZN(n97) );
  ND2OPTIBD1BWP30P140 U133 ( .A1(n102), .A2(i_data_bus[48]), .ZN(n96) );
  OAI21D1BWP30P140 U134 ( .A1(n1), .A2(n97), .B(n96), .ZN(N335) );
  ND2OPTIBD1BWP30P140 U135 ( .A1(n102), .A2(i_data_bus[49]), .ZN(n98) );
  OAI21D1BWP30P140 U136 ( .A1(n1), .A2(n99), .B(n98), .ZN(N336) );
  ND2OPTIBD1BWP30P140 U137 ( .A1(n102), .A2(i_data_bus[50]), .ZN(n100) );
  OAI21D1BWP30P140 U138 ( .A1(n1), .A2(n101), .B(n100), .ZN(N337) );
  OAI21D1BWP30P140 U139 ( .A1(n1), .A2(n104), .B(n103), .ZN(N350) );
  INVD1BWP30P140 U140 ( .I(i_data_bus[33]), .ZN(n106) );
  INVD1BWP30P140 U141 ( .I(i_data_bus[32]), .ZN(n108) );
  IND2D2BWP30P140 U142 ( .A1(n126), .B1(i_data_bus[0]), .ZN(n107) );
  INVD1BWP30P140 U143 ( .I(n114), .ZN(n116) );
  OAI21D1BWP30P140 U144 ( .A1(n116), .A2(i_cmd[1]), .B(n115), .ZN(N354) );
  INVD1BWP30P140 U145 ( .I(i_data_bus[39]), .ZN(n117) );
  OAI22D1BWP30P140 U146 ( .A1(n126), .A2(n118), .B1(n124), .B2(n117), .ZN(N294) );
  INVD1BWP30P140 U147 ( .I(i_data_bus[38]), .ZN(n119) );
  OAI22D1BWP30P140 U148 ( .A1(n126), .A2(n120), .B1(n124), .B2(n119), .ZN(N293) );
  INVD1BWP30P140 U149 ( .I(i_data_bus[36]), .ZN(n121) );
  OAI22D1BWP30P140 U150 ( .A1(n126), .A2(n122), .B1(n124), .B2(n121), .ZN(N291) );
  INVD1BWP30P140 U151 ( .I(i_data_bus[35]), .ZN(n123) );
  OAI22D1BWP30P140 U152 ( .A1(n126), .A2(n125), .B1(n124), .B2(n123), .ZN(N290) );
  INVD1BWP30P140 U153 ( .I(i_data_bus[60]), .ZN(n127) );
  MOAI22D1BWP30P140 U154 ( .A1(n147), .A2(n127), .B1(n145), .B2(i_data_bus[28]), .ZN(N315) );
  INVD1BWP30P140 U155 ( .I(i_data_bus[48]), .ZN(n128) );
  MOAI22D1BWP30P140 U156 ( .A1(n147), .A2(n128), .B1(n145), .B2(i_data_bus[16]), .ZN(N303) );
  INVD1BWP30P140 U157 ( .I(i_data_bus[34]), .ZN(n129) );
  MOAI22D1BWP30P140 U158 ( .A1(n147), .A2(n129), .B1(n145), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140 U159 ( .I(i_data_bus[59]), .ZN(n130) );
  MOAI22D1BWP30P140 U160 ( .A1(n147), .A2(n130), .B1(n145), .B2(i_data_bus[27]), .ZN(N314) );
  INVD1BWP30P140 U161 ( .I(i_data_bus[47]), .ZN(n131) );
  MOAI22D1BWP30P140 U162 ( .A1(n147), .A2(n131), .B1(n145), .B2(i_data_bus[15]), .ZN(N302) );
  INVD1BWP30P140 U163 ( .I(i_data_bus[58]), .ZN(n132) );
  MOAI22D1BWP30P140 U164 ( .A1(n147), .A2(n132), .B1(n145), .B2(i_data_bus[26]), .ZN(N313) );
  INVD1BWP30P140 U165 ( .I(i_data_bus[46]), .ZN(n133) );
  MOAI22D1BWP30P140 U166 ( .A1(n147), .A2(n133), .B1(n145), .B2(i_data_bus[14]), .ZN(N301) );
  INVD1BWP30P140 U167 ( .I(i_data_bus[57]), .ZN(n134) );
  MOAI22D1BWP30P140 U168 ( .A1(n147), .A2(n134), .B1(n145), .B2(i_data_bus[25]), .ZN(N312) );
  INVD1BWP30P140 U169 ( .I(i_data_bus[45]), .ZN(n135) );
  MOAI22D1BWP30P140 U170 ( .A1(n147), .A2(n135), .B1(n145), .B2(i_data_bus[13]), .ZN(N300) );
  INVD1BWP30P140 U171 ( .I(i_data_bus[56]), .ZN(n136) );
  MOAI22D1BWP30P140 U172 ( .A1(n147), .A2(n136), .B1(n145), .B2(i_data_bus[24]), .ZN(N311) );
  INVD1BWP30P140 U173 ( .I(i_data_bus[44]), .ZN(n137) );
  MOAI22D1BWP30P140 U174 ( .A1(n147), .A2(n137), .B1(n145), .B2(i_data_bus[12]), .ZN(N299) );
  INVD1BWP30P140 U175 ( .I(i_data_bus[55]), .ZN(n138) );
  MOAI22D1BWP30P140 U176 ( .A1(n147), .A2(n138), .B1(n145), .B2(i_data_bus[23]), .ZN(N310) );
  INVD1BWP30P140 U177 ( .I(i_data_bus[43]), .ZN(n139) );
  MOAI22D1BWP30P140 U178 ( .A1(n147), .A2(n139), .B1(n145), .B2(i_data_bus[11]), .ZN(N298) );
  INVD1BWP30P140 U179 ( .I(i_data_bus[54]), .ZN(n140) );
  MOAI22D1BWP30P140 U180 ( .A1(n147), .A2(n140), .B1(n145), .B2(i_data_bus[22]), .ZN(N309) );
  INVD1BWP30P140 U181 ( .I(i_data_bus[42]), .ZN(n141) );
  MOAI22D1BWP30P140 U182 ( .A1(n147), .A2(n141), .B1(n145), .B2(i_data_bus[10]), .ZN(N297) );
  INVD1BWP30P140 U183 ( .I(i_data_bus[53]), .ZN(n142) );
  MOAI22D1BWP30P140 U184 ( .A1(n147), .A2(n142), .B1(n145), .B2(i_data_bus[21]), .ZN(N308) );
  INVD1BWP30P140 U185 ( .I(i_data_bus[41]), .ZN(n143) );
  MOAI22D1BWP30P140 U186 ( .A1(n147), .A2(n143), .B1(n145), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140 U187 ( .I(i_data_bus[52]), .ZN(n144) );
  MOAI22D1BWP30P140 U188 ( .A1(n147), .A2(n144), .B1(n145), .B2(i_data_bus[20]), .ZN(N307) );
  INVD1BWP30P140 U189 ( .I(i_data_bus[40]), .ZN(n146) );
  MOAI22D1BWP30P140 U190 ( .A1(n147), .A2(n146), .B1(n145), .B2(i_data_bus[8]), 
        .ZN(N295) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_1 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90;

  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n25), .Z(n88) );
  INR2D1BWP30P140 U4 ( .A1(i_cmd[1]), .B1(i_valid[1]), .ZN(n6) );
  NR2D1BWP30P140 U5 ( .A1(n48), .A2(i_cmd[1]), .ZN(n52) );
  INVD4BWP30P140 U6 ( .I(n10), .ZN(n1) );
  ND2OPTIBD1BWP30P140 U7 ( .A1(i_cmd[0]), .A2(n25), .ZN(n4) );
  NR2D1BWP30P140 U8 ( .A1(i_valid[0]), .A2(i_cmd[1]), .ZN(n5) );
  INVD1BWP30P140 U9 ( .I(n3), .ZN(n8) );
  ND2OPTIBD1BWP30P140 U10 ( .A1(n24), .A2(n23), .ZN(n3) );
  INVD1BWP30P140 U11 ( .I(i_valid[0]), .ZN(n50) );
  INVD1BWP30P140 U12 ( .I(n72), .ZN(n61) );
  ND2D1BWP30P140 U13 ( .A1(n2), .A2(i_en), .ZN(n48) );
  INVD1BWP30P140 U14 ( .I(i_cmd[0]), .ZN(n23) );
  OAI22D1BWP30P140 U15 ( .A1(n47), .A2(n64), .B1(n1), .B2(n7), .ZN(N297) );
  INVD1BWP30P140 U16 ( .I(n88), .ZN(n26) );
  INVD1BWP30P140 U17 ( .I(rst), .ZN(n2) );
  INR2D2BWP30P140 U18 ( .A1(i_valid[0]), .B1(n48), .ZN(n24) );
  INVD2BWP30P140 U19 ( .I(n8), .ZN(n47) );
  INVD1BWP30P140 U20 ( .I(i_data_bus[10]), .ZN(n64) );
  NR3D1BWP30P140 U21 ( .A1(n6), .A2(n5), .A3(n4), .ZN(n10) );
  INVD1BWP30P140 U22 ( .I(i_data_bus[42]), .ZN(n7) );
  INVD1BWP30P140 U23 ( .I(i_data_bus[51]), .ZN(n9) );
  INVD2BWP30P140 U24 ( .I(n8), .ZN(n22) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[19]), .ZN(n71) );
  OAI22D1BWP30P140 U26 ( .A1(n1), .A2(n9), .B1(n22), .B2(n71), .ZN(N306) );
  INVD1BWP30P140 U27 ( .I(i_data_bus[52]), .ZN(n11) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[20]), .ZN(n73) );
  OAI22D1BWP30P140 U29 ( .A1(n1), .A2(n11), .B1(n22), .B2(n73), .ZN(N307) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[53]), .ZN(n12) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[21]), .ZN(n74) );
  OAI22D1BWP30P140 U32 ( .A1(n1), .A2(n12), .B1(n22), .B2(n74), .ZN(N308) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[55]), .ZN(n13) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[23]), .ZN(n76) );
  OAI22D1BWP30P140 U35 ( .A1(n1), .A2(n13), .B1(n22), .B2(n76), .ZN(N310) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[57]), .ZN(n14) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[25]), .ZN(n85) );
  OAI22D1BWP30P140 U38 ( .A1(n1), .A2(n14), .B1(n22), .B2(n85), .ZN(N312) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[59]), .ZN(n15) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[27]), .ZN(n86) );
  OAI22D1BWP30P140 U41 ( .A1(n1), .A2(n15), .B1(n22), .B2(n86), .ZN(N314) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[61]), .ZN(n16) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[29]), .ZN(n87) );
  OAI22D1BWP30P140 U44 ( .A1(n1), .A2(n16), .B1(n22), .B2(n87), .ZN(N316) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[63]), .ZN(n17) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[31]), .ZN(n90) );
  OAI22D1BWP30P140 U47 ( .A1(n1), .A2(n17), .B1(n22), .B2(n90), .ZN(N318) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[33]), .ZN(n18) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[1]), .ZN(n58) );
  OAI22D1BWP30P140 U50 ( .A1(n1), .A2(n18), .B1(n22), .B2(n58), .ZN(N288) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[34]), .ZN(n19) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[2]), .ZN(n55) );
  OAI22D1BWP30P140 U53 ( .A1(n1), .A2(n19), .B1(n22), .B2(n55), .ZN(N289) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[35]), .ZN(n20) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[3]), .ZN(n59) );
  OAI22D1BWP30P140 U56 ( .A1(n1), .A2(n20), .B1(n22), .B2(n59), .ZN(N290) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[32]), .ZN(n21) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[0]), .ZN(n54) );
  OAI22D1BWP30P140 U59 ( .A1(n1), .A2(n21), .B1(n22), .B2(n54), .ZN(N287) );
  INVD2BWP30P140 U60 ( .I(i_valid[1]), .ZN(n49) );
  OAI31D1BWP30P140 U61 ( .A1(n48), .A2(n49), .A3(n23), .B(n22), .ZN(N353) );
  INVD1BWP30P140 U62 ( .I(n24), .ZN(n27) );
  INVD1BWP30P140 U63 ( .I(n48), .ZN(n25) );
  OAI21D1BWP30P140 U64 ( .A1(n27), .A2(i_cmd[1]), .B(n26), .ZN(N354) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[7]), .ZN(n62) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[39]), .ZN(n28) );
  OAI22D1BWP30P140 U67 ( .A1(n47), .A2(n62), .B1(n1), .B2(n28), .ZN(N294) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[6]), .ZN(n57) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[38]), .ZN(n29) );
  OAI22D1BWP30P140 U70 ( .A1(n47), .A2(n57), .B1(n1), .B2(n29), .ZN(N293) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[5]), .ZN(n60) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[37]), .ZN(n30) );
  OAI22D1BWP30P140 U73 ( .A1(n47), .A2(n60), .B1(n1), .B2(n30), .ZN(N292) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[4]), .ZN(n56) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[36]), .ZN(n31) );
  OAI22D1BWP30P140 U76 ( .A1(n47), .A2(n56), .B1(n1), .B2(n31), .ZN(N291) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[30]), .ZN(n80) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[62]), .ZN(n32) );
  OAI22D1BWP30P140 U79 ( .A1(n47), .A2(n80), .B1(n1), .B2(n32), .ZN(N317) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[28]), .ZN(n79) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[60]), .ZN(n33) );
  OAI22D1BWP30P140 U82 ( .A1(n47), .A2(n79), .B1(n1), .B2(n33), .ZN(N315) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[26]), .ZN(n78) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[58]), .ZN(n34) );
  OAI22D1BWP30P140 U85 ( .A1(n47), .A2(n78), .B1(n1), .B2(n34), .ZN(N313) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[24]), .ZN(n77) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[56]), .ZN(n35) );
  OAI22D1BWP30P140 U88 ( .A1(n47), .A2(n77), .B1(n1), .B2(n35), .ZN(N311) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[22]), .ZN(n75) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[54]), .ZN(n36) );
  OAI22D1BWP30P140 U91 ( .A1(n47), .A2(n75), .B1(n1), .B2(n36), .ZN(N309) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[18]), .ZN(n70) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[50]), .ZN(n37) );
  OAI22D1BWP30P140 U94 ( .A1(n47), .A2(n70), .B1(n1), .B2(n37), .ZN(N305) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[17]), .ZN(n69) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[49]), .ZN(n38) );
  OAI22D1BWP30P140 U97 ( .A1(n47), .A2(n69), .B1(n1), .B2(n38), .ZN(N304) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[16]), .ZN(n68) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[48]), .ZN(n39) );
  OAI22D1BWP30P140 U100 ( .A1(n47), .A2(n68), .B1(n1), .B2(n39), .ZN(N303) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[15]), .ZN(n67) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[47]), .ZN(n40) );
  OAI22D1BWP30P140 U103 ( .A1(n47), .A2(n67), .B1(n1), .B2(n40), .ZN(N302) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[8]), .ZN(n63) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[40]), .ZN(n41) );
  OAI22D1BWP30P140 U106 ( .A1(n47), .A2(n63), .B1(n1), .B2(n41), .ZN(N295) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[13]), .ZN(n84) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[45]), .ZN(n42) );
  OAI22D1BWP30P140 U109 ( .A1(n47), .A2(n84), .B1(n1), .B2(n42), .ZN(N300) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[12]), .ZN(n65) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[44]), .ZN(n43) );
  OAI22D1BWP30P140 U112 ( .A1(n47), .A2(n65), .B1(n1), .B2(n43), .ZN(N299) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[9]), .ZN(n81) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[41]), .ZN(n44) );
  OAI22D1BWP30P140 U115 ( .A1(n47), .A2(n81), .B1(n1), .B2(n44), .ZN(N296) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[14]), .ZN(n66) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[46]), .ZN(n45) );
  OAI22D1BWP30P140 U118 ( .A1(n47), .A2(n66), .B1(n1), .B2(n45), .ZN(N301) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[11]), .ZN(n82) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[43]), .ZN(n46) );
  OAI22D1BWP30P140 U121 ( .A1(n47), .A2(n82), .B1(n1), .B2(n46), .ZN(N298) );
  MUX2NUD1BWP30P140 U122 ( .I0(n50), .I1(n49), .S(i_cmd[0]), .ZN(n51) );
  ND2OPTIBD1BWP30P140 U123 ( .A1(n52), .A2(n51), .ZN(n53) );
  INVD2BWP30P140 U124 ( .I(n53), .ZN(n72) );
  MOAI22D1BWP30P140 U125 ( .A1(n54), .A2(n89), .B1(i_data_bus[32]), .B2(n88), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U126 ( .A1(n55), .A2(n61), .B1(i_data_bus[34]), .B2(n88), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n61), .B1(i_data_bus[36]), .B2(n88), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n61), .B1(i_data_bus[38]), .B2(n88), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n61), .B1(i_data_bus[33]), .B2(n88), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n61), .B1(i_data_bus[35]), .B2(n88), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n61), .B1(i_data_bus[37]), .B2(n88), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n61), .B1(i_data_bus[39]), .B2(n88), 
        .ZN(N326) );
  INVD2BWP30P140 U133 ( .I(n72), .ZN(n83) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n83), .B1(i_data_bus[40]), .B2(n88), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n83), .B1(i_data_bus[42]), .B2(n88), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n83), .B1(i_data_bus[44]), .B2(n88), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n83), .B1(i_data_bus[46]), .B2(n88), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n83), .B1(i_data_bus[47]), .B2(n88), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n83), .B1(i_data_bus[48]), .B2(n88), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n83), .B1(i_data_bus[49]), .B2(n88), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n83), .B1(i_data_bus[50]), .B2(n88), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n83), .B1(i_data_bus[51]), .B2(n88), 
        .ZN(N338) );
  INVD2BWP30P140 U143 ( .I(n72), .ZN(n89) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n89), .B1(i_data_bus[52]), .B2(n88), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n89), .B1(i_data_bus[53]), .B2(n88), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n89), .B1(i_data_bus[54]), .B2(n88), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n89), .B1(i_data_bus[55]), .B2(n88), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n89), .B1(i_data_bus[56]), .B2(n88), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n89), .B1(i_data_bus[58]), .B2(n88), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n89), .B1(i_data_bus[60]), .B2(n88), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n89), .B1(i_data_bus[62]), .B2(n88), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n83), .B1(i_data_bus[41]), .B2(n88), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n83), .B1(i_data_bus[43]), .B2(n88), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n83), .B1(i_data_bus[45]), .B2(n88), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n89), .B1(i_data_bus[57]), .B2(n88), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n89), .B1(i_data_bus[59]), .B2(n88), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n89), .B1(i_data_bus[61]), .B2(n88), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U158 ( .A1(n90), .A2(n89), .B1(i_data_bus[63]), .B2(n88), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_2 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91;

  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n46), .Z(n89) );
  ND2OPTIBD1BWP30P140 U4 ( .A1(n45), .A2(n44), .ZN(n5) );
  NR2D1BWP30P140 U5 ( .A1(n49), .A2(i_cmd[1]), .ZN(n53) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n49), .ZN(n45) );
  INVD1BWP30P140 U7 ( .I(i_cmd[0]), .ZN(n44) );
  INVD2BWP30P140 U8 ( .I(n4), .ZN(n16) );
  INVD2BWP30P140 U9 ( .I(n28), .ZN(n43) );
  INVD4BWP30P140 U10 ( .I(n28), .ZN(n26) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n3), .A2(n2), .ZN(n4) );
  NR2D1BWP30P140 U12 ( .A1(n49), .A2(n44), .ZN(n2) );
  MUX2NUD1BWP30P140 U13 ( .I0(n51), .I1(n50), .S(i_cmd[1]), .ZN(n3) );
  ND2D1BWP30P140 U14 ( .A1(n1), .A2(i_en), .ZN(n49) );
  INVD1BWP30P140 U15 ( .I(n89), .ZN(n47) );
  INVD1BWP30P140 U16 ( .I(i_valid[0]), .ZN(n51) );
  INVD1BWP30P140 U17 ( .I(rst), .ZN(n1) );
  INVD2BWP30P140 U18 ( .I(n16), .ZN(n38) );
  INVD1BWP30P140 U19 ( .I(i_data_bus[40]), .ZN(n6) );
  INVD2BWP30P140 U20 ( .I(n5), .ZN(n28) );
  INVD1BWP30P140 U21 ( .I(i_data_bus[8]), .ZN(n87) );
  OAI22D1BWP30P140 U22 ( .A1(n38), .A2(n6), .B1(n26), .B2(n87), .ZN(N295) );
  INVD1BWP30P140 U23 ( .I(i_data_bus[42]), .ZN(n7) );
  INVD1BWP30P140 U24 ( .I(i_data_bus[10]), .ZN(n88) );
  OAI22D1BWP30P140 U25 ( .A1(n38), .A2(n7), .B1(n26), .B2(n88), .ZN(N297) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[43]), .ZN(n8) );
  INVD1BWP30P140 U27 ( .I(i_data_bus[11]), .ZN(n78) );
  OAI22D1BWP30P140 U28 ( .A1(n38), .A2(n8), .B1(n26), .B2(n78), .ZN(N298) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[44]), .ZN(n9) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[12]), .ZN(n91) );
  OAI22D1BWP30P140 U31 ( .A1(n38), .A2(n9), .B1(n26), .B2(n91), .ZN(N299) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[45]), .ZN(n10) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[13]), .ZN(n79) );
  OAI22D1BWP30P140 U34 ( .A1(n38), .A2(n10), .B1(n26), .B2(n79), .ZN(N300) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[46]), .ZN(n11) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[14]), .ZN(n86) );
  OAI22D1BWP30P140 U37 ( .A1(n38), .A2(n11), .B1(n26), .B2(n86), .ZN(N301) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[47]), .ZN(n12) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[15]), .ZN(n85) );
  OAI22D1BWP30P140 U40 ( .A1(n38), .A2(n12), .B1(n26), .B2(n85), .ZN(N302) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[48]), .ZN(n13) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[16]), .ZN(n64) );
  OAI22D1BWP30P140 U43 ( .A1(n38), .A2(n13), .B1(n26), .B2(n64), .ZN(N303) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[49]), .ZN(n14) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[17]), .ZN(n65) );
  OAI22D1BWP30P140 U46 ( .A1(n38), .A2(n14), .B1(n26), .B2(n65), .ZN(N304) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[50]), .ZN(n15) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[18]), .ZN(n66) );
  OAI22D1BWP30P140 U49 ( .A1(n38), .A2(n15), .B1(n26), .B2(n66), .ZN(N305) );
  INVD2BWP30P140 U50 ( .I(n16), .ZN(n42) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[54]), .ZN(n17) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[22]), .ZN(n71) );
  OAI22D1BWP30P140 U53 ( .A1(n42), .A2(n17), .B1(n26), .B2(n71), .ZN(N309) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[56]), .ZN(n18) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[24]), .ZN(n73) );
  OAI22D1BWP30P140 U56 ( .A1(n42), .A2(n18), .B1(n26), .B2(n73), .ZN(N311) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[58]), .ZN(n19) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[26]), .ZN(n74) );
  OAI22D1BWP30P140 U59 ( .A1(n42), .A2(n19), .B1(n26), .B2(n74), .ZN(N313) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[60]), .ZN(n20) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[28]), .ZN(n75) );
  OAI22D1BWP30P140 U62 ( .A1(n42), .A2(n20), .B1(n26), .B2(n75), .ZN(N315) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[62]), .ZN(n21) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[30]), .ZN(n76) );
  OAI22D1BWP30P140 U65 ( .A1(n42), .A2(n21), .B1(n26), .B2(n76), .ZN(N317) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[36]), .ZN(n22) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[4]), .ZN(n57) );
  OAI22D1BWP30P140 U68 ( .A1(n38), .A2(n22), .B1(n26), .B2(n57), .ZN(N291) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[37]), .ZN(n23) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[5]), .ZN(n61) );
  OAI22D1BWP30P140 U71 ( .A1(n42), .A2(n23), .B1(n26), .B2(n61), .ZN(N292) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[41]), .ZN(n24) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[9]), .ZN(n77) );
  OAI22D1BWP30P140 U74 ( .A1(n38), .A2(n24), .B1(n26), .B2(n77), .ZN(N296) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[38]), .ZN(n25) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[6]), .ZN(n58) );
  OAI22D1BWP30P140 U77 ( .A1(n38), .A2(n25), .B1(n26), .B2(n58), .ZN(N293) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[39]), .ZN(n27) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[7]), .ZN(n63) );
  OAI22D1BWP30P140 U80 ( .A1(n42), .A2(n27), .B1(n26), .B2(n63), .ZN(N294) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[35]), .ZN(n29) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[3]), .ZN(n60) );
  OAI22D1BWP30P140 U83 ( .A1(n42), .A2(n29), .B1(n43), .B2(n60), .ZN(N290) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[34]), .ZN(n30) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[2]), .ZN(n56) );
  OAI22D1BWP30P140 U86 ( .A1(n38), .A2(n30), .B1(n43), .B2(n56), .ZN(N289) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[33]), .ZN(n31) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[1]), .ZN(n59) );
  OAI22D1BWP30P140 U89 ( .A1(n42), .A2(n31), .B1(n43), .B2(n59), .ZN(N288) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[32]), .ZN(n32) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[0]), .ZN(n55) );
  OAI22D1BWP30P140 U92 ( .A1(n38), .A2(n32), .B1(n43), .B2(n55), .ZN(N287) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[63]), .ZN(n33) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[31]), .ZN(n84) );
  OAI22D1BWP30P140 U95 ( .A1(n42), .A2(n33), .B1(n43), .B2(n84), .ZN(N318) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[61]), .ZN(n34) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[29]), .ZN(n82) );
  OAI22D1BWP30P140 U98 ( .A1(n42), .A2(n34), .B1(n43), .B2(n82), .ZN(N316) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[59]), .ZN(n35) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[27]), .ZN(n81) );
  OAI22D1BWP30P140 U101 ( .A1(n42), .A2(n35), .B1(n43), .B2(n81), .ZN(N314) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[52]), .ZN(n36) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[20]), .ZN(n69) );
  OAI22D1BWP30P140 U104 ( .A1(n42), .A2(n36), .B1(n43), .B2(n69), .ZN(N307) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[51]), .ZN(n37) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[19]), .ZN(n67) );
  OAI22D1BWP30P140 U107 ( .A1(n38), .A2(n37), .B1(n43), .B2(n67), .ZN(N306) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[55]), .ZN(n39) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[23]), .ZN(n72) );
  OAI22D1BWP30P140 U110 ( .A1(n42), .A2(n39), .B1(n43), .B2(n72), .ZN(N310) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[57]), .ZN(n40) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[25]), .ZN(n80) );
  OAI22D1BWP30P140 U113 ( .A1(n42), .A2(n40), .B1(n26), .B2(n80), .ZN(N312) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[53]), .ZN(n41) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[21]), .ZN(n70) );
  OAI22D1BWP30P140 U116 ( .A1(n42), .A2(n41), .B1(n26), .B2(n70), .ZN(N308) );
  INVD2BWP30P140 U117 ( .I(i_valid[1]), .ZN(n50) );
  OAI31D1BWP30P140 U118 ( .A1(n49), .A2(n50), .A3(n44), .B(n26), .ZN(N353) );
  INVD1BWP30P140 U119 ( .I(n45), .ZN(n48) );
  INVD1BWP30P140 U120 ( .I(n49), .ZN(n46) );
  OAI21D1BWP30P140 U121 ( .A1(n48), .A2(i_cmd[1]), .B(n47), .ZN(N354) );
  MUX2NUD1BWP30P140 U122 ( .I0(n51), .I1(n50), .S(i_cmd[0]), .ZN(n52) );
  ND2OPTIBD1BWP30P140 U123 ( .A1(n53), .A2(n52), .ZN(n54) );
  INVD2BWP30P140 U124 ( .I(n54), .ZN(n68) );
  INVD2BWP30P140 U125 ( .I(n68), .ZN(n62) );
  MOAI22D1BWP30P140 U126 ( .A1(n55), .A2(n62), .B1(i_data_bus[32]), .B2(n89), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n62), .B1(i_data_bus[34]), .B2(n89), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n62), .B1(i_data_bus[36]), .B2(n89), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n62), .B1(i_data_bus[38]), .B2(n89), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n62), .B1(i_data_bus[33]), .B2(n89), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n62), .B1(i_data_bus[35]), .B2(n89), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n62), .B1(i_data_bus[37]), .B2(n89), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n62), .B1(i_data_bus[39]), .B2(n89), 
        .ZN(N326) );
  INVD2BWP30P140 U134 ( .I(n68), .ZN(n90) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n90), .B1(i_data_bus[48]), .B2(n89), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n90), .B1(i_data_bus[49]), .B2(n89), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n90), .B1(i_data_bus[50]), .B2(n89), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n90), .B1(i_data_bus[51]), .B2(n89), 
        .ZN(N338) );
  INVD2BWP30P140 U139 ( .I(n68), .ZN(n83) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n83), .B1(i_data_bus[52]), .B2(n89), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n83), .B1(i_data_bus[53]), .B2(n89), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n83), .B1(i_data_bus[54]), .B2(n89), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n83), .B1(i_data_bus[55]), .B2(n89), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n83), .B1(i_data_bus[56]), .B2(n89), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n83), .B1(i_data_bus[58]), .B2(n89), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n83), .B1(i_data_bus[60]), .B2(n89), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n83), .B1(i_data_bus[62]), .B2(n89), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n90), .B1(i_data_bus[41]), .B2(n89), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n90), .B1(i_data_bus[43]), .B2(n89), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n90), .B1(i_data_bus[45]), .B2(n89), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n83), .B1(i_data_bus[57]), .B2(n89), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n83), .B1(i_data_bus[59]), .B2(n89), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n83), .B1(i_data_bus[61]), .B2(n89), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n83), .B1(i_data_bus[63]), .B2(n89), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n90), .B1(i_data_bus[47]), .B2(n89), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n90), .B1(i_data_bus[46]), .B2(n89), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n90), .B1(i_data_bus[40]), .B2(n89), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n90), .B1(i_data_bus[42]), .B2(n89), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n91), .A2(n90), .B1(i_data_bus[44]), .B2(n89), 
        .ZN(N331) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_3 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91;

  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n46), .Z(n89) );
  NR2D1BWP30P140 U4 ( .A1(n49), .A2(i_cmd[1]), .ZN(n53) );
  OAI31D0BWP30P140 U5 ( .A1(n49), .A2(n50), .A3(n44), .B(n26), .ZN(N353) );
  INVD2BWP30P140 U6 ( .I(n4), .ZN(n7) );
  ND2OPTIBD1BWP30P140 U7 ( .A1(n3), .A2(n2), .ZN(n4) );
  NR2D1BWP30P140 U8 ( .A1(n49), .A2(n44), .ZN(n2) );
  MUX2NUD1BWP30P140 U9 ( .I0(n51), .I1(n50), .S(i_cmd[1]), .ZN(n3) );
  INVD2BWP30P140 U10 ( .I(n28), .ZN(n26) );
  INVD1BWP30P140 U11 ( .I(i_cmd[0]), .ZN(n44) );
  ND2D1BWP30P140 U12 ( .A1(n1), .A2(i_en), .ZN(n49) );
  OAI22D1BWP30P140 U13 ( .A1(n40), .A2(n6), .B1(n26), .B2(n64), .ZN(N295) );
  INVD1BWP30P140 U14 ( .I(n89), .ZN(n47) );
  INVD1BWP30P140 U15 ( .I(i_valid[0]), .ZN(n51) );
  INVD1BWP30P140 U16 ( .I(rst), .ZN(n1) );
  INVD2BWP30P140 U17 ( .I(n7), .ZN(n40) );
  INVD1BWP30P140 U18 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D2BWP30P140 U19 ( .A1(i_valid[0]), .B1(n49), .ZN(n45) );
  CKND2D2BWP30P140 U20 ( .A1(n45), .A2(n44), .ZN(n5) );
  INVD2BWP30P140 U21 ( .I(n5), .ZN(n28) );
  INVD1BWP30P140 U22 ( .I(i_data_bus[8]), .ZN(n64) );
  INVD2BWP30P140 U23 ( .I(n7), .ZN(n42) );
  INVD1BWP30P140 U24 ( .I(i_data_bus[39]), .ZN(n8) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[7]), .ZN(n55) );
  OAI22D1BWP30P140 U26 ( .A1(n42), .A2(n8), .B1(n43), .B2(n55), .ZN(N294) );
  INVD1BWP30P140 U27 ( .I(i_data_bus[38]), .ZN(n9) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[6]), .ZN(n58) );
  OAI22D1BWP30P140 U29 ( .A1(n40), .A2(n9), .B1(n26), .B2(n58), .ZN(N293) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[37]), .ZN(n10) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[5]), .ZN(n63) );
  OAI22D1BWP30P140 U32 ( .A1(n42), .A2(n10), .B1(n43), .B2(n63), .ZN(N292) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[36]), .ZN(n11) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[4]), .ZN(n59) );
  OAI22D1BWP30P140 U35 ( .A1(n40), .A2(n11), .B1(n26), .B2(n59), .ZN(N291) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[62]), .ZN(n12) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[30]), .ZN(n81) );
  OAI22D1BWP30P140 U38 ( .A1(n42), .A2(n12), .B1(n43), .B2(n81), .ZN(N317) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[60]), .ZN(n13) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[28]), .ZN(n80) );
  OAI22D1BWP30P140 U41 ( .A1(n42), .A2(n13), .B1(n26), .B2(n80), .ZN(N315) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[58]), .ZN(n14) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[26]), .ZN(n79) );
  OAI22D1BWP30P140 U44 ( .A1(n42), .A2(n14), .B1(n43), .B2(n79), .ZN(N313) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[56]), .ZN(n15) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[24]), .ZN(n78) );
  OAI22D1BWP30P140 U47 ( .A1(n42), .A2(n15), .B1(n26), .B2(n78), .ZN(N311) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[54]), .ZN(n16) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[22]), .ZN(n76) );
  OAI22D1BWP30P140 U50 ( .A1(n42), .A2(n16), .B1(n43), .B2(n76), .ZN(N309) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[50]), .ZN(n17) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[18]), .ZN(n71) );
  OAI22D1BWP30P140 U53 ( .A1(n40), .A2(n17), .B1(n26), .B2(n71), .ZN(N305) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[49]), .ZN(n18) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[17]), .ZN(n70) );
  OAI22D1BWP30P140 U56 ( .A1(n40), .A2(n18), .B1(n43), .B2(n70), .ZN(N304) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[48]), .ZN(n19) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[16]), .ZN(n69) );
  OAI22D1BWP30P140 U59 ( .A1(n40), .A2(n19), .B1(n26), .B2(n69), .ZN(N303) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[47]), .ZN(n20) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n68) );
  OAI22D1BWP30P140 U62 ( .A1(n40), .A2(n20), .B1(n43), .B2(n68), .ZN(N302) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[46]), .ZN(n21) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[14]), .ZN(n67) );
  OAI22D1BWP30P140 U65 ( .A1(n40), .A2(n21), .B1(n26), .B2(n67), .ZN(N301) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[45]), .ZN(n22) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[13]), .ZN(n85) );
  OAI22D1BWP30P140 U68 ( .A1(n40), .A2(n22), .B1(n43), .B2(n85), .ZN(N300) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[44]), .ZN(n23) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[12]), .ZN(n66) );
  OAI22D1BWP30P140 U71 ( .A1(n40), .A2(n23), .B1(n26), .B2(n66), .ZN(N299) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[43]), .ZN(n24) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[11]), .ZN(n83) );
  OAI22D1BWP30P140 U74 ( .A1(n40), .A2(n24), .B1(n43), .B2(n83), .ZN(N298) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[42]), .ZN(n25) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[10]), .ZN(n65) );
  OAI22D1BWP30P140 U77 ( .A1(n40), .A2(n25), .B1(n26), .B2(n65), .ZN(N297) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[41]), .ZN(n27) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[9]), .ZN(n82) );
  OAI22D1BWP30P140 U80 ( .A1(n40), .A2(n27), .B1(n43), .B2(n82), .ZN(N296) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[61]), .ZN(n29) );
  INVD2BWP30P140 U82 ( .I(n28), .ZN(n43) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[29]), .ZN(n88) );
  OAI22D1BWP30P140 U84 ( .A1(n42), .A2(n29), .B1(n26), .B2(n88), .ZN(N316) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[63]), .ZN(n30) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[31]), .ZN(n91) );
  OAI22D1BWP30P140 U87 ( .A1(n42), .A2(n30), .B1(n43), .B2(n91), .ZN(N318) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[35]), .ZN(n31) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[3]), .ZN(n56) );
  OAI22D1BWP30P140 U90 ( .A1(n42), .A2(n31), .B1(n26), .B2(n56), .ZN(N290) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[59]), .ZN(n32) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[27]), .ZN(n87) );
  OAI22D1BWP30P140 U93 ( .A1(n42), .A2(n32), .B1(n43), .B2(n87), .ZN(N314) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[34]), .ZN(n33) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[2]), .ZN(n60) );
  OAI22D1BWP30P140 U96 ( .A1(n40), .A2(n33), .B1(n26), .B2(n60), .ZN(N289) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[55]), .ZN(n34) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[23]), .ZN(n77) );
  OAI22D1BWP30P140 U99 ( .A1(n42), .A2(n34), .B1(n43), .B2(n77), .ZN(N310) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[53]), .ZN(n35) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[21]), .ZN(n75) );
  OAI22D1BWP30P140 U102 ( .A1(n42), .A2(n35), .B1(n26), .B2(n75), .ZN(N308) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[51]), .ZN(n36) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[19]), .ZN(n72) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n36), .B1(n43), .B2(n72), .ZN(N306) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[57]), .ZN(n37) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[25]), .ZN(n86) );
  OAI22D1BWP30P140 U108 ( .A1(n42), .A2(n37), .B1(n26), .B2(n86), .ZN(N312) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[33]), .ZN(n38) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[1]), .ZN(n57) );
  OAI22D1BWP30P140 U111 ( .A1(n42), .A2(n38), .B1(n43), .B2(n57), .ZN(N288) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[32]), .ZN(n39) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[0]), .ZN(n61) );
  OAI22D1BWP30P140 U114 ( .A1(n40), .A2(n39), .B1(n26), .B2(n61), .ZN(N287) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[52]), .ZN(n41) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[20]), .ZN(n74) );
  OAI22D1BWP30P140 U117 ( .A1(n42), .A2(n41), .B1(n43), .B2(n74), .ZN(N307) );
  INVD2BWP30P140 U118 ( .I(i_valid[1]), .ZN(n50) );
  INVD1BWP30P140 U119 ( .I(n45), .ZN(n48) );
  INVD1BWP30P140 U120 ( .I(n49), .ZN(n46) );
  OAI21D1BWP30P140 U121 ( .A1(n48), .A2(i_cmd[1]), .B(n47), .ZN(N354) );
  MUX2NUD1BWP30P140 U122 ( .I0(n51), .I1(n50), .S(i_cmd[0]), .ZN(n52) );
  ND2OPTIBD1BWP30P140 U123 ( .A1(n53), .A2(n52), .ZN(n54) );
  INVD2BWP30P140 U124 ( .I(n54), .ZN(n73) );
  INVD2BWP30P140 U125 ( .I(n73), .ZN(n62) );
  MOAI22D1BWP30P140 U126 ( .A1(n55), .A2(n62), .B1(i_data_bus[39]), .B2(n89), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n62), .B1(i_data_bus[35]), .B2(n89), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n62), .B1(i_data_bus[33]), .B2(n89), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n62), .B1(i_data_bus[38]), .B2(n89), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n62), .B1(i_data_bus[36]), .B2(n89), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n62), .B1(i_data_bus[34]), .B2(n89), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n62), .B1(i_data_bus[32]), .B2(n89), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n62), .B1(i_data_bus[37]), .B2(n89), 
        .ZN(N324) );
  INVD2BWP30P140 U134 ( .I(n73), .ZN(n84) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n84), .B1(i_data_bus[40]), .B2(n89), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n84), .B1(i_data_bus[42]), .B2(n89), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n84), .B1(i_data_bus[44]), .B2(n89), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n84), .B1(i_data_bus[46]), .B2(n89), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n84), .B1(i_data_bus[47]), .B2(n89), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n84), .B1(i_data_bus[48]), .B2(n89), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n84), .B1(i_data_bus[49]), .B2(n89), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n84), .B1(i_data_bus[50]), .B2(n89), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n84), .B1(i_data_bus[51]), .B2(n89), 
        .ZN(N338) );
  INVD2BWP30P140 U144 ( .I(n73), .ZN(n90) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n90), .B1(i_data_bus[52]), .B2(n89), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n90), .B1(i_data_bus[53]), .B2(n89), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n90), .B1(i_data_bus[54]), .B2(n89), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n90), .B1(i_data_bus[55]), .B2(n89), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n90), .B1(i_data_bus[56]), .B2(n89), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n90), .B1(i_data_bus[58]), .B2(n89), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n90), .B1(i_data_bus[60]), .B2(n89), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n90), .B1(i_data_bus[62]), .B2(n89), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n84), .B1(i_data_bus[41]), .B2(n89), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n84), .B1(i_data_bus[43]), .B2(n89), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n84), .B1(i_data_bus[45]), .B2(n89), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n90), .B1(i_data_bus[57]), .B2(n89), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n90), .B1(i_data_bus[59]), .B2(n89), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n90), .B1(i_data_bus[61]), .B2(n89), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n91), .A2(n90), .B1(i_data_bus[63]), .B2(n89), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_4 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91;

  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n46), .Z(n89) );
  NR2D1BWP30P140 U4 ( .A1(n49), .A2(i_cmd[1]), .ZN(n53) );
  OAI31D0BWP30P140 U5 ( .A1(n49), .A2(n50), .A3(n44), .B(n26), .ZN(N353) );
  INVD2BWP30P140 U6 ( .I(n4), .ZN(n7) );
  ND2OPTIBD1BWP30P140 U7 ( .A1(n3), .A2(n2), .ZN(n4) );
  NR2D1BWP30P140 U8 ( .A1(n49), .A2(n44), .ZN(n2) );
  MUX2NUD1BWP30P140 U9 ( .I0(n51), .I1(n50), .S(i_cmd[1]), .ZN(n3) );
  INVD2BWP30P140 U10 ( .I(n28), .ZN(n26) );
  INVD1BWP30P140 U11 ( .I(i_cmd[0]), .ZN(n44) );
  ND2D1BWP30P140 U12 ( .A1(n1), .A2(i_en), .ZN(n49) );
  OAI22D1BWP30P140 U13 ( .A1(n40), .A2(n6), .B1(n26), .B2(n79), .ZN(N313) );
  INVD1BWP30P140 U14 ( .I(n89), .ZN(n47) );
  INVD1BWP30P140 U15 ( .I(i_valid[0]), .ZN(n51) );
  INVD1BWP30P140 U16 ( .I(rst), .ZN(n1) );
  INVD2BWP30P140 U17 ( .I(n7), .ZN(n40) );
  INVD1BWP30P140 U18 ( .I(i_data_bus[58]), .ZN(n6) );
  INR2D2BWP30P140 U19 ( .A1(i_valid[0]), .B1(n49), .ZN(n45) );
  CKND2D2BWP30P140 U20 ( .A1(n45), .A2(n44), .ZN(n5) );
  INVD2BWP30P140 U21 ( .I(n5), .ZN(n28) );
  INVD1BWP30P140 U22 ( .I(i_data_bus[26]), .ZN(n79) );
  INVD2BWP30P140 U23 ( .I(n7), .ZN(n42) );
  INVD1BWP30P140 U24 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[10]), .ZN(n65) );
  OAI22D1BWP30P140 U26 ( .A1(n42), .A2(n8), .B1(n43), .B2(n65), .ZN(N297) );
  INVD1BWP30P140 U27 ( .I(i_data_bus[40]), .ZN(n9) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[8]), .ZN(n64) );
  OAI22D1BWP30P140 U29 ( .A1(n42), .A2(n9), .B1(n26), .B2(n64), .ZN(N295) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[41]), .ZN(n10) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[9]), .ZN(n82) );
  OAI22D1BWP30P140 U32 ( .A1(n42), .A2(n10), .B1(n43), .B2(n82), .ZN(N296) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[39]), .ZN(n11) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[7]), .ZN(n55) );
  OAI22D1BWP30P140 U35 ( .A1(n40), .A2(n11), .B1(n26), .B2(n55), .ZN(N294) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[38]), .ZN(n12) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[6]), .ZN(n59) );
  OAI22D1BWP30P140 U38 ( .A1(n42), .A2(n12), .B1(n43), .B2(n59), .ZN(N293) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[37]), .ZN(n13) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[5]), .ZN(n56) );
  OAI22D1BWP30P140 U41 ( .A1(n40), .A2(n13), .B1(n26), .B2(n56), .ZN(N292) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[54]), .ZN(n14) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[22]), .ZN(n76) );
  OAI22D1BWP30P140 U44 ( .A1(n40), .A2(n14), .B1(n43), .B2(n76), .ZN(N309) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[44]), .ZN(n15) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[12]), .ZN(n66) );
  OAI22D1BWP30P140 U47 ( .A1(n42), .A2(n15), .B1(n26), .B2(n66), .ZN(N299) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[45]), .ZN(n16) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[13]), .ZN(n85) );
  OAI22D1BWP30P140 U50 ( .A1(n42), .A2(n16), .B1(n43), .B2(n85), .ZN(N300) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[46]), .ZN(n17) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[14]), .ZN(n67) );
  OAI22D1BWP30P140 U53 ( .A1(n42), .A2(n17), .B1(n26), .B2(n67), .ZN(N301) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[36]), .ZN(n18) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[4]), .ZN(n60) );
  OAI22D1BWP30P140 U56 ( .A1(n42), .A2(n18), .B1(n43), .B2(n60), .ZN(N291) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[62]), .ZN(n19) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[30]), .ZN(n81) );
  OAI22D1BWP30P140 U59 ( .A1(n40), .A2(n19), .B1(n26), .B2(n81), .ZN(N317) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[49]), .ZN(n20) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[17]), .ZN(n70) );
  OAI22D1BWP30P140 U62 ( .A1(n42), .A2(n20), .B1(n43), .B2(n70), .ZN(N304) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[50]), .ZN(n21) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[18]), .ZN(n71) );
  OAI22D1BWP30P140 U65 ( .A1(n42), .A2(n21), .B1(n26), .B2(n71), .ZN(N305) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[43]), .ZN(n22) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[11]), .ZN(n83) );
  OAI22D1BWP30P140 U68 ( .A1(n42), .A2(n22), .B1(n43), .B2(n83), .ZN(N298) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[47]), .ZN(n23) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[15]), .ZN(n68) );
  OAI22D1BWP30P140 U71 ( .A1(n42), .A2(n23), .B1(n26), .B2(n68), .ZN(N302) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[48]), .ZN(n24) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[16]), .ZN(n69) );
  OAI22D1BWP30P140 U74 ( .A1(n42), .A2(n24), .B1(n43), .B2(n69), .ZN(N303) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[60]), .ZN(n25) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[28]), .ZN(n80) );
  OAI22D1BWP30P140 U77 ( .A1(n40), .A2(n25), .B1(n26), .B2(n80), .ZN(N315) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[56]), .ZN(n27) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[24]), .ZN(n78) );
  OAI22D1BWP30P140 U80 ( .A1(n40), .A2(n27), .B1(n43), .B2(n78), .ZN(N311) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[34]), .ZN(n29) );
  INVD2BWP30P140 U82 ( .I(n28), .ZN(n43) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[2]), .ZN(n61) );
  OAI22D1BWP30P140 U84 ( .A1(n42), .A2(n29), .B1(n26), .B2(n61), .ZN(N289) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[35]), .ZN(n30) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[3]), .ZN(n57) );
  OAI22D1BWP30P140 U87 ( .A1(n40), .A2(n30), .B1(n43), .B2(n57), .ZN(N290) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[33]), .ZN(n31) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[1]), .ZN(n58) );
  OAI22D1BWP30P140 U90 ( .A1(n40), .A2(n31), .B1(n26), .B2(n58), .ZN(N288) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[32]), .ZN(n32) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[0]), .ZN(n63) );
  OAI22D1BWP30P140 U93 ( .A1(n42), .A2(n32), .B1(n43), .B2(n63), .ZN(N287) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[63]), .ZN(n33) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[31]), .ZN(n91) );
  OAI22D1BWP30P140 U96 ( .A1(n40), .A2(n33), .B1(n26), .B2(n91), .ZN(N318) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[61]), .ZN(n34) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[29]), .ZN(n88) );
  OAI22D1BWP30P140 U99 ( .A1(n40), .A2(n34), .B1(n43), .B2(n88), .ZN(N316) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[59]), .ZN(n35) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[27]), .ZN(n87) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n35), .B1(n26), .B2(n87), .ZN(N314) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[57]), .ZN(n36) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[25]), .ZN(n86) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n36), .B1(n43), .B2(n86), .ZN(N312) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[55]), .ZN(n37) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[23]), .ZN(n77) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n37), .B1(n26), .B2(n77), .ZN(N310) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[53]), .ZN(n38) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[21]), .ZN(n75) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n38), .B1(n43), .B2(n75), .ZN(N308) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[52]), .ZN(n39) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[20]), .ZN(n74) );
  OAI22D1BWP30P140 U114 ( .A1(n40), .A2(n39), .B1(n26), .B2(n74), .ZN(N307) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[51]), .ZN(n41) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[19]), .ZN(n72) );
  OAI22D1BWP30P140 U117 ( .A1(n42), .A2(n41), .B1(n43), .B2(n72), .ZN(N306) );
  INVD2BWP30P140 U118 ( .I(i_valid[1]), .ZN(n50) );
  INVD1BWP30P140 U119 ( .I(n45), .ZN(n48) );
  INVD1BWP30P140 U120 ( .I(n49), .ZN(n46) );
  OAI21D1BWP30P140 U121 ( .A1(n48), .A2(i_cmd[1]), .B(n47), .ZN(N354) );
  MUX2NUD1BWP30P140 U122 ( .I0(n51), .I1(n50), .S(i_cmd[0]), .ZN(n52) );
  ND2OPTIBD1BWP30P140 U123 ( .A1(n53), .A2(n52), .ZN(n54) );
  INVD2BWP30P140 U124 ( .I(n54), .ZN(n73) );
  INVD2BWP30P140 U125 ( .I(n73), .ZN(n62) );
  MOAI22D1BWP30P140 U126 ( .A1(n55), .A2(n62), .B1(i_data_bus[39]), .B2(n89), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n62), .B1(i_data_bus[37]), .B2(n89), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n62), .B1(i_data_bus[35]), .B2(n89), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n62), .B1(i_data_bus[33]), .B2(n89), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n62), .B1(i_data_bus[38]), .B2(n89), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n62), .B1(i_data_bus[36]), .B2(n89), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n62), .B1(i_data_bus[34]), .B2(n89), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n62), .B1(i_data_bus[32]), .B2(n89), 
        .ZN(N319) );
  INVD2BWP30P140 U134 ( .I(n73), .ZN(n84) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n84), .B1(i_data_bus[40]), .B2(n89), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n84), .B1(i_data_bus[42]), .B2(n89), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n84), .B1(i_data_bus[44]), .B2(n89), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n84), .B1(i_data_bus[46]), .B2(n89), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n84), .B1(i_data_bus[47]), .B2(n89), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n84), .B1(i_data_bus[48]), .B2(n89), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n84), .B1(i_data_bus[49]), .B2(n89), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n84), .B1(i_data_bus[50]), .B2(n89), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n84), .B1(i_data_bus[51]), .B2(n89), 
        .ZN(N338) );
  INVD2BWP30P140 U144 ( .I(n73), .ZN(n90) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n90), .B1(i_data_bus[52]), .B2(n89), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n90), .B1(i_data_bus[53]), .B2(n89), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n90), .B1(i_data_bus[54]), .B2(n89), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n90), .B1(i_data_bus[55]), .B2(n89), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n90), .B1(i_data_bus[56]), .B2(n89), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n90), .B1(i_data_bus[58]), .B2(n89), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n90), .B1(i_data_bus[60]), .B2(n89), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n90), .B1(i_data_bus[62]), .B2(n89), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n84), .B1(i_data_bus[41]), .B2(n89), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n84), .B1(i_data_bus[43]), .B2(n89), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n84), .B1(i_data_bus[45]), .B2(n89), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n90), .B1(i_data_bus[57]), .B2(n89), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n90), .B1(i_data_bus[59]), .B2(n89), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n90), .B1(i_data_bus[61]), .B2(n89), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n91), .A2(n90), .B1(i_data_bus[63]), .B2(n89), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_5 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91;

  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n46), .Z(n89) );
  NR2D1BWP30P140 U4 ( .A1(n49), .A2(i_cmd[1]), .ZN(n53) );
  OAI31D0BWP30P140 U5 ( .A1(n49), .A2(n50), .A3(n44), .B(n26), .ZN(N353) );
  INVD2BWP30P140 U6 ( .I(n4), .ZN(n7) );
  ND2OPTIBD1BWP30P140 U7 ( .A1(n3), .A2(n2), .ZN(n4) );
  NR2D1BWP30P140 U8 ( .A1(n49), .A2(n44), .ZN(n2) );
  MUX2NUD1BWP30P140 U9 ( .I0(n51), .I1(n50), .S(i_cmd[1]), .ZN(n3) );
  INVD2BWP30P140 U10 ( .I(n28), .ZN(n26) );
  INVD1BWP30P140 U11 ( .I(i_cmd[0]), .ZN(n44) );
  ND2D1BWP30P140 U12 ( .A1(n1), .A2(i_en), .ZN(n49) );
  OAI22D1BWP30P140 U13 ( .A1(n40), .A2(n6), .B1(n26), .B2(n55), .ZN(N294) );
  INVD1BWP30P140 U14 ( .I(n89), .ZN(n47) );
  INVD1BWP30P140 U15 ( .I(i_valid[0]), .ZN(n51) );
  INVD1BWP30P140 U16 ( .I(rst), .ZN(n1) );
  INVD2BWP30P140 U17 ( .I(n7), .ZN(n40) );
  INVD1BWP30P140 U18 ( .I(i_data_bus[39]), .ZN(n6) );
  INR2D2BWP30P140 U19 ( .A1(i_valid[0]), .B1(n49), .ZN(n45) );
  CKND2D2BWP30P140 U20 ( .A1(n45), .A2(n44), .ZN(n5) );
  INVD2BWP30P140 U21 ( .I(n5), .ZN(n28) );
  INVD1BWP30P140 U22 ( .I(i_data_bus[7]), .ZN(n55) );
  INVD2BWP30P140 U23 ( .I(n7), .ZN(n42) );
  INVD1BWP30P140 U24 ( .I(i_data_bus[40]), .ZN(n8) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[8]), .ZN(n64) );
  OAI22D1BWP30P140 U26 ( .A1(n42), .A2(n8), .B1(n43), .B2(n64), .ZN(N295) );
  INVD1BWP30P140 U27 ( .I(i_data_bus[41]), .ZN(n9) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[9]), .ZN(n82) );
  OAI22D1BWP30P140 U29 ( .A1(n42), .A2(n9), .B1(n26), .B2(n82), .ZN(N296) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[42]), .ZN(n10) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[10]), .ZN(n65) );
  OAI22D1BWP30P140 U32 ( .A1(n42), .A2(n10), .B1(n43), .B2(n65), .ZN(N297) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[43]), .ZN(n11) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[11]), .ZN(n83) );
  OAI22D1BWP30P140 U35 ( .A1(n42), .A2(n11), .B1(n26), .B2(n83), .ZN(N298) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[44]), .ZN(n12) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[12]), .ZN(n66) );
  OAI22D1BWP30P140 U38 ( .A1(n42), .A2(n12), .B1(n43), .B2(n66), .ZN(N299) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[45]), .ZN(n13) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[13]), .ZN(n85) );
  OAI22D1BWP30P140 U41 ( .A1(n42), .A2(n13), .B1(n26), .B2(n85), .ZN(N300) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[46]), .ZN(n14) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[14]), .ZN(n67) );
  OAI22D1BWP30P140 U44 ( .A1(n42), .A2(n14), .B1(n43), .B2(n67), .ZN(N301) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[47]), .ZN(n15) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[15]), .ZN(n68) );
  OAI22D1BWP30P140 U47 ( .A1(n42), .A2(n15), .B1(n26), .B2(n68), .ZN(N302) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[48]), .ZN(n16) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[16]), .ZN(n69) );
  OAI22D1BWP30P140 U50 ( .A1(n42), .A2(n16), .B1(n43), .B2(n69), .ZN(N303) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[49]), .ZN(n17) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[17]), .ZN(n70) );
  OAI22D1BWP30P140 U53 ( .A1(n42), .A2(n17), .B1(n26), .B2(n70), .ZN(N304) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[50]), .ZN(n18) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[18]), .ZN(n71) );
  OAI22D1BWP30P140 U56 ( .A1(n42), .A2(n18), .B1(n43), .B2(n71), .ZN(N305) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[54]), .ZN(n19) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[22]), .ZN(n76) );
  OAI22D1BWP30P140 U59 ( .A1(n40), .A2(n19), .B1(n26), .B2(n76), .ZN(N309) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[56]), .ZN(n20) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[24]), .ZN(n78) );
  OAI22D1BWP30P140 U62 ( .A1(n40), .A2(n20), .B1(n43), .B2(n78), .ZN(N311) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[58]), .ZN(n21) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[26]), .ZN(n79) );
  OAI22D1BWP30P140 U65 ( .A1(n40), .A2(n21), .B1(n26), .B2(n79), .ZN(N313) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[60]), .ZN(n22) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[28]), .ZN(n80) );
  OAI22D1BWP30P140 U68 ( .A1(n40), .A2(n22), .B1(n43), .B2(n80), .ZN(N315) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[62]), .ZN(n23) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[30]), .ZN(n81) );
  OAI22D1BWP30P140 U71 ( .A1(n40), .A2(n23), .B1(n26), .B2(n81), .ZN(N317) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[36]), .ZN(n24) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[4]), .ZN(n60) );
  OAI22D1BWP30P140 U74 ( .A1(n42), .A2(n24), .B1(n43), .B2(n60), .ZN(N291) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[37]), .ZN(n25) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[5]), .ZN(n56) );
  OAI22D1BWP30P140 U77 ( .A1(n40), .A2(n25), .B1(n26), .B2(n56), .ZN(N292) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[38]), .ZN(n27) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[6]), .ZN(n59) );
  OAI22D1BWP30P140 U80 ( .A1(n42), .A2(n27), .B1(n43), .B2(n59), .ZN(N293) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[35]), .ZN(n29) );
  INVD2BWP30P140 U82 ( .I(n28), .ZN(n43) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[3]), .ZN(n57) );
  OAI22D1BWP30P140 U84 ( .A1(n40), .A2(n29), .B1(n26), .B2(n57), .ZN(N290) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[34]), .ZN(n30) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[2]), .ZN(n61) );
  OAI22D1BWP30P140 U87 ( .A1(n42), .A2(n30), .B1(n43), .B2(n61), .ZN(N289) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[33]), .ZN(n31) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[1]), .ZN(n58) );
  OAI22D1BWP30P140 U90 ( .A1(n40), .A2(n31), .B1(n26), .B2(n58), .ZN(N288) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[32]), .ZN(n32) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[0]), .ZN(n63) );
  OAI22D1BWP30P140 U93 ( .A1(n42), .A2(n32), .B1(n43), .B2(n63), .ZN(N287) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[63]), .ZN(n33) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[31]), .ZN(n88) );
  OAI22D1BWP30P140 U96 ( .A1(n40), .A2(n33), .B1(n26), .B2(n88), .ZN(N318) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[61]), .ZN(n34) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[29]), .ZN(n91) );
  OAI22D1BWP30P140 U99 ( .A1(n40), .A2(n34), .B1(n43), .B2(n91), .ZN(N316) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[59]), .ZN(n35) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[27]), .ZN(n87) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n35), .B1(n26), .B2(n87), .ZN(N314) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[57]), .ZN(n36) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[25]), .ZN(n86) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n36), .B1(n43), .B2(n86), .ZN(N312) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[55]), .ZN(n37) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[23]), .ZN(n77) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n37), .B1(n26), .B2(n77), .ZN(N310) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[53]), .ZN(n38) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[21]), .ZN(n75) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n38), .B1(n43), .B2(n75), .ZN(N308) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[52]), .ZN(n39) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[20]), .ZN(n74) );
  OAI22D1BWP30P140 U114 ( .A1(n40), .A2(n39), .B1(n26), .B2(n74), .ZN(N307) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[51]), .ZN(n41) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[19]), .ZN(n72) );
  OAI22D1BWP30P140 U117 ( .A1(n42), .A2(n41), .B1(n43), .B2(n72), .ZN(N306) );
  INVD2BWP30P140 U118 ( .I(i_valid[1]), .ZN(n50) );
  INVD1BWP30P140 U119 ( .I(n45), .ZN(n48) );
  INVD1BWP30P140 U120 ( .I(n49), .ZN(n46) );
  OAI21D1BWP30P140 U121 ( .A1(n48), .A2(i_cmd[1]), .B(n47), .ZN(N354) );
  MUX2NUD1BWP30P140 U122 ( .I0(n51), .I1(n50), .S(i_cmd[0]), .ZN(n52) );
  ND2OPTIBD1BWP30P140 U123 ( .A1(n53), .A2(n52), .ZN(n54) );
  INVD2BWP30P140 U124 ( .I(n54), .ZN(n73) );
  INVD2BWP30P140 U125 ( .I(n73), .ZN(n62) );
  MOAI22D1BWP30P140 U126 ( .A1(n55), .A2(n62), .B1(i_data_bus[39]), .B2(n89), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n62), .B1(i_data_bus[37]), .B2(n89), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n62), .B1(i_data_bus[35]), .B2(n89), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n62), .B1(i_data_bus[33]), .B2(n89), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n62), .B1(i_data_bus[38]), .B2(n89), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n62), .B1(i_data_bus[36]), .B2(n89), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n62), .B1(i_data_bus[34]), .B2(n89), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n62), .B1(i_data_bus[32]), .B2(n89), 
        .ZN(N319) );
  INVD2BWP30P140 U134 ( .I(n73), .ZN(n84) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n84), .B1(i_data_bus[40]), .B2(n89), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n84), .B1(i_data_bus[42]), .B2(n89), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n84), .B1(i_data_bus[44]), .B2(n89), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n84), .B1(i_data_bus[46]), .B2(n89), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n84), .B1(i_data_bus[47]), .B2(n89), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n84), .B1(i_data_bus[48]), .B2(n89), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n84), .B1(i_data_bus[49]), .B2(n89), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n84), .B1(i_data_bus[50]), .B2(n89), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n84), .B1(i_data_bus[51]), .B2(n89), 
        .ZN(N338) );
  INVD2BWP30P140 U144 ( .I(n73), .ZN(n90) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n90), .B1(i_data_bus[52]), .B2(n89), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n90), .B1(i_data_bus[53]), .B2(n89), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n90), .B1(i_data_bus[54]), .B2(n89), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n90), .B1(i_data_bus[55]), .B2(n89), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n90), .B1(i_data_bus[56]), .B2(n89), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n90), .B1(i_data_bus[58]), .B2(n89), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n90), .B1(i_data_bus[60]), .B2(n89), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n90), .B1(i_data_bus[62]), .B2(n89), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n84), .B1(i_data_bus[41]), .B2(n89), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n84), .B1(i_data_bus[43]), .B2(n89), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n84), .B1(i_data_bus[45]), .B2(n89), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n90), .B1(i_data_bus[57]), .B2(n89), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n90), .B1(i_data_bus[59]), .B2(n89), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n90), .B1(i_data_bus[63]), .B2(n89), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U159 ( .A1(n91), .A2(n90), .B1(i_data_bus[61]), .B2(n89), 
        .ZN(N348) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_6 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91;

  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n46), .Z(n89) );
  NR2D1BWP30P140 U4 ( .A1(n49), .A2(i_cmd[1]), .ZN(n53) );
  OAI31D0BWP30P140 U5 ( .A1(n49), .A2(n50), .A3(n44), .B(n26), .ZN(N353) );
  INVD2BWP30P140 U6 ( .I(n4), .ZN(n15) );
  ND2OPTIBD1BWP30P140 U7 ( .A1(n3), .A2(n2), .ZN(n4) );
  NR2D1BWP30P140 U8 ( .A1(n49), .A2(n44), .ZN(n2) );
  MUX2NUD1BWP30P140 U9 ( .I0(n51), .I1(n50), .S(i_cmd[1]), .ZN(n3) );
  INVD2BWP30P140 U10 ( .I(n28), .ZN(n26) );
  INVD1BWP30P140 U11 ( .I(i_cmd[0]), .ZN(n44) );
  ND2D1BWP30P140 U12 ( .A1(n1), .A2(i_en), .ZN(n49) );
  OAI22D1BWP30P140 U13 ( .A1(n34), .A2(n6), .B1(n26), .B2(n69), .ZN(N303) );
  INVD1BWP30P140 U14 ( .I(n89), .ZN(n47) );
  INVD1BWP30P140 U15 ( .I(i_valid[0]), .ZN(n51) );
  INVD1BWP30P140 U16 ( .I(rst), .ZN(n1) );
  INVD2BWP30P140 U17 ( .I(n15), .ZN(n34) );
  INVD1BWP30P140 U18 ( .I(i_data_bus[48]), .ZN(n6) );
  INR2D2BWP30P140 U19 ( .A1(i_valid[0]), .B1(n49), .ZN(n45) );
  CKND2D2BWP30P140 U20 ( .A1(n45), .A2(n44), .ZN(n5) );
  INVD2BWP30P140 U21 ( .I(n5), .ZN(n28) );
  INVD1BWP30P140 U22 ( .I(i_data_bus[16]), .ZN(n69) );
  INVD1BWP30P140 U23 ( .I(i_data_bus[40]), .ZN(n7) );
  INVD1BWP30P140 U24 ( .I(i_data_bus[8]), .ZN(n64) );
  OAI22D1BWP30P140 U25 ( .A1(n34), .A2(n7), .B1(n43), .B2(n64), .ZN(N295) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[41]), .ZN(n8) );
  INVD1BWP30P140 U27 ( .I(i_data_bus[9]), .ZN(n82) );
  OAI22D1BWP30P140 U28 ( .A1(n34), .A2(n8), .B1(n26), .B2(n82), .ZN(N296) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[11]), .ZN(n83) );
  OAI22D1BWP30P140 U31 ( .A1(n34), .A2(n9), .B1(n43), .B2(n83), .ZN(N298) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[45]), .ZN(n10) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[13]), .ZN(n85) );
  OAI22D1BWP30P140 U34 ( .A1(n34), .A2(n10), .B1(n26), .B2(n85), .ZN(N300) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[46]), .ZN(n11) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[14]), .ZN(n67) );
  OAI22D1BWP30P140 U37 ( .A1(n34), .A2(n11), .B1(n43), .B2(n67), .ZN(N301) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[47]), .ZN(n12) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[15]), .ZN(n68) );
  OAI22D1BWP30P140 U40 ( .A1(n34), .A2(n12), .B1(n26), .B2(n68), .ZN(N302) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[49]), .ZN(n13) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[17]), .ZN(n70) );
  OAI22D1BWP30P140 U43 ( .A1(n34), .A2(n13), .B1(n43), .B2(n70), .ZN(N304) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[50]), .ZN(n14) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[18]), .ZN(n71) );
  OAI22D1BWP30P140 U46 ( .A1(n34), .A2(n14), .B1(n26), .B2(n71), .ZN(N305) );
  INVD2BWP30P140 U47 ( .I(n15), .ZN(n42) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[54]), .ZN(n16) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[22]), .ZN(n76) );
  OAI22D1BWP30P140 U50 ( .A1(n42), .A2(n16), .B1(n43), .B2(n76), .ZN(N309) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[56]), .ZN(n17) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[24]), .ZN(n78) );
  OAI22D1BWP30P140 U53 ( .A1(n42), .A2(n17), .B1(n26), .B2(n78), .ZN(N311) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[58]), .ZN(n18) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[26]), .ZN(n79) );
  OAI22D1BWP30P140 U56 ( .A1(n42), .A2(n18), .B1(n43), .B2(n79), .ZN(N313) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[60]), .ZN(n19) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[28]), .ZN(n80) );
  OAI22D1BWP30P140 U59 ( .A1(n42), .A2(n19), .B1(n26), .B2(n80), .ZN(N315) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[62]), .ZN(n20) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[30]), .ZN(n81) );
  OAI22D1BWP30P140 U62 ( .A1(n42), .A2(n20), .B1(n43), .B2(n81), .ZN(N317) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[42]), .ZN(n21) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[10]), .ZN(n65) );
  OAI22D1BWP30P140 U65 ( .A1(n34), .A2(n21), .B1(n26), .B2(n65), .ZN(N297) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[36]), .ZN(n22) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[4]), .ZN(n60) );
  OAI22D1BWP30P140 U68 ( .A1(n34), .A2(n22), .B1(n43), .B2(n60), .ZN(N291) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[44]), .ZN(n23) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[12]), .ZN(n66) );
  OAI22D1BWP30P140 U71 ( .A1(n34), .A2(n23), .B1(n26), .B2(n66), .ZN(N299) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[37]), .ZN(n24) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[5]), .ZN(n56) );
  OAI22D1BWP30P140 U74 ( .A1(n42), .A2(n24), .B1(n43), .B2(n56), .ZN(N292) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[38]), .ZN(n25) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[6]), .ZN(n59) );
  OAI22D1BWP30P140 U77 ( .A1(n34), .A2(n25), .B1(n26), .B2(n59), .ZN(N293) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[39]), .ZN(n27) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[7]), .ZN(n55) );
  OAI22D1BWP30P140 U80 ( .A1(n42), .A2(n27), .B1(n43), .B2(n55), .ZN(N294) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[51]), .ZN(n29) );
  INVD2BWP30P140 U82 ( .I(n28), .ZN(n43) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[19]), .ZN(n72) );
  OAI22D1BWP30P140 U84 ( .A1(n34), .A2(n29), .B1(n26), .B2(n72), .ZN(N306) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[35]), .ZN(n30) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[3]), .ZN(n57) );
  OAI22D1BWP30P140 U87 ( .A1(n42), .A2(n30), .B1(n43), .B2(n57), .ZN(N290) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[34]), .ZN(n31) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[2]), .ZN(n61) );
  OAI22D1BWP30P140 U90 ( .A1(n34), .A2(n31), .B1(n26), .B2(n61), .ZN(N289) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[33]), .ZN(n32) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[1]), .ZN(n58) );
  OAI22D1BWP30P140 U93 ( .A1(n42), .A2(n32), .B1(n43), .B2(n58), .ZN(N288) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[32]), .ZN(n33) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[0]), .ZN(n63) );
  OAI22D1BWP30P140 U96 ( .A1(n34), .A2(n33), .B1(n26), .B2(n63), .ZN(N287) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[61]), .ZN(n35) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[29]), .ZN(n88) );
  OAI22D1BWP30P140 U99 ( .A1(n42), .A2(n35), .B1(n43), .B2(n88), .ZN(N316) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[59]), .ZN(n36) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[27]), .ZN(n87) );
  OAI22D1BWP30P140 U102 ( .A1(n42), .A2(n36), .B1(n26), .B2(n87), .ZN(N314) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[57]), .ZN(n37) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[25]), .ZN(n86) );
  OAI22D1BWP30P140 U105 ( .A1(n42), .A2(n37), .B1(n43), .B2(n86), .ZN(N312) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[55]), .ZN(n38) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[23]), .ZN(n77) );
  OAI22D1BWP30P140 U108 ( .A1(n42), .A2(n38), .B1(n26), .B2(n77), .ZN(N310) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[53]), .ZN(n39) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[21]), .ZN(n75) );
  OAI22D1BWP30P140 U111 ( .A1(n42), .A2(n39), .B1(n43), .B2(n75), .ZN(N308) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[52]), .ZN(n40) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[20]), .ZN(n74) );
  OAI22D1BWP30P140 U114 ( .A1(n42), .A2(n40), .B1(n26), .B2(n74), .ZN(N307) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[63]), .ZN(n41) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[31]), .ZN(n91) );
  OAI22D1BWP30P140 U117 ( .A1(n42), .A2(n41), .B1(n43), .B2(n91), .ZN(N318) );
  INVD2BWP30P140 U118 ( .I(i_valid[1]), .ZN(n50) );
  INVD1BWP30P140 U119 ( .I(n45), .ZN(n48) );
  INVD1BWP30P140 U120 ( .I(n49), .ZN(n46) );
  OAI21D1BWP30P140 U121 ( .A1(n48), .A2(i_cmd[1]), .B(n47), .ZN(N354) );
  MUX2NUD1BWP30P140 U122 ( .I0(n51), .I1(n50), .S(i_cmd[0]), .ZN(n52) );
  ND2OPTIBD1BWP30P140 U123 ( .A1(n53), .A2(n52), .ZN(n54) );
  INVD2BWP30P140 U124 ( .I(n54), .ZN(n73) );
  INVD2BWP30P140 U125 ( .I(n73), .ZN(n62) );
  MOAI22D1BWP30P140 U126 ( .A1(n55), .A2(n62), .B1(i_data_bus[39]), .B2(n89), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n62), .B1(i_data_bus[37]), .B2(n89), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n62), .B1(i_data_bus[35]), .B2(n89), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n62), .B1(i_data_bus[33]), .B2(n89), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n62), .B1(i_data_bus[38]), .B2(n89), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n62), .B1(i_data_bus[36]), .B2(n89), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n62), .B1(i_data_bus[34]), .B2(n89), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n62), .B1(i_data_bus[32]), .B2(n89), 
        .ZN(N319) );
  INVD2BWP30P140 U134 ( .I(n73), .ZN(n84) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n84), .B1(i_data_bus[40]), .B2(n89), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n84), .B1(i_data_bus[42]), .B2(n89), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n84), .B1(i_data_bus[44]), .B2(n89), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n84), .B1(i_data_bus[46]), .B2(n89), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n84), .B1(i_data_bus[47]), .B2(n89), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n84), .B1(i_data_bus[48]), .B2(n89), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n84), .B1(i_data_bus[49]), .B2(n89), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n84), .B1(i_data_bus[50]), .B2(n89), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n84), .B1(i_data_bus[51]), .B2(n89), 
        .ZN(N338) );
  INVD2BWP30P140 U144 ( .I(n73), .ZN(n90) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n90), .B1(i_data_bus[52]), .B2(n89), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n90), .B1(i_data_bus[53]), .B2(n89), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n90), .B1(i_data_bus[54]), .B2(n89), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n90), .B1(i_data_bus[55]), .B2(n89), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n90), .B1(i_data_bus[56]), .B2(n89), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n90), .B1(i_data_bus[58]), .B2(n89), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n90), .B1(i_data_bus[60]), .B2(n89), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n90), .B1(i_data_bus[62]), .B2(n89), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n84), .B1(i_data_bus[41]), .B2(n89), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n84), .B1(i_data_bus[43]), .B2(n89), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n84), .B1(i_data_bus[45]), .B2(n89), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n90), .B1(i_data_bus[57]), .B2(n89), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n90), .B1(i_data_bus[59]), .B2(n89), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n90), .B1(i_data_bus[61]), .B2(n89), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n91), .A2(n90), .B1(i_data_bus[63]), .B2(n89), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_7 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91;

  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n46), .Z(n89) );
  NR2D1BWP30P140 U4 ( .A1(n49), .A2(i_cmd[1]), .ZN(n53) );
  OAI31D0BWP30P140 U5 ( .A1(n49), .A2(n50), .A3(n44), .B(n26), .ZN(N353) );
  INVD2BWP30P140 U6 ( .I(n4), .ZN(n7) );
  ND2OPTIBD1BWP30P140 U7 ( .A1(n3), .A2(n2), .ZN(n4) );
  NR2D1BWP30P140 U8 ( .A1(n49), .A2(n44), .ZN(n2) );
  MUX2NUD1BWP30P140 U9 ( .I0(n51), .I1(n50), .S(i_cmd[1]), .ZN(n3) );
  INVD2BWP30P140 U10 ( .I(n28), .ZN(n26) );
  INVD1BWP30P140 U11 ( .I(i_cmd[0]), .ZN(n44) );
  ND2D1BWP30P140 U12 ( .A1(n1), .A2(i_en), .ZN(n49) );
  OAI22D1BWP30P140 U13 ( .A1(n40), .A2(n6), .B1(n26), .B2(n78), .ZN(N300) );
  INVD1BWP30P140 U14 ( .I(n89), .ZN(n47) );
  INVD1BWP30P140 U15 ( .I(i_valid[0]), .ZN(n51) );
  INVD1BWP30P140 U16 ( .I(rst), .ZN(n1) );
  INVD2BWP30P140 U17 ( .I(n7), .ZN(n40) );
  INVD1BWP30P140 U18 ( .I(i_data_bus[45]), .ZN(n6) );
  INR2D2BWP30P140 U19 ( .A1(i_valid[0]), .B1(n49), .ZN(n45) );
  CKND2D2BWP30P140 U20 ( .A1(n45), .A2(n44), .ZN(n5) );
  INVD2BWP30P140 U21 ( .I(n5), .ZN(n28) );
  INVD1BWP30P140 U22 ( .I(i_data_bus[13]), .ZN(n78) );
  INVD2BWP30P140 U23 ( .I(n7), .ZN(n42) );
  INVD1BWP30P140 U24 ( .I(i_data_bus[37]), .ZN(n8) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[5]), .ZN(n56) );
  OAI22D1BWP30P140 U26 ( .A1(n42), .A2(n8), .B1(n43), .B2(n56), .ZN(N292) );
  INVD1BWP30P140 U27 ( .I(i_data_bus[58]), .ZN(n9) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[26]), .ZN(n73) );
  OAI22D1BWP30P140 U29 ( .A1(n42), .A2(n9), .B1(n26), .B2(n73), .ZN(N313) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[62]), .ZN(n10) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[30]), .ZN(n75) );
  OAI22D1BWP30P140 U32 ( .A1(n42), .A2(n10), .B1(n43), .B2(n75), .ZN(N317) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[36]), .ZN(n11) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[4]), .ZN(n60) );
  OAI22D1BWP30P140 U35 ( .A1(n40), .A2(n11), .B1(n26), .B2(n60), .ZN(N291) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[38]), .ZN(n12) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[6]), .ZN(n59) );
  OAI22D1BWP30P140 U38 ( .A1(n40), .A2(n12), .B1(n43), .B2(n59), .ZN(N293) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[39]), .ZN(n13) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[7]), .ZN(n55) );
  OAI22D1BWP30P140 U41 ( .A1(n42), .A2(n13), .B1(n26), .B2(n55), .ZN(N294) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[60]), .ZN(n14) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[28]), .ZN(n74) );
  OAI22D1BWP30P140 U44 ( .A1(n42), .A2(n14), .B1(n43), .B2(n74), .ZN(N315) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[54]), .ZN(n15) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[22]), .ZN(n70) );
  OAI22D1BWP30P140 U47 ( .A1(n42), .A2(n15), .B1(n26), .B2(n70), .ZN(N309) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[56]), .ZN(n16) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[24]), .ZN(n72) );
  OAI22D1BWP30P140 U50 ( .A1(n42), .A2(n16), .B1(n43), .B2(n72), .ZN(N311) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[40]), .ZN(n17) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[8]), .ZN(n86) );
  OAI22D1BWP30P140 U53 ( .A1(n40), .A2(n17), .B1(n26), .B2(n86), .ZN(N295) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[41]), .ZN(n18) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[9]), .ZN(n76) );
  OAI22D1BWP30P140 U56 ( .A1(n40), .A2(n18), .B1(n43), .B2(n76), .ZN(N296) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[42]), .ZN(n19) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[10]), .ZN(n87) );
  OAI22D1BWP30P140 U59 ( .A1(n40), .A2(n19), .B1(n26), .B2(n87), .ZN(N297) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[43]), .ZN(n20) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[11]), .ZN(n77) );
  OAI22D1BWP30P140 U62 ( .A1(n40), .A2(n20), .B1(n43), .B2(n77), .ZN(N298) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[44]), .ZN(n21) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[12]), .ZN(n88) );
  OAI22D1BWP30P140 U65 ( .A1(n40), .A2(n21), .B1(n26), .B2(n88), .ZN(N299) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[50]), .ZN(n22) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[18]), .ZN(n65) );
  OAI22D1BWP30P140 U68 ( .A1(n40), .A2(n22), .B1(n43), .B2(n65), .ZN(N305) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[49]), .ZN(n23) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[17]), .ZN(n64) );
  OAI22D1BWP30P140 U71 ( .A1(n40), .A2(n23), .B1(n26), .B2(n64), .ZN(N304) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[48]), .ZN(n24) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[16]), .ZN(n84) );
  OAI22D1BWP30P140 U74 ( .A1(n40), .A2(n24), .B1(n43), .B2(n84), .ZN(N303) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[47]), .ZN(n25) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[15]), .ZN(n85) );
  OAI22D1BWP30P140 U77 ( .A1(n40), .A2(n25), .B1(n26), .B2(n85), .ZN(N302) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[46]), .ZN(n27) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[14]), .ZN(n91) );
  OAI22D1BWP30P140 U80 ( .A1(n40), .A2(n27), .B1(n43), .B2(n91), .ZN(N301) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[51]), .ZN(n29) );
  INVD2BWP30P140 U82 ( .I(n28), .ZN(n43) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[19]), .ZN(n66) );
  OAI22D1BWP30P140 U84 ( .A1(n40), .A2(n29), .B1(n26), .B2(n66), .ZN(N306) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[52]), .ZN(n30) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[20]), .ZN(n68) );
  OAI22D1BWP30P140 U87 ( .A1(n42), .A2(n30), .B1(n43), .B2(n68), .ZN(N307) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[53]), .ZN(n31) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[21]), .ZN(n69) );
  OAI22D1BWP30P140 U90 ( .A1(n42), .A2(n31), .B1(n26), .B2(n69), .ZN(N308) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[55]), .ZN(n32) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[23]), .ZN(n71) );
  OAI22D1BWP30P140 U93 ( .A1(n42), .A2(n32), .B1(n43), .B2(n71), .ZN(N310) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[57]), .ZN(n33) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[25]), .ZN(n79) );
  OAI22D1BWP30P140 U96 ( .A1(n42), .A2(n33), .B1(n26), .B2(n79), .ZN(N312) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[59]), .ZN(n34) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[27]), .ZN(n80) );
  OAI22D1BWP30P140 U99 ( .A1(n42), .A2(n34), .B1(n43), .B2(n80), .ZN(N314) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[61]), .ZN(n35) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[29]), .ZN(n81) );
  OAI22D1BWP30P140 U102 ( .A1(n42), .A2(n35), .B1(n26), .B2(n81), .ZN(N316) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[63]), .ZN(n36) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[31]), .ZN(n83) );
  OAI22D1BWP30P140 U105 ( .A1(n42), .A2(n36), .B1(n43), .B2(n83), .ZN(N318) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[32]), .ZN(n37) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[0]), .ZN(n63) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n37), .B1(n26), .B2(n63), .ZN(N287) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[33]), .ZN(n38) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[1]), .ZN(n58) );
  OAI22D1BWP30P140 U111 ( .A1(n42), .A2(n38), .B1(n43), .B2(n58), .ZN(N288) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[34]), .ZN(n39) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[2]), .ZN(n61) );
  OAI22D1BWP30P140 U114 ( .A1(n40), .A2(n39), .B1(n26), .B2(n61), .ZN(N289) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[35]), .ZN(n41) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[3]), .ZN(n57) );
  OAI22D1BWP30P140 U117 ( .A1(n42), .A2(n41), .B1(n43), .B2(n57), .ZN(N290) );
  INVD2BWP30P140 U118 ( .I(i_valid[1]), .ZN(n50) );
  INVD1BWP30P140 U119 ( .I(n45), .ZN(n48) );
  INVD1BWP30P140 U120 ( .I(n49), .ZN(n46) );
  OAI21D1BWP30P140 U121 ( .A1(n48), .A2(i_cmd[1]), .B(n47), .ZN(N354) );
  MUX2NUD1BWP30P140 U122 ( .I0(n51), .I1(n50), .S(i_cmd[0]), .ZN(n52) );
  ND2OPTIBD1BWP30P140 U123 ( .A1(n53), .A2(n52), .ZN(n54) );
  INVD2BWP30P140 U124 ( .I(n54), .ZN(n67) );
  INVD2BWP30P140 U125 ( .I(n67), .ZN(n62) );
  MOAI22D1BWP30P140 U126 ( .A1(n55), .A2(n62), .B1(i_data_bus[39]), .B2(n89), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n62), .B1(i_data_bus[37]), .B2(n89), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n62), .B1(i_data_bus[35]), .B2(n89), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n62), .B1(i_data_bus[33]), .B2(n89), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n62), .B1(i_data_bus[38]), .B2(n89), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n62), .B1(i_data_bus[36]), .B2(n89), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n62), .B1(i_data_bus[34]), .B2(n89), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n62), .B1(i_data_bus[32]), .B2(n89), 
        .ZN(N319) );
  INVD2BWP30P140 U134 ( .I(n67), .ZN(n90) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n90), .B1(i_data_bus[49]), .B2(n89), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n90), .B1(i_data_bus[50]), .B2(n89), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n90), .B1(i_data_bus[51]), .B2(n89), 
        .ZN(N338) );
  INVD2BWP30P140 U138 ( .I(n67), .ZN(n82) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n82), .B1(i_data_bus[52]), .B2(n89), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n82), .B1(i_data_bus[53]), .B2(n89), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n82), .B1(i_data_bus[54]), .B2(n89), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n82), .B1(i_data_bus[55]), .B2(n89), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n82), .B1(i_data_bus[56]), .B2(n89), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n82), .B1(i_data_bus[58]), .B2(n89), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n82), .B1(i_data_bus[60]), .B2(n89), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n82), .B1(i_data_bus[62]), .B2(n89), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n90), .B1(i_data_bus[41]), .B2(n89), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n90), .B1(i_data_bus[43]), .B2(n89), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n90), .B1(i_data_bus[45]), .B2(n89), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n82), .B1(i_data_bus[57]), .B2(n89), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n82), .B1(i_data_bus[59]), .B2(n89), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n82), .B1(i_data_bus[61]), .B2(n89), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n82), .B1(i_data_bus[63]), .B2(n89), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n90), .B1(i_data_bus[48]), .B2(n89), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n90), .B1(i_data_bus[47]), .B2(n89), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n90), .B1(i_data_bus[40]), .B2(n89), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n90), .B1(i_data_bus[42]), .B2(n89), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n90), .B1(i_data_bus[44]), .B2(n89), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U159 ( .A1(n91), .A2(n90), .B1(i_data_bus[46]), .B2(n89), 
        .ZN(N333) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_8 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96;

  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  INVD2BWP30P140 U3 ( .I(n15), .ZN(n59) );
  INVD3BWP30P140 U4 ( .I(n60), .ZN(n87) );
  NR2D1BWP30P140 U5 ( .A1(n42), .A2(n36), .ZN(n4) );
  INVD1BWP30P140 U6 ( .I(i_cmd[0]), .ZN(n36) );
  INVD2BWP30P140 U7 ( .I(i_valid[0]), .ZN(n5) );
  INVD1BWP30P140 U8 ( .I(n89), .ZN(n60) );
  ND2D1BWP30P140 U9 ( .A1(n7), .A2(n6), .ZN(N313) );
  INR2D2BWP30P140 U10 ( .A1(n37), .B1(i_cmd[0]), .ZN(n15) );
  INVD1BWP30P140 U11 ( .I(n24), .ZN(n34) );
  CKND2D2BWP30P140 U12 ( .A1(n44), .A2(n43), .ZN(n89) );
  NR2D1BWP30P140 U13 ( .A1(i_cmd[1]), .A2(n42), .ZN(n43) );
  INVD2BWP30P140 U14 ( .I(n24), .ZN(n58) );
  INVD2BWP30P140 U15 ( .I(n15), .ZN(n55) );
  BUFFD1BWP30P140 U16 ( .I(n89), .Z(n95) );
  INR2D2BWP30P140 U17 ( .A1(n38), .B1(n5), .ZN(n37) );
  ND2D1BWP30P140 U18 ( .A1(n1), .A2(i_en), .ZN(n42) );
  OAI22D1BWP30P140 U19 ( .A1(n32), .A2(n30), .B1(n59), .B2(n29), .ZN(N306) );
  OAI22D1BWP30P140 U20 ( .A1(n32), .A2(n31), .B1(n59), .B2(n81), .ZN(N307) );
  OAI22D1BWP30P140 U21 ( .A1(n34), .A2(n33), .B1(n59), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U22 ( .A1(n58), .A2(n35), .B1(n59), .B2(n79), .ZN(N309) );
  ND2OPTIBD1BWP30P140 U23 ( .A1(n15), .A2(i_data_bus[26]), .ZN(n6) );
  ND2OPTIBD1BWP30P140 U24 ( .A1(n24), .A2(i_data_bus[58]), .ZN(n7) );
  OAI22D1BWP30P140 U25 ( .A1(n34), .A2(n8), .B1(n59), .B2(n92), .ZN(N310) );
  OAI22D1BWP30P140 U26 ( .A1(n34), .A2(n9), .B1(n59), .B2(n91), .ZN(N311) );
  OAI22D1BWP30P140 U27 ( .A1(n34), .A2(n10), .B1(n59), .B2(n71), .ZN(N312) );
  OAI22D1BWP30P140 U28 ( .A1(n34), .A2(n11), .B1(n59), .B2(n83), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n34), .A2(n12), .B1(n59), .B2(n70), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n34), .A2(n13), .B1(n59), .B2(n72), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n34), .A2(n14), .B1(n59), .B2(n82), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n34), .A2(n61), .B1(n59), .B2(n63), .ZN(N318) );
  OAI22D1BWP30P140 U33 ( .A1(n32), .A2(n28), .B1(n55), .B2(n85), .ZN(N295) );
  OAI22D1BWP30P140 U34 ( .A1(n32), .A2(n27), .B1(n55), .B2(n65), .ZN(N296) );
  OAI22D1BWP30P140 U35 ( .A1(n32), .A2(n26), .B1(n55), .B2(n86), .ZN(N297) );
  OAI22D1BWP30P140 U36 ( .A1(n58), .A2(n25), .B1(n55), .B2(n67), .ZN(N298) );
  OAI22D1BWP30P140 U37 ( .A1(n32), .A2(n21), .B1(n55), .B2(n76), .ZN(N299) );
  OAI22D1BWP30P140 U38 ( .A1(n32), .A2(n20), .B1(n55), .B2(n75), .ZN(N300) );
  OAI22D1BWP30P140 U39 ( .A1(n32), .A2(n23), .B1(n55), .B2(n74), .ZN(N301) );
  OAI22D1BWP30P140 U40 ( .A1(n32), .A2(n22), .B1(n55), .B2(n78), .ZN(N302) );
  OAI22D1BWP30P140 U41 ( .A1(n32), .A2(n17), .B1(n55), .B2(n66), .ZN(N303) );
  OAI22D1BWP30P140 U42 ( .A1(n32), .A2(n16), .B1(n55), .B2(n77), .ZN(N304) );
  OAI22D1BWP30P140 U43 ( .A1(n32), .A2(n19), .B1(n55), .B2(n18), .ZN(N305) );
  ND2D1BWP30P140 U44 ( .A1(n46), .A2(n45), .ZN(N337) );
  ND2D1BWP30P140 U45 ( .A1(n94), .A2(i_data_bus[50]), .ZN(n45) );
  IND2D1BWP30P140 U46 ( .A1(n89), .B1(i_data_bus[18]), .ZN(n46) );
  ND2D1BWP30P140 U47 ( .A1(n48), .A2(n47), .ZN(N338) );
  ND2D1BWP30P140 U48 ( .A1(n94), .A2(i_data_bus[51]), .ZN(n47) );
  IND2D1BWP30P140 U49 ( .A1(n89), .B1(i_data_bus[19]), .ZN(n48) );
  INR2D6BWP30P140 U50 ( .A1(i_cmd[1]), .B1(n39), .ZN(n94) );
  INVD1BWP30P140 U51 ( .I(n94), .ZN(n62) );
  INVD1BWP30P140 U52 ( .I(rst), .ZN(n1) );
  INVD2BWP30P140 U53 ( .I(i_valid[1]), .ZN(n41) );
  MUX2NUD1BWP30P140 U54 ( .I0(n5), .I1(n41), .S(i_cmd[1]), .ZN(n2) );
  INVD2BWP30P140 U55 ( .I(n2), .ZN(n3) );
  INR2D4BWP30P140 U56 ( .A1(n4), .B1(n3), .ZN(n24) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[26]), .ZN(n84) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[55]), .ZN(n8) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[23]), .ZN(n92) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[56]), .ZN(n9) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[24]), .ZN(n91) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[57]), .ZN(n10) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[25]), .ZN(n71) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[59]), .ZN(n11) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[27]), .ZN(n83) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[60]), .ZN(n12) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[28]), .ZN(n70) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[61]), .ZN(n13) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[29]), .ZN(n72) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[62]), .ZN(n14) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[30]), .ZN(n82) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[63]), .ZN(n61) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[31]), .ZN(n63) );
  INVD2BWP30P140 U74 ( .I(n24), .ZN(n32) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[49]), .ZN(n16) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[17]), .ZN(n77) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[48]), .ZN(n17) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[16]), .ZN(n66) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[50]), .ZN(n19) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[18]), .ZN(n18) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[45]), .ZN(n20) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[13]), .ZN(n75) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[44]), .ZN(n21) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[12]), .ZN(n76) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[47]), .ZN(n22) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[15]), .ZN(n78) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[46]), .ZN(n23) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[14]), .ZN(n74) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[43]), .ZN(n25) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[11]), .ZN(n67) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[42]), .ZN(n26) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[10]), .ZN(n86) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[41]), .ZN(n27) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[9]), .ZN(n65) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[40]), .ZN(n28) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[8]), .ZN(n85) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[51]), .ZN(n30) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[19]), .ZN(n29) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[52]), .ZN(n31) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[20]), .ZN(n81) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[53]), .ZN(n33) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[54]), .ZN(n35) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[22]), .ZN(n79) );
  OAI31D1BWP30P140 U105 ( .A1(n42), .A2(n41), .A3(n36), .B(n59), .ZN(N353) );
  INVD1BWP30P140 U106 ( .I(n37), .ZN(n40) );
  INVD1BWP30P140 U107 ( .I(n42), .ZN(n38) );
  ND2OPTIBD1BWP30P140 U108 ( .A1(i_valid[1]), .A2(n38), .ZN(n39) );
  OAI21D1BWP30P140 U109 ( .A1(n40), .A2(i_cmd[1]), .B(n62), .ZN(N354) );
  MUX2NUD1BWP30P140 U110 ( .I0(n5), .I1(n41), .S(i_cmd[0]), .ZN(n44) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[39]), .ZN(n49) );
  OAI22D1BWP30P140 U113 ( .A1(n55), .A2(n64), .B1(n58), .B2(n49), .ZN(N294) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[0]), .ZN(n93) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[32]), .ZN(n50) );
  OAI22D1BWP30P140 U116 ( .A1(n59), .A2(n93), .B1(n58), .B2(n50), .ZN(N287) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[3]), .ZN(n90) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[35]), .ZN(n51) );
  OAI22D1BWP30P140 U119 ( .A1(n59), .A2(n90), .B1(n58), .B2(n51), .ZN(N290) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[4]), .ZN(n88) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[36]), .ZN(n52) );
  OAI22D1BWP30P140 U122 ( .A1(n55), .A2(n88), .B1(n58), .B2(n52), .ZN(N291) );
  INVD1BWP30P140 U123 ( .I(i_data_bus[2]), .ZN(n96) );
  INVD1BWP30P140 U124 ( .I(i_data_bus[34]), .ZN(n53) );
  OAI22D1BWP30P140 U125 ( .A1(n59), .A2(n96), .B1(n58), .B2(n53), .ZN(N289) );
  INVD1BWP30P140 U126 ( .I(i_data_bus[6]), .ZN(n73) );
  INVD1BWP30P140 U127 ( .I(i_data_bus[38]), .ZN(n54) );
  OAI22D1BWP30P140 U128 ( .A1(n55), .A2(n73), .B1(n58), .B2(n54), .ZN(N293) );
  INVD1BWP30P140 U129 ( .I(i_data_bus[5]), .ZN(n68) );
  INVD1BWP30P140 U130 ( .I(i_data_bus[37]), .ZN(n56) );
  OAI22D1BWP30P140 U131 ( .A1(n59), .A2(n68), .B1(n58), .B2(n56), .ZN(N292) );
  INVD1BWP30P140 U132 ( .I(i_data_bus[1]), .ZN(n69) );
  INVD1BWP30P140 U133 ( .I(i_data_bus[33]), .ZN(n57) );
  OAI22D1BWP30P140 U134 ( .A1(n59), .A2(n69), .B1(n58), .B2(n57), .ZN(N288) );
  OAI22D1BWP30P140 U135 ( .A1(n87), .A2(n63), .B1(n62), .B2(n61), .ZN(N350) );
  MOAI22D1BWP30P140 U136 ( .A1(n64), .A2(n87), .B1(i_data_bus[39]), .B2(n94), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U137 ( .A1(n65), .A2(n95), .B1(i_data_bus[41]), .B2(n94), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n66), .A2(n87), .B1(i_data_bus[48]), .B2(n94), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U139 ( .A1(n67), .A2(n87), .B1(i_data_bus[43]), .B2(n94), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n68), .A2(n87), .B1(i_data_bus[37]), .B2(n94), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U141 ( .A1(n69), .A2(n87), .B1(i_data_bus[33]), .B2(n94), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U142 ( .A1(n70), .A2(n87), .B1(i_data_bus[60]), .B2(n94), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U143 ( .A1(n71), .A2(n87), .B1(i_data_bus[57]), .B2(n94), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U144 ( .A1(n72), .A2(n87), .B1(i_data_bus[61]), .B2(n94), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U145 ( .A1(n73), .A2(n87), .B1(i_data_bus[38]), .B2(n94), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U146 ( .A1(n74), .A2(n87), .B1(i_data_bus[46]), .B2(n94), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U147 ( .A1(n75), .A2(n87), .B1(i_data_bus[45]), .B2(n94), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U148 ( .A1(n76), .A2(n87), .B1(i_data_bus[44]), .B2(n94), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U149 ( .A1(n77), .A2(n95), .B1(i_data_bus[49]), .B2(n94), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U150 ( .A1(n78), .A2(n87), .B1(i_data_bus[47]), .B2(n94), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U151 ( .A1(n79), .A2(n87), .B1(i_data_bus[54]), .B2(n94), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n80), .A2(n87), .B1(i_data_bus[53]), .B2(n94), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U153 ( .A1(n81), .A2(n87), .B1(i_data_bus[52]), .B2(n94), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U154 ( .A1(n82), .A2(n87), .B1(i_data_bus[62]), .B2(n94), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U155 ( .A1(n83), .A2(n87), .B1(i_data_bus[59]), .B2(n94), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U156 ( .A1(n84), .A2(n87), .B1(i_data_bus[58]), .B2(n94), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U157 ( .A1(n85), .A2(n87), .B1(i_data_bus[40]), .B2(n94), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U158 ( .A1(n86), .A2(n87), .B1(i_data_bus[42]), .B2(n94), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n88), .A2(n95), .B1(i_data_bus[36]), .B2(n94), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n87), .B1(i_data_bus[35]), .B2(n94), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U161 ( .A1(n91), .A2(n87), .B1(i_data_bus[56]), .B2(n94), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U162 ( .A1(n92), .A2(n87), .B1(i_data_bus[55]), .B2(n94), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U163 ( .A1(n93), .A2(n87), .B1(i_data_bus[32]), .B2(n94), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U164 ( .A1(n96), .A2(n87), .B1(i_data_bus[34]), .B2(n94), 
        .ZN(N321) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_9 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n18), .Z(n89) );
  CKND2D3BWP30P140 U4 ( .A1(n5), .A2(n4), .ZN(n47) );
  NR2D1BWP30P140 U5 ( .A1(n49), .A2(i_cmd[1]), .ZN(n53) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n49), .ZN(n17) );
  INVD1BWP30P140 U7 ( .I(i_cmd[0]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U8 ( .A1(n17), .A2(n3), .ZN(n2) );
  ND2D1BWP30P140 U9 ( .A1(n1), .A2(i_en), .ZN(n49) );
  INVD1BWP30P140 U10 ( .I(n47), .ZN(n6) );
  INVD1BWP30P140 U11 ( .I(n77), .ZN(n62) );
  INVD1BWP30P140 U12 ( .I(n89), .ZN(n19) );
  INVD1BWP30P140 U13 ( .I(n2), .ZN(n11) );
  INVD1BWP30P140 U14 ( .I(rst), .ZN(n1) );
  INVD2BWP30P140 U15 ( .I(i_valid[1]), .ZN(n50) );
  INVD2BWP30P140 U16 ( .I(n11), .ZN(n48) );
  OAI31D1BWP30P140 U17 ( .A1(n49), .A2(n50), .A3(n3), .B(n48), .ZN(N353) );
  INVD1BWP30P140 U18 ( .I(i_data_bus[0]), .ZN(n55) );
  INVD1BWP30P140 U19 ( .I(i_valid[0]), .ZN(n51) );
  MUX2NOPTD2BWP30P140 U20 ( .I0(n51), .I1(n50), .S(i_cmd[1]), .ZN(n5) );
  NR2OPTPAD1BWP30P140 U21 ( .A1(n49), .A2(n3), .ZN(n4) );
  INVD2BWP30P140 U22 ( .I(n6), .ZN(n16) );
  INVD1BWP30P140 U23 ( .I(i_data_bus[32]), .ZN(n7) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n55), .B1(n16), .B2(n7), .ZN(N287) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[1]), .ZN(n56) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[33]), .ZN(n8) );
  OAI22D1BWP30P140 U27 ( .A1(n48), .A2(n56), .B1(n16), .B2(n8), .ZN(N288) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[34]), .ZN(n9) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n59), .B1(n16), .B2(n9), .ZN(N289) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[35]), .ZN(n10) );
  OAI22D1BWP30P140 U33 ( .A1(n48), .A2(n60), .B1(n16), .B2(n10), .ZN(N290) );
  INVD2BWP30P140 U34 ( .I(n11), .ZN(n32) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[36]), .ZN(n12) );
  OAI22D1BWP30P140 U37 ( .A1(n32), .A2(n61), .B1(n16), .B2(n12), .ZN(N291) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[5]), .ZN(n63) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[37]), .ZN(n13) );
  OAI22D1BWP30P140 U40 ( .A1(n32), .A2(n63), .B1(n16), .B2(n13), .ZN(N292) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[38]), .ZN(n14) );
  OAI22D1BWP30P140 U43 ( .A1(n32), .A2(n58), .B1(n16), .B2(n14), .ZN(N293) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[39]), .ZN(n15) );
  OAI22D1BWP30P140 U46 ( .A1(n32), .A2(n57), .B1(n16), .B2(n15), .ZN(N294) );
  INVD1BWP30P140 U47 ( .I(n17), .ZN(n20) );
  INVD1BWP30P140 U48 ( .I(n49), .ZN(n18) );
  OAI21D1BWP30P140 U49 ( .A1(n20), .A2(i_cmd[1]), .B(n19), .ZN(N354) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[8]), .ZN(n64) );
  BUFFD4BWP30P140 U51 ( .I(n47), .Z(n44) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[40]), .ZN(n21) );
  OAI22D1BWP30P140 U53 ( .A1(n32), .A2(n64), .B1(n44), .B2(n21), .ZN(N295) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[9]), .ZN(n65) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[41]), .ZN(n22) );
  OAI22D1BWP30P140 U56 ( .A1(n32), .A2(n65), .B1(n44), .B2(n22), .ZN(N296) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[10]), .ZN(n66) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[42]), .ZN(n23) );
  OAI22D1BWP30P140 U59 ( .A1(n32), .A2(n66), .B1(n44), .B2(n23), .ZN(N297) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[11]), .ZN(n67) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[43]), .ZN(n24) );
  OAI22D1BWP30P140 U62 ( .A1(n32), .A2(n67), .B1(n44), .B2(n24), .ZN(N298) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[12]), .ZN(n68) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[44]), .ZN(n25) );
  OAI22D1BWP30P140 U65 ( .A1(n32), .A2(n68), .B1(n44), .B2(n25), .ZN(N299) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[13]), .ZN(n69) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[45]), .ZN(n26) );
  OAI22D1BWP30P140 U68 ( .A1(n32), .A2(n69), .B1(n44), .B2(n26), .ZN(N300) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[14]), .ZN(n70) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[46]), .ZN(n27) );
  OAI22D1BWP30P140 U71 ( .A1(n32), .A2(n70), .B1(n44), .B2(n27), .ZN(N301) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[15]), .ZN(n71) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[47]), .ZN(n28) );
  OAI22D1BWP30P140 U74 ( .A1(n32), .A2(n71), .B1(n44), .B2(n28), .ZN(N302) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[16]), .ZN(n72) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[48]), .ZN(n29) );
  OAI22D1BWP30P140 U77 ( .A1(n32), .A2(n72), .B1(n44), .B2(n29), .ZN(N303) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[17]), .ZN(n73) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[49]), .ZN(n30) );
  OAI22D1BWP30P140 U80 ( .A1(n32), .A2(n73), .B1(n44), .B2(n30), .ZN(N304) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[18]), .ZN(n74) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[50]), .ZN(n31) );
  OAI22D1BWP30P140 U83 ( .A1(n32), .A2(n74), .B1(n44), .B2(n31), .ZN(N305) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[19]), .ZN(n76) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[51]), .ZN(n33) );
  OAI22D1BWP30P140 U86 ( .A1(n48), .A2(n76), .B1(n44), .B2(n33), .ZN(N306) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[20]), .ZN(n78) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[52]), .ZN(n34) );
  OAI22D1BWP30P140 U89 ( .A1(n48), .A2(n78), .B1(n44), .B2(n34), .ZN(N307) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[21]), .ZN(n79) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[53]), .ZN(n35) );
  OAI22D1BWP30P140 U92 ( .A1(n48), .A2(n79), .B1(n44), .B2(n35), .ZN(N308) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[22]), .ZN(n80) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[54]), .ZN(n36) );
  OAI22D1BWP30P140 U95 ( .A1(n48), .A2(n80), .B1(n44), .B2(n36), .ZN(N309) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[23]), .ZN(n81) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[55]), .ZN(n37) );
  OAI22D1BWP30P140 U98 ( .A1(n48), .A2(n81), .B1(n44), .B2(n37), .ZN(N310) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[24]), .ZN(n82) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[56]), .ZN(n38) );
  OAI22D1BWP30P140 U101 ( .A1(n48), .A2(n82), .B1(n44), .B2(n38), .ZN(N311) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[25]), .ZN(n83) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[57]), .ZN(n39) );
  OAI22D1BWP30P140 U104 ( .A1(n48), .A2(n83), .B1(n44), .B2(n39), .ZN(N312) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[26]), .ZN(n84) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[58]), .ZN(n40) );
  OAI22D1BWP30P140 U107 ( .A1(n48), .A2(n84), .B1(n44), .B2(n40), .ZN(N313) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[27]), .ZN(n85) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[59]), .ZN(n41) );
  OAI22D1BWP30P140 U110 ( .A1(n48), .A2(n85), .B1(n44), .B2(n41), .ZN(N314) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[28]), .ZN(n86) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[60]), .ZN(n42) );
  OAI22D1BWP30P140 U113 ( .A1(n48), .A2(n86), .B1(n44), .B2(n42), .ZN(N315) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[29]), .ZN(n87) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[61]), .ZN(n43) );
  OAI22D1BWP30P140 U116 ( .A1(n48), .A2(n87), .B1(n44), .B2(n43), .ZN(N316) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[30]), .ZN(n88) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[62]), .ZN(n45) );
  OAI22D1BWP30P140 U119 ( .A1(n48), .A2(n88), .B1(n47), .B2(n45), .ZN(N317) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[31]), .ZN(n91) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[63]), .ZN(n46) );
  OAI22D1BWP30P140 U122 ( .A1(n48), .A2(n91), .B1(n47), .B2(n46), .ZN(N318) );
  MUX2NUD1BWP30P140 U123 ( .I0(n51), .I1(n50), .S(i_cmd[0]), .ZN(n52) );
  ND2OPTIBD1BWP30P140 U124 ( .A1(n53), .A2(n52), .ZN(n54) );
  INVD2BWP30P140 U125 ( .I(n54), .ZN(n77) );
  MOAI22D1BWP30P140 U126 ( .A1(n55), .A2(n62), .B1(i_data_bus[32]), .B2(n89), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n62), .B1(i_data_bus[33]), .B2(n89), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n62), .B1(i_data_bus[39]), .B2(n89), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n62), .B1(i_data_bus[38]), .B2(n89), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n62), .B1(i_data_bus[34]), .B2(n89), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n62), .B1(i_data_bus[35]), .B2(n89), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n90), .B1(i_data_bus[36]), .B2(n89), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n75), .B1(i_data_bus[37]), .B2(n89), 
        .ZN(N324) );
  INVD2BWP30P140 U134 ( .I(n77), .ZN(n75) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n90), .B1(i_data_bus[40]), .B2(n89), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n75), .B1(i_data_bus[41]), .B2(n89), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n90), .B1(i_data_bus[42]), .B2(n89), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n75), .B1(i_data_bus[43]), .B2(n89), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n90), .B1(i_data_bus[44]), .B2(n89), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n75), .B1(i_data_bus[45]), .B2(n89), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n90), .B1(i_data_bus[46]), .B2(n89), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n75), .B1(i_data_bus[47]), .B2(n89), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n90), .B1(i_data_bus[48]), .B2(n89), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n75), .B1(i_data_bus[49]), .B2(n89), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n90), .B1(i_data_bus[50]), .B2(n89), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U146 ( .A1(n76), .A2(n75), .B1(i_data_bus[51]), .B2(n89), 
        .ZN(N338) );
  INVD2BWP30P140 U147 ( .I(n77), .ZN(n90) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n90), .B1(i_data_bus[52]), .B2(n89), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n75), .B1(i_data_bus[53]), .B2(n89), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n90), .B1(i_data_bus[54]), .B2(n89), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n75), .B1(i_data_bus[55]), .B2(n89), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n90), .B1(i_data_bus[56]), .B2(n89), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n75), .B1(i_data_bus[57]), .B2(n89), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n90), .B1(i_data_bus[58]), .B2(n89), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n75), .B1(i_data_bus[59]), .B2(n89), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n90), .B1(i_data_bus[60]), .B2(n89), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n75), .B1(i_data_bus[61]), .B2(n89), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n90), .B1(i_data_bus[62]), .B2(n89), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U159 ( .A1(n91), .A2(n75), .B1(i_data_bus[63]), .B2(n89), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_10 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n18), .Z(n89) );
  CKND2D3BWP30P140 U4 ( .A1(n5), .A2(n4), .ZN(n47) );
  NR2D1BWP30P140 U5 ( .A1(n49), .A2(i_cmd[1]), .ZN(n53) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n49), .ZN(n17) );
  NR2D1BWP30P140 U7 ( .A1(n49), .A2(n3), .ZN(n4) );
  ND2OPTIBD1BWP30P140 U8 ( .A1(n17), .A2(n3), .ZN(n2) );
  ND2D1BWP30P140 U9 ( .A1(n1), .A2(i_en), .ZN(n49) );
  INVD1BWP30P140 U10 ( .I(n47), .ZN(n6) );
  INVD1BWP30P140 U11 ( .I(n77), .ZN(n62) );
  INVD1BWP30P140 U12 ( .I(n89), .ZN(n19) );
  INVD1BWP30P140 U13 ( .I(n2), .ZN(n11) );
  INVD1BWP30P140 U14 ( .I(rst), .ZN(n1) );
  INVD2BWP30P140 U15 ( .I(i_valid[1]), .ZN(n50) );
  INVD2BWP30P140 U16 ( .I(i_cmd[0]), .ZN(n3) );
  INVD2BWP30P140 U17 ( .I(n11), .ZN(n48) );
  OAI31D1BWP30P140 U18 ( .A1(n49), .A2(n50), .A3(n3), .B(n48), .ZN(N353) );
  INVD1BWP30P140 U19 ( .I(i_data_bus[0]), .ZN(n55) );
  INVD1BWP30P140 U20 ( .I(i_valid[0]), .ZN(n51) );
  MUX2NOPTD2BWP30P140 U21 ( .I0(n51), .I1(n50), .S(i_cmd[1]), .ZN(n5) );
  INVD2BWP30P140 U22 ( .I(n6), .ZN(n16) );
  INVD1BWP30P140 U23 ( .I(i_data_bus[32]), .ZN(n7) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n55), .B1(n16), .B2(n7), .ZN(N287) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[1]), .ZN(n56) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[33]), .ZN(n8) );
  OAI22D1BWP30P140 U27 ( .A1(n48), .A2(n56), .B1(n16), .B2(n8), .ZN(N288) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[2]), .ZN(n57) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[34]), .ZN(n9) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n57), .B1(n16), .B2(n9), .ZN(N289) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[3]), .ZN(n58) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[35]), .ZN(n10) );
  OAI22D1BWP30P140 U33 ( .A1(n48), .A2(n58), .B1(n16), .B2(n10), .ZN(N290) );
  INVD2BWP30P140 U34 ( .I(n11), .ZN(n32) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[36]), .ZN(n12) );
  OAI22D1BWP30P140 U37 ( .A1(n32), .A2(n59), .B1(n16), .B2(n12), .ZN(N291) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[5]), .ZN(n60) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[37]), .ZN(n13) );
  OAI22D1BWP30P140 U40 ( .A1(n32), .A2(n60), .B1(n16), .B2(n13), .ZN(N292) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[6]), .ZN(n61) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[38]), .ZN(n14) );
  OAI22D1BWP30P140 U43 ( .A1(n32), .A2(n61), .B1(n16), .B2(n14), .ZN(N293) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[7]), .ZN(n63) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[39]), .ZN(n15) );
  OAI22D1BWP30P140 U46 ( .A1(n32), .A2(n63), .B1(n16), .B2(n15), .ZN(N294) );
  INVD1BWP30P140 U47 ( .I(n17), .ZN(n20) );
  INVD1BWP30P140 U48 ( .I(n49), .ZN(n18) );
  OAI21D1BWP30P140 U49 ( .A1(n20), .A2(i_cmd[1]), .B(n19), .ZN(N354) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[8]), .ZN(n91) );
  BUFFD4BWP30P140 U51 ( .I(n47), .Z(n44) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[40]), .ZN(n21) );
  OAI22D1BWP30P140 U53 ( .A1(n32), .A2(n91), .B1(n44), .B2(n21), .ZN(N295) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[9]), .ZN(n88) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[41]), .ZN(n22) );
  OAI22D1BWP30P140 U56 ( .A1(n32), .A2(n88), .B1(n44), .B2(n22), .ZN(N296) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[10]), .ZN(n87) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[42]), .ZN(n23) );
  OAI22D1BWP30P140 U59 ( .A1(n32), .A2(n87), .B1(n44), .B2(n23), .ZN(N297) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[11]), .ZN(n86) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[43]), .ZN(n24) );
  OAI22D1BWP30P140 U62 ( .A1(n32), .A2(n86), .B1(n44), .B2(n24), .ZN(N298) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[12]), .ZN(n85) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[44]), .ZN(n25) );
  OAI22D1BWP30P140 U65 ( .A1(n32), .A2(n85), .B1(n44), .B2(n25), .ZN(N299) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[13]), .ZN(n84) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[45]), .ZN(n26) );
  OAI22D1BWP30P140 U68 ( .A1(n32), .A2(n84), .B1(n44), .B2(n26), .ZN(N300) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[14]), .ZN(n83) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[46]), .ZN(n27) );
  OAI22D1BWP30P140 U71 ( .A1(n32), .A2(n83), .B1(n44), .B2(n27), .ZN(N301) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[15]), .ZN(n82) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[47]), .ZN(n28) );
  OAI22D1BWP30P140 U74 ( .A1(n32), .A2(n82), .B1(n44), .B2(n28), .ZN(N302) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[16]), .ZN(n81) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[48]), .ZN(n29) );
  OAI22D1BWP30P140 U77 ( .A1(n32), .A2(n81), .B1(n44), .B2(n29), .ZN(N303) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[17]), .ZN(n80) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[49]), .ZN(n30) );
  OAI22D1BWP30P140 U80 ( .A1(n32), .A2(n80), .B1(n44), .B2(n30), .ZN(N304) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[18]), .ZN(n79) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[50]), .ZN(n31) );
  OAI22D1BWP30P140 U83 ( .A1(n32), .A2(n79), .B1(n44), .B2(n31), .ZN(N305) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[51]), .ZN(n33) );
  OAI22D1BWP30P140 U86 ( .A1(n48), .A2(n78), .B1(n44), .B2(n33), .ZN(N306) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[20]), .ZN(n76) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[52]), .ZN(n34) );
  OAI22D1BWP30P140 U89 ( .A1(n48), .A2(n76), .B1(n44), .B2(n34), .ZN(N307) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[21]), .ZN(n74) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[53]), .ZN(n35) );
  OAI22D1BWP30P140 U92 ( .A1(n48), .A2(n74), .B1(n44), .B2(n35), .ZN(N308) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[22]), .ZN(n73) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[54]), .ZN(n36) );
  OAI22D1BWP30P140 U95 ( .A1(n48), .A2(n73), .B1(n44), .B2(n36), .ZN(N309) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[23]), .ZN(n72) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[55]), .ZN(n37) );
  OAI22D1BWP30P140 U98 ( .A1(n48), .A2(n72), .B1(n44), .B2(n37), .ZN(N310) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[24]), .ZN(n71) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[56]), .ZN(n38) );
  OAI22D1BWP30P140 U101 ( .A1(n48), .A2(n71), .B1(n44), .B2(n38), .ZN(N311) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[25]), .ZN(n70) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[57]), .ZN(n39) );
  OAI22D1BWP30P140 U104 ( .A1(n48), .A2(n70), .B1(n44), .B2(n39), .ZN(N312) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[26]), .ZN(n69) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[58]), .ZN(n40) );
  OAI22D1BWP30P140 U107 ( .A1(n48), .A2(n69), .B1(n44), .B2(n40), .ZN(N313) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[27]), .ZN(n68) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[59]), .ZN(n41) );
  OAI22D1BWP30P140 U110 ( .A1(n48), .A2(n68), .B1(n44), .B2(n41), .ZN(N314) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[28]), .ZN(n67) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[60]), .ZN(n42) );
  OAI22D1BWP30P140 U113 ( .A1(n48), .A2(n67), .B1(n44), .B2(n42), .ZN(N315) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[29]), .ZN(n66) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[61]), .ZN(n43) );
  OAI22D1BWP30P140 U116 ( .A1(n48), .A2(n66), .B1(n44), .B2(n43), .ZN(N316) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[30]), .ZN(n65) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[62]), .ZN(n45) );
  OAI22D1BWP30P140 U119 ( .A1(n48), .A2(n65), .B1(n47), .B2(n45), .ZN(N317) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[31]), .ZN(n64) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[63]), .ZN(n46) );
  OAI22D1BWP30P140 U122 ( .A1(n48), .A2(n64), .B1(n47), .B2(n46), .ZN(N318) );
  MUX2NUD1BWP30P140 U123 ( .I0(n51), .I1(n50), .S(i_cmd[0]), .ZN(n52) );
  ND2OPTIBD1BWP30P140 U124 ( .A1(n53), .A2(n52), .ZN(n54) );
  INVD2BWP30P140 U125 ( .I(n54), .ZN(n77) );
  MOAI22D1BWP30P140 U126 ( .A1(n55), .A2(n62), .B1(i_data_bus[32]), .B2(n89), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n62), .B1(i_data_bus[33]), .B2(n89), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n62), .B1(i_data_bus[34]), .B2(n89), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n62), .B1(i_data_bus[35]), .B2(n89), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n62), .B1(i_data_bus[36]), .B2(n89), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n62), .B1(i_data_bus[37]), .B2(n89), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n90), .B1(i_data_bus[38]), .B2(n89), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n75), .B1(i_data_bus[39]), .B2(n89), 
        .ZN(N326) );
  INVD2BWP30P140 U134 ( .I(n77), .ZN(n75) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n90), .B1(i_data_bus[63]), .B2(n89), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n75), .B1(i_data_bus[62]), .B2(n89), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n90), .B1(i_data_bus[61]), .B2(n89), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n75), .B1(i_data_bus[60]), .B2(n89), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n90), .B1(i_data_bus[59]), .B2(n89), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n75), .B1(i_data_bus[58]), .B2(n89), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n90), .B1(i_data_bus[57]), .B2(n89), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n75), .B1(i_data_bus[56]), .B2(n89), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n90), .B1(i_data_bus[55]), .B2(n89), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n75), .B1(i_data_bus[54]), .B2(n89), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n90), .B1(i_data_bus[53]), .B2(n89), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U146 ( .A1(n76), .A2(n75), .B1(i_data_bus[52]), .B2(n89), 
        .ZN(N339) );
  INVD2BWP30P140 U147 ( .I(n77), .ZN(n90) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n90), .B1(i_data_bus[51]), .B2(n89), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n75), .B1(i_data_bus[50]), .B2(n89), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n90), .B1(i_data_bus[49]), .B2(n89), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n75), .B1(i_data_bus[48]), .B2(n89), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n90), .B1(i_data_bus[47]), .B2(n89), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n75), .B1(i_data_bus[46]), .B2(n89), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n90), .B1(i_data_bus[45]), .B2(n89), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n75), .B1(i_data_bus[44]), .B2(n89), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n90), .B1(i_data_bus[43]), .B2(n89), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n75), .B1(i_data_bus[42]), .B2(n89), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n90), .B1(i_data_bus[41]), .B2(n89), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U159 ( .A1(n91), .A2(n75), .B1(i_data_bus[40]), .B2(n89), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_11 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n18), .Z(n89) );
  CKND2D3BWP30P140 U4 ( .A1(n5), .A2(n4), .ZN(n47) );
  NR2D1BWP30P140 U5 ( .A1(n49), .A2(i_cmd[1]), .ZN(n53) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n49), .ZN(n17) );
  INVD1BWP30P140 U7 ( .I(i_cmd[0]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U8 ( .A1(n17), .A2(n3), .ZN(n2) );
  ND2D1BWP30P140 U9 ( .A1(n1), .A2(i_en), .ZN(n49) );
  INVD1BWP30P140 U10 ( .I(n47), .ZN(n6) );
  INVD1BWP30P140 U11 ( .I(n77), .ZN(n62) );
  INVD1BWP30P140 U12 ( .I(n89), .ZN(n19) );
  INVD1BWP30P140 U13 ( .I(n2), .ZN(n11) );
  INVD1BWP30P140 U14 ( .I(rst), .ZN(n1) );
  INVD2BWP30P140 U15 ( .I(i_valid[1]), .ZN(n50) );
  INVD2BWP30P140 U16 ( .I(n11), .ZN(n48) );
  OAI31D1BWP30P140 U17 ( .A1(n49), .A2(n50), .A3(n3), .B(n48), .ZN(N353) );
  INVD1BWP30P140 U18 ( .I(i_data_bus[0]), .ZN(n55) );
  INVD1BWP30P140 U19 ( .I(i_valid[0]), .ZN(n51) );
  MUX2NOPTD2BWP30P140 U20 ( .I0(n51), .I1(n50), .S(i_cmd[1]), .ZN(n5) );
  NR2OPTPAD1BWP30P140 U21 ( .A1(n49), .A2(n3), .ZN(n4) );
  INVD2BWP30P140 U22 ( .I(n6), .ZN(n16) );
  INVD1BWP30P140 U23 ( .I(i_data_bus[32]), .ZN(n7) );
  OAI22D1BWP30P140 U24 ( .A1(n41), .A2(n55), .B1(n16), .B2(n7), .ZN(N287) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[1]), .ZN(n56) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[33]), .ZN(n8) );
  OAI22D1BWP30P140 U27 ( .A1(n48), .A2(n56), .B1(n16), .B2(n8), .ZN(N288) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[2]), .ZN(n57) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[34]), .ZN(n9) );
  OAI22D1BWP30P140 U30 ( .A1(n41), .A2(n57), .B1(n16), .B2(n9), .ZN(N289) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[3]), .ZN(n58) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[35]), .ZN(n10) );
  OAI22D1BWP30P140 U33 ( .A1(n48), .A2(n58), .B1(n16), .B2(n10), .ZN(N290) );
  INVD2BWP30P140 U34 ( .I(n11), .ZN(n41) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[36]), .ZN(n12) );
  OAI22D1BWP30P140 U37 ( .A1(n41), .A2(n59), .B1(n16), .B2(n12), .ZN(N291) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[5]), .ZN(n60) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[37]), .ZN(n13) );
  OAI22D1BWP30P140 U40 ( .A1(n41), .A2(n60), .B1(n16), .B2(n13), .ZN(N292) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[6]), .ZN(n61) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[38]), .ZN(n14) );
  OAI22D1BWP30P140 U43 ( .A1(n41), .A2(n61), .B1(n16), .B2(n14), .ZN(N293) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[7]), .ZN(n63) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[39]), .ZN(n15) );
  OAI22D1BWP30P140 U46 ( .A1(n41), .A2(n63), .B1(n16), .B2(n15), .ZN(N294) );
  INVD1BWP30P140 U47 ( .I(n17), .ZN(n20) );
  INVD1BWP30P140 U48 ( .I(n49), .ZN(n18) );
  OAI21D1BWP30P140 U49 ( .A1(n20), .A2(i_cmd[1]), .B(n19), .ZN(N354) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[24]), .ZN(n71) );
  BUFFD4BWP30P140 U51 ( .I(n47), .Z(n44) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[56]), .ZN(n21) );
  OAI22D1BWP30P140 U53 ( .A1(n48), .A2(n71), .B1(n44), .B2(n21), .ZN(N311) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[25]), .ZN(n70) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[57]), .ZN(n22) );
  OAI22D1BWP30P140 U56 ( .A1(n48), .A2(n70), .B1(n44), .B2(n22), .ZN(N312) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[26]), .ZN(n69) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[58]), .ZN(n23) );
  OAI22D1BWP30P140 U59 ( .A1(n48), .A2(n69), .B1(n44), .B2(n23), .ZN(N313) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[27]), .ZN(n68) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[59]), .ZN(n24) );
  OAI22D1BWP30P140 U62 ( .A1(n48), .A2(n68), .B1(n44), .B2(n24), .ZN(N314) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[28]), .ZN(n67) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[60]), .ZN(n25) );
  OAI22D1BWP30P140 U65 ( .A1(n48), .A2(n67), .B1(n44), .B2(n25), .ZN(N315) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[29]), .ZN(n66) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[61]), .ZN(n26) );
  OAI22D1BWP30P140 U68 ( .A1(n48), .A2(n66), .B1(n44), .B2(n26), .ZN(N316) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[30]), .ZN(n65) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[62]), .ZN(n27) );
  OAI22D1BWP30P140 U71 ( .A1(n48), .A2(n65), .B1(n44), .B2(n27), .ZN(N317) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[31]), .ZN(n64) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[63]), .ZN(n28) );
  OAI22D1BWP30P140 U74 ( .A1(n48), .A2(n64), .B1(n44), .B2(n28), .ZN(N318) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[23]), .ZN(n72) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[55]), .ZN(n29) );
  OAI22D1BWP30P140 U77 ( .A1(n48), .A2(n72), .B1(n44), .B2(n29), .ZN(N310) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[8]), .ZN(n91) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[40]), .ZN(n30) );
  OAI22D1BWP30P140 U80 ( .A1(n41), .A2(n91), .B1(n44), .B2(n30), .ZN(N295) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[9]), .ZN(n88) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[41]), .ZN(n31) );
  OAI22D1BWP30P140 U83 ( .A1(n41), .A2(n88), .B1(n44), .B2(n31), .ZN(N296) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[10]), .ZN(n87) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[42]), .ZN(n32) );
  OAI22D1BWP30P140 U86 ( .A1(n41), .A2(n87), .B1(n44), .B2(n32), .ZN(N297) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[11]), .ZN(n86) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[43]), .ZN(n33) );
  OAI22D1BWP30P140 U89 ( .A1(n41), .A2(n86), .B1(n44), .B2(n33), .ZN(N298) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[12]), .ZN(n85) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[44]), .ZN(n34) );
  OAI22D1BWP30P140 U92 ( .A1(n41), .A2(n85), .B1(n44), .B2(n34), .ZN(N299) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[13]), .ZN(n84) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[45]), .ZN(n35) );
  OAI22D1BWP30P140 U95 ( .A1(n41), .A2(n84), .B1(n44), .B2(n35), .ZN(N300) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[14]), .ZN(n83) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[46]), .ZN(n36) );
  OAI22D1BWP30P140 U98 ( .A1(n41), .A2(n83), .B1(n44), .B2(n36), .ZN(N301) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[15]), .ZN(n82) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[47]), .ZN(n37) );
  OAI22D1BWP30P140 U101 ( .A1(n41), .A2(n82), .B1(n44), .B2(n37), .ZN(N302) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[16]), .ZN(n81) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[48]), .ZN(n38) );
  OAI22D1BWP30P140 U104 ( .A1(n41), .A2(n81), .B1(n44), .B2(n38), .ZN(N303) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[17]), .ZN(n80) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[49]), .ZN(n39) );
  OAI22D1BWP30P140 U107 ( .A1(n41), .A2(n80), .B1(n44), .B2(n39), .ZN(N304) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[18]), .ZN(n79) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[50]), .ZN(n40) );
  OAI22D1BWP30P140 U110 ( .A1(n41), .A2(n79), .B1(n44), .B2(n40), .ZN(N305) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[51]), .ZN(n42) );
  OAI22D1BWP30P140 U113 ( .A1(n48), .A2(n78), .B1(n44), .B2(n42), .ZN(N306) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[20]), .ZN(n76) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[52]), .ZN(n43) );
  OAI22D1BWP30P140 U116 ( .A1(n48), .A2(n76), .B1(n44), .B2(n43), .ZN(N307) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[21]), .ZN(n74) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[53]), .ZN(n45) );
  OAI22D1BWP30P140 U119 ( .A1(n48), .A2(n74), .B1(n47), .B2(n45), .ZN(N308) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[22]), .ZN(n73) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[54]), .ZN(n46) );
  OAI22D1BWP30P140 U122 ( .A1(n48), .A2(n73), .B1(n47), .B2(n46), .ZN(N309) );
  MUX2NUD1BWP30P140 U123 ( .I0(n51), .I1(n50), .S(i_cmd[0]), .ZN(n52) );
  ND2OPTIBD1BWP30P140 U124 ( .A1(n53), .A2(n52), .ZN(n54) );
  INVD2BWP30P140 U125 ( .I(n54), .ZN(n77) );
  MOAI22D1BWP30P140 U126 ( .A1(n55), .A2(n62), .B1(i_data_bus[32]), .B2(n89), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n62), .B1(i_data_bus[33]), .B2(n89), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n62), .B1(i_data_bus[34]), .B2(n89), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n62), .B1(i_data_bus[35]), .B2(n89), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n62), .B1(i_data_bus[36]), .B2(n89), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n62), .B1(i_data_bus[37]), .B2(n89), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n90), .B1(i_data_bus[38]), .B2(n89), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n75), .B1(i_data_bus[39]), .B2(n89), 
        .ZN(N326) );
  INVD2BWP30P140 U134 ( .I(n77), .ZN(n75) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n90), .B1(i_data_bus[63]), .B2(n89), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n75), .B1(i_data_bus[62]), .B2(n89), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n90), .B1(i_data_bus[61]), .B2(n89), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n75), .B1(i_data_bus[60]), .B2(n89), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n90), .B1(i_data_bus[59]), .B2(n89), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n75), .B1(i_data_bus[58]), .B2(n89), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n90), .B1(i_data_bus[57]), .B2(n89), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n75), .B1(i_data_bus[56]), .B2(n89), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n90), .B1(i_data_bus[55]), .B2(n89), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n75), .B1(i_data_bus[54]), .B2(n89), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n90), .B1(i_data_bus[53]), .B2(n89), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U146 ( .A1(n76), .A2(n75), .B1(i_data_bus[52]), .B2(n89), 
        .ZN(N339) );
  INVD2BWP30P140 U147 ( .I(n77), .ZN(n90) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n90), .B1(i_data_bus[51]), .B2(n89), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n75), .B1(i_data_bus[50]), .B2(n89), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n90), .B1(i_data_bus[49]), .B2(n89), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n75), .B1(i_data_bus[48]), .B2(n89), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n90), .B1(i_data_bus[47]), .B2(n89), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n75), .B1(i_data_bus[46]), .B2(n89), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n90), .B1(i_data_bus[45]), .B2(n89), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n75), .B1(i_data_bus[44]), .B2(n89), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n90), .B1(i_data_bus[43]), .B2(n89), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n75), .B1(i_data_bus[42]), .B2(n89), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n90), .B1(i_data_bus[41]), .B2(n89), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U159 ( .A1(n91), .A2(n75), .B1(i_data_bus[40]), .B2(n89), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_12 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n18), .Z(n89) );
  CKND2D3BWP30P140 U4 ( .A1(n5), .A2(n4), .ZN(n47) );
  NR2D1BWP30P140 U5 ( .A1(n49), .A2(i_cmd[1]), .ZN(n53) );
  NR2D1BWP30P140 U6 ( .A1(n49), .A2(n3), .ZN(n4) );
  ND2OPTIBD1BWP30P140 U7 ( .A1(n17), .A2(n3), .ZN(n2) );
  ND2D1BWP30P140 U8 ( .A1(n1), .A2(i_en), .ZN(n49) );
  INVD1BWP30P140 U9 ( .I(n47), .ZN(n6) );
  INVD1BWP30P140 U10 ( .I(n75), .ZN(n62) );
  INVD1BWP30P140 U11 ( .I(n89), .ZN(n19) );
  INVD1BWP30P140 U12 ( .I(n2), .ZN(n11) );
  INVD1BWP30P140 U13 ( .I(rst), .ZN(n1) );
  INVD2BWP30P140 U14 ( .I(i_valid[1]), .ZN(n50) );
  INVD2BWP30P140 U15 ( .I(i_cmd[0]), .ZN(n3) );
  INR2D2BWP30P140 U16 ( .A1(i_valid[0]), .B1(n49), .ZN(n17) );
  INVD2BWP30P140 U17 ( .I(n11), .ZN(n48) );
  OAI31D1BWP30P140 U18 ( .A1(n49), .A2(n50), .A3(n3), .B(n48), .ZN(N353) );
  INVD1BWP30P140 U19 ( .I(i_data_bus[0]), .ZN(n55) );
  INVD1BWP30P140 U20 ( .I(i_valid[0]), .ZN(n51) );
  MUX2NOPTD2BWP30P140 U21 ( .I0(n51), .I1(n50), .S(i_cmd[1]), .ZN(n5) );
  INVD2BWP30P140 U22 ( .I(n6), .ZN(n16) );
  INVD1BWP30P140 U23 ( .I(i_data_bus[32]), .ZN(n7) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n55), .B1(n16), .B2(n7), .ZN(N287) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[1]), .ZN(n56) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[33]), .ZN(n8) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n56), .B1(n16), .B2(n8), .ZN(N288) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[2]), .ZN(n57) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[34]), .ZN(n9) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n57), .B1(n16), .B2(n9), .ZN(N289) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[3]), .ZN(n58) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[35]), .ZN(n10) );
  OAI22D1BWP30P140 U33 ( .A1(n32), .A2(n58), .B1(n16), .B2(n10), .ZN(N290) );
  INVD2BWP30P140 U34 ( .I(n11), .ZN(n32) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[36]), .ZN(n12) );
  OAI22D1BWP30P140 U37 ( .A1(n32), .A2(n59), .B1(n16), .B2(n12), .ZN(N291) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[5]), .ZN(n60) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[37]), .ZN(n13) );
  OAI22D1BWP30P140 U40 ( .A1(n32), .A2(n60), .B1(n16), .B2(n13), .ZN(N292) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[6]), .ZN(n61) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[38]), .ZN(n14) );
  OAI22D1BWP30P140 U43 ( .A1(n32), .A2(n61), .B1(n16), .B2(n14), .ZN(N293) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[7]), .ZN(n63) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[39]), .ZN(n15) );
  OAI22D1BWP30P140 U46 ( .A1(n32), .A2(n63), .B1(n16), .B2(n15), .ZN(N294) );
  INVD1BWP30P140 U47 ( .I(n17), .ZN(n20) );
  INVD1BWP30P140 U48 ( .I(n49), .ZN(n18) );
  OAI21D1BWP30P140 U49 ( .A1(n20), .A2(i_cmd[1]), .B(n19), .ZN(N354) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[8]), .ZN(n74) );
  BUFFD4BWP30P140 U51 ( .I(n47), .Z(n44) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[40]), .ZN(n21) );
  OAI22D1BWP30P140 U53 ( .A1(n32), .A2(n74), .B1(n44), .B2(n21), .ZN(N295) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[9]), .ZN(n73) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[41]), .ZN(n22) );
  OAI22D1BWP30P140 U56 ( .A1(n32), .A2(n73), .B1(n44), .B2(n22), .ZN(N296) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[10]), .ZN(n72) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[42]), .ZN(n23) );
  OAI22D1BWP30P140 U59 ( .A1(n32), .A2(n72), .B1(n44), .B2(n23), .ZN(N297) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[11]), .ZN(n71) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[43]), .ZN(n24) );
  OAI22D1BWP30P140 U62 ( .A1(n32), .A2(n71), .B1(n44), .B2(n24), .ZN(N298) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[12]), .ZN(n70) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[44]), .ZN(n25) );
  OAI22D1BWP30P140 U65 ( .A1(n32), .A2(n70), .B1(n44), .B2(n25), .ZN(N299) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[13]), .ZN(n69) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[45]), .ZN(n26) );
  OAI22D1BWP30P140 U68 ( .A1(n32), .A2(n69), .B1(n44), .B2(n26), .ZN(N300) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[14]), .ZN(n68) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[46]), .ZN(n27) );
  OAI22D1BWP30P140 U71 ( .A1(n32), .A2(n68), .B1(n44), .B2(n27), .ZN(N301) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[15]), .ZN(n67) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[47]), .ZN(n28) );
  OAI22D1BWP30P140 U74 ( .A1(n32), .A2(n67), .B1(n44), .B2(n28), .ZN(N302) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[16]), .ZN(n66) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[48]), .ZN(n29) );
  OAI22D1BWP30P140 U77 ( .A1(n32), .A2(n66), .B1(n44), .B2(n29), .ZN(N303) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[17]), .ZN(n65) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[49]), .ZN(n30) );
  OAI22D1BWP30P140 U80 ( .A1(n32), .A2(n65), .B1(n44), .B2(n30), .ZN(N304) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[18]), .ZN(n64) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[50]), .ZN(n31) );
  OAI22D1BWP30P140 U83 ( .A1(n32), .A2(n64), .B1(n44), .B2(n31), .ZN(N305) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[19]), .ZN(n91) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[51]), .ZN(n33) );
  OAI22D1BWP30P140 U86 ( .A1(n48), .A2(n91), .B1(n44), .B2(n33), .ZN(N306) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[20]), .ZN(n88) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[52]), .ZN(n34) );
  OAI22D1BWP30P140 U89 ( .A1(n48), .A2(n88), .B1(n44), .B2(n34), .ZN(N307) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[21]), .ZN(n86) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[53]), .ZN(n35) );
  OAI22D1BWP30P140 U92 ( .A1(n48), .A2(n86), .B1(n44), .B2(n35), .ZN(N308) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[22]), .ZN(n85) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[54]), .ZN(n36) );
  OAI22D1BWP30P140 U95 ( .A1(n48), .A2(n85), .B1(n44), .B2(n36), .ZN(N309) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[23]), .ZN(n84) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[55]), .ZN(n37) );
  OAI22D1BWP30P140 U98 ( .A1(n48), .A2(n84), .B1(n44), .B2(n37), .ZN(N310) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[56]), .ZN(n38) );
  OAI22D1BWP30P140 U101 ( .A1(n48), .A2(n83), .B1(n44), .B2(n38), .ZN(N311) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[25]), .ZN(n82) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[57]), .ZN(n39) );
  OAI22D1BWP30P140 U104 ( .A1(n48), .A2(n82), .B1(n44), .B2(n39), .ZN(N312) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[26]), .ZN(n81) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[58]), .ZN(n40) );
  OAI22D1BWP30P140 U107 ( .A1(n48), .A2(n81), .B1(n44), .B2(n40), .ZN(N313) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[27]), .ZN(n80) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[59]), .ZN(n41) );
  OAI22D1BWP30P140 U110 ( .A1(n48), .A2(n80), .B1(n44), .B2(n41), .ZN(N314) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[28]), .ZN(n79) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[60]), .ZN(n42) );
  OAI22D1BWP30P140 U113 ( .A1(n48), .A2(n79), .B1(n44), .B2(n42), .ZN(N315) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[29]), .ZN(n78) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[61]), .ZN(n43) );
  OAI22D1BWP30P140 U116 ( .A1(n48), .A2(n78), .B1(n44), .B2(n43), .ZN(N316) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[30]), .ZN(n77) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[62]), .ZN(n45) );
  OAI22D1BWP30P140 U119 ( .A1(n48), .A2(n77), .B1(n47), .B2(n45), .ZN(N317) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[31]), .ZN(n76) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[63]), .ZN(n46) );
  OAI22D1BWP30P140 U122 ( .A1(n48), .A2(n76), .B1(n47), .B2(n46), .ZN(N318) );
  MUX2NUD1BWP30P140 U123 ( .I0(n51), .I1(n50), .S(i_cmd[0]), .ZN(n52) );
  ND2OPTIBD1BWP30P140 U124 ( .A1(n53), .A2(n52), .ZN(n54) );
  INVD2BWP30P140 U125 ( .I(n54), .ZN(n75) );
  MOAI22D1BWP30P140 U126 ( .A1(n55), .A2(n62), .B1(i_data_bus[32]), .B2(n89), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n62), .B1(i_data_bus[33]), .B2(n89), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n62), .B1(i_data_bus[34]), .B2(n89), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n62), .B1(i_data_bus[35]), .B2(n89), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n62), .B1(i_data_bus[36]), .B2(n89), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n62), .B1(i_data_bus[37]), .B2(n89), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n87), .B1(i_data_bus[38]), .B2(n89), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n90), .B1(i_data_bus[39]), .B2(n89), 
        .ZN(N326) );
  INVD2BWP30P140 U134 ( .I(n75), .ZN(n90) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n87), .B1(i_data_bus[50]), .B2(n89), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n90), .B1(i_data_bus[49]), .B2(n89), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n87), .B1(i_data_bus[48]), .B2(n89), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n90), .B1(i_data_bus[47]), .B2(n89), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n87), .B1(i_data_bus[46]), .B2(n89), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n90), .B1(i_data_bus[45]), .B2(n89), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n87), .B1(i_data_bus[44]), .B2(n89), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n90), .B1(i_data_bus[43]), .B2(n89), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n87), .B1(i_data_bus[42]), .B2(n89), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n90), .B1(i_data_bus[41]), .B2(n89), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n87), .B1(i_data_bus[40]), .B2(n89), 
        .ZN(N327) );
  INVD2BWP30P140 U146 ( .I(n75), .ZN(n87) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n87), .B1(i_data_bus[63]), .B2(n89), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n90), .B1(i_data_bus[62]), .B2(n89), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n87), .B1(i_data_bus[61]), .B2(n89), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n90), .B1(i_data_bus[60]), .B2(n89), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n87), .B1(i_data_bus[59]), .B2(n89), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n90), .B1(i_data_bus[58]), .B2(n89), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n87), .B1(i_data_bus[57]), .B2(n89), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n90), .B1(i_data_bus[56]), .B2(n89), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n87), .B1(i_data_bus[55]), .B2(n89), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U156 ( .A1(n85), .A2(n90), .B1(i_data_bus[54]), .B2(n89), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U157 ( .A1(n86), .A2(n87), .B1(i_data_bus[53]), .B2(n89), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n90), .B1(i_data_bus[52]), .B2(n89), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U159 ( .A1(n91), .A2(n90), .B1(i_data_bus[51]), .B2(n89), 
        .ZN(N338) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_13 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n18), .Z(n89) );
  CKND2D3BWP30P140 U4 ( .A1(n5), .A2(n4), .ZN(n47) );
  NR2D1BWP30P140 U5 ( .A1(n49), .A2(i_cmd[1]), .ZN(n53) );
  INVD1BWP30P140 U6 ( .I(i_cmd[0]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U7 ( .A1(n17), .A2(n3), .ZN(n2) );
  ND2D1BWP30P140 U8 ( .A1(n1), .A2(i_en), .ZN(n49) );
  INVD1BWP30P140 U9 ( .I(n47), .ZN(n6) );
  INVD1BWP30P140 U10 ( .I(n77), .ZN(n62) );
  INVD1BWP30P140 U11 ( .I(n89), .ZN(n19) );
  INVD1BWP30P140 U12 ( .I(n2), .ZN(n11) );
  INVD1BWP30P140 U13 ( .I(rst), .ZN(n1) );
  INVD2BWP30P140 U14 ( .I(i_valid[1]), .ZN(n50) );
  INR2D2BWP30P140 U15 ( .A1(i_valid[0]), .B1(n49), .ZN(n17) );
  INVD2BWP30P140 U16 ( .I(n11), .ZN(n48) );
  OAI31D1BWP30P140 U17 ( .A1(n49), .A2(n50), .A3(n3), .B(n48), .ZN(N353) );
  INVD1BWP30P140 U18 ( .I(i_data_bus[0]), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(i_valid[0]), .ZN(n51) );
  MUX2NOPTD2BWP30P140 U20 ( .I0(n51), .I1(n50), .S(i_cmd[1]), .ZN(n5) );
  NR2OPTPAD1BWP30P140 U21 ( .A1(n49), .A2(n3), .ZN(n4) );
  INVD2BWP30P140 U22 ( .I(n6), .ZN(n16) );
  INVD1BWP30P140 U23 ( .I(i_data_bus[32]), .ZN(n7) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n63), .B1(n16), .B2(n7), .ZN(N287) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[1]), .ZN(n61) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[33]), .ZN(n8) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n61), .B1(n16), .B2(n8), .ZN(N288) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[34]), .ZN(n9) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n60), .B1(n16), .B2(n9), .ZN(N289) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[3]), .ZN(n59) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[35]), .ZN(n10) );
  OAI22D1BWP30P140 U33 ( .A1(n32), .A2(n59), .B1(n16), .B2(n10), .ZN(N290) );
  INVD2BWP30P140 U34 ( .I(n11), .ZN(n32) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[4]), .ZN(n58) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[36]), .ZN(n12) );
  OAI22D1BWP30P140 U37 ( .A1(n32), .A2(n58), .B1(n16), .B2(n12), .ZN(N291) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[5]), .ZN(n57) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[37]), .ZN(n13) );
  OAI22D1BWP30P140 U40 ( .A1(n32), .A2(n57), .B1(n16), .B2(n13), .ZN(N292) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[6]), .ZN(n56) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[38]), .ZN(n14) );
  OAI22D1BWP30P140 U43 ( .A1(n32), .A2(n56), .B1(n16), .B2(n14), .ZN(N293) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[7]), .ZN(n55) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[39]), .ZN(n15) );
  OAI22D1BWP30P140 U46 ( .A1(n32), .A2(n55), .B1(n16), .B2(n15), .ZN(N294) );
  INVD1BWP30P140 U47 ( .I(n17), .ZN(n20) );
  INVD1BWP30P140 U48 ( .I(n49), .ZN(n18) );
  OAI21D1BWP30P140 U49 ( .A1(n20), .A2(i_cmd[1]), .B(n19), .ZN(N354) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[8]), .ZN(n91) );
  BUFFD4BWP30P140 U51 ( .I(n47), .Z(n44) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[40]), .ZN(n21) );
  OAI22D1BWP30P140 U53 ( .A1(n32), .A2(n91), .B1(n44), .B2(n21), .ZN(N295) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[9]), .ZN(n88) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[41]), .ZN(n22) );
  OAI22D1BWP30P140 U56 ( .A1(n32), .A2(n88), .B1(n44), .B2(n22), .ZN(N296) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[10]), .ZN(n87) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[42]), .ZN(n23) );
  OAI22D1BWP30P140 U59 ( .A1(n32), .A2(n87), .B1(n44), .B2(n23), .ZN(N297) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[11]), .ZN(n86) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[43]), .ZN(n24) );
  OAI22D1BWP30P140 U62 ( .A1(n32), .A2(n86), .B1(n44), .B2(n24), .ZN(N298) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[12]), .ZN(n85) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[44]), .ZN(n25) );
  OAI22D1BWP30P140 U65 ( .A1(n32), .A2(n85), .B1(n44), .B2(n25), .ZN(N299) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[13]), .ZN(n84) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[45]), .ZN(n26) );
  OAI22D1BWP30P140 U68 ( .A1(n32), .A2(n84), .B1(n44), .B2(n26), .ZN(N300) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[14]), .ZN(n83) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[46]), .ZN(n27) );
  OAI22D1BWP30P140 U71 ( .A1(n32), .A2(n83), .B1(n44), .B2(n27), .ZN(N301) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[15]), .ZN(n82) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[47]), .ZN(n28) );
  OAI22D1BWP30P140 U74 ( .A1(n32), .A2(n82), .B1(n44), .B2(n28), .ZN(N302) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[16]), .ZN(n81) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[48]), .ZN(n29) );
  OAI22D1BWP30P140 U77 ( .A1(n32), .A2(n81), .B1(n44), .B2(n29), .ZN(N303) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[17]), .ZN(n80) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[49]), .ZN(n30) );
  OAI22D1BWP30P140 U80 ( .A1(n32), .A2(n80), .B1(n44), .B2(n30), .ZN(N304) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[18]), .ZN(n79) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[50]), .ZN(n31) );
  OAI22D1BWP30P140 U83 ( .A1(n32), .A2(n79), .B1(n44), .B2(n31), .ZN(N305) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[51]), .ZN(n33) );
  OAI22D1BWP30P140 U86 ( .A1(n48), .A2(n78), .B1(n44), .B2(n33), .ZN(N306) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[20]), .ZN(n76) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[52]), .ZN(n34) );
  OAI22D1BWP30P140 U89 ( .A1(n48), .A2(n76), .B1(n44), .B2(n34), .ZN(N307) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[21]), .ZN(n74) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[53]), .ZN(n35) );
  OAI22D1BWP30P140 U92 ( .A1(n48), .A2(n74), .B1(n44), .B2(n35), .ZN(N308) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[22]), .ZN(n73) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[54]), .ZN(n36) );
  OAI22D1BWP30P140 U95 ( .A1(n48), .A2(n73), .B1(n44), .B2(n36), .ZN(N309) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[23]), .ZN(n72) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[55]), .ZN(n37) );
  OAI22D1BWP30P140 U98 ( .A1(n48), .A2(n72), .B1(n44), .B2(n37), .ZN(N310) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[24]), .ZN(n71) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[56]), .ZN(n38) );
  OAI22D1BWP30P140 U101 ( .A1(n48), .A2(n71), .B1(n44), .B2(n38), .ZN(N311) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[25]), .ZN(n70) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[57]), .ZN(n39) );
  OAI22D1BWP30P140 U104 ( .A1(n48), .A2(n70), .B1(n44), .B2(n39), .ZN(N312) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[26]), .ZN(n69) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[58]), .ZN(n40) );
  OAI22D1BWP30P140 U107 ( .A1(n48), .A2(n69), .B1(n44), .B2(n40), .ZN(N313) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[27]), .ZN(n68) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[59]), .ZN(n41) );
  OAI22D1BWP30P140 U110 ( .A1(n48), .A2(n68), .B1(n44), .B2(n41), .ZN(N314) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[28]), .ZN(n67) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[60]), .ZN(n42) );
  OAI22D1BWP30P140 U113 ( .A1(n48), .A2(n67), .B1(n44), .B2(n42), .ZN(N315) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[29]), .ZN(n66) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[61]), .ZN(n43) );
  OAI22D1BWP30P140 U116 ( .A1(n48), .A2(n66), .B1(n44), .B2(n43), .ZN(N316) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[30]), .ZN(n65) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[62]), .ZN(n45) );
  OAI22D1BWP30P140 U119 ( .A1(n48), .A2(n65), .B1(n47), .B2(n45), .ZN(N317) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[31]), .ZN(n64) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[63]), .ZN(n46) );
  OAI22D1BWP30P140 U122 ( .A1(n48), .A2(n64), .B1(n47), .B2(n46), .ZN(N318) );
  MUX2NUD1BWP30P140 U123 ( .I0(n51), .I1(n50), .S(i_cmd[0]), .ZN(n52) );
  ND2OPTIBD1BWP30P140 U124 ( .A1(n53), .A2(n52), .ZN(n54) );
  INVD2BWP30P140 U125 ( .I(n54), .ZN(n77) );
  MOAI22D1BWP30P140 U126 ( .A1(n55), .A2(n62), .B1(i_data_bus[39]), .B2(n89), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n62), .B1(i_data_bus[38]), .B2(n89), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n62), .B1(i_data_bus[37]), .B2(n89), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n62), .B1(i_data_bus[36]), .B2(n89), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n62), .B1(i_data_bus[35]), .B2(n89), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n62), .B1(i_data_bus[34]), .B2(n89), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n90), .B1(i_data_bus[33]), .B2(n89), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n75), .B1(i_data_bus[32]), .B2(n89), 
        .ZN(N319) );
  INVD2BWP30P140 U134 ( .I(n77), .ZN(n75) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n90), .B1(i_data_bus[63]), .B2(n89), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n75), .B1(i_data_bus[62]), .B2(n89), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n90), .B1(i_data_bus[61]), .B2(n89), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n75), .B1(i_data_bus[60]), .B2(n89), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n90), .B1(i_data_bus[59]), .B2(n89), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n75), .B1(i_data_bus[58]), .B2(n89), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n90), .B1(i_data_bus[57]), .B2(n89), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n75), .B1(i_data_bus[56]), .B2(n89), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n90), .B1(i_data_bus[55]), .B2(n89), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n75), .B1(i_data_bus[54]), .B2(n89), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n90), .B1(i_data_bus[53]), .B2(n89), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U146 ( .A1(n76), .A2(n75), .B1(i_data_bus[52]), .B2(n89), 
        .ZN(N339) );
  INVD2BWP30P140 U147 ( .I(n77), .ZN(n90) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n90), .B1(i_data_bus[51]), .B2(n89), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n75), .B1(i_data_bus[50]), .B2(n89), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n90), .B1(i_data_bus[49]), .B2(n89), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n75), .B1(i_data_bus[48]), .B2(n89), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n90), .B1(i_data_bus[47]), .B2(n89), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n75), .B1(i_data_bus[46]), .B2(n89), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n90), .B1(i_data_bus[45]), .B2(n89), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n75), .B1(i_data_bus[44]), .B2(n89), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n90), .B1(i_data_bus[43]), .B2(n89), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n75), .B1(i_data_bus[42]), .B2(n89), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n90), .B1(i_data_bus[41]), .B2(n89), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U159 ( .A1(n91), .A2(n75), .B1(i_data_bus[40]), .B2(n89), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_14 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n18), .Z(n89) );
  CKND2D3BWP30P140 U4 ( .A1(n5), .A2(n4), .ZN(n47) );
  NR2D1BWP30P140 U5 ( .A1(n49), .A2(i_cmd[1]), .ZN(n53) );
  INVD1BWP30P140 U6 ( .I(i_cmd[0]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U7 ( .A1(n17), .A2(n3), .ZN(n2) );
  ND2D1BWP30P140 U8 ( .A1(n1), .A2(i_en), .ZN(n49) );
  INVD1BWP30P140 U9 ( .I(n47), .ZN(n6) );
  INVD1BWP30P140 U10 ( .I(n77), .ZN(n62) );
  INVD1BWP30P140 U11 ( .I(n89), .ZN(n19) );
  INVD1BWP30P140 U12 ( .I(n2), .ZN(n11) );
  INVD1BWP30P140 U13 ( .I(rst), .ZN(n1) );
  INVD2BWP30P140 U14 ( .I(i_valid[1]), .ZN(n50) );
  INR2D2BWP30P140 U15 ( .A1(i_valid[0]), .B1(n49), .ZN(n17) );
  INVD2BWP30P140 U16 ( .I(n11), .ZN(n48) );
  OAI31D1BWP30P140 U17 ( .A1(n49), .A2(n50), .A3(n3), .B(n48), .ZN(N353) );
  INVD2BWP30P140 U18 ( .I(n11), .ZN(n32) );
  INVD1BWP30P140 U19 ( .I(i_data_bus[4]), .ZN(n63) );
  INVD1BWP30P140 U20 ( .I(i_valid[0]), .ZN(n51) );
  MUX2NOPTD2BWP30P140 U21 ( .I0(n51), .I1(n50), .S(i_cmd[1]), .ZN(n5) );
  NR2OPTPAD1BWP30P140 U22 ( .A1(n49), .A2(n3), .ZN(n4) );
  INVD2BWP30P140 U23 ( .I(n6), .ZN(n16) );
  INVD1BWP30P140 U24 ( .I(i_data_bus[36]), .ZN(n7) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n63), .B1(n16), .B2(n7), .ZN(N291) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[5]), .ZN(n55) );
  INVD1BWP30P140 U27 ( .I(i_data_bus[37]), .ZN(n8) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n55), .B1(n16), .B2(n8), .ZN(N292) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[38]), .ZN(n9) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n58), .B1(n16), .B2(n9), .ZN(N293) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[39]), .ZN(n10) );
  OAI22D1BWP30P140 U34 ( .A1(n32), .A2(n57), .B1(n16), .B2(n10), .ZN(N294) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[2]), .ZN(n56) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[34]), .ZN(n12) );
  OAI22D1BWP30P140 U37 ( .A1(n32), .A2(n56), .B1(n16), .B2(n12), .ZN(N289) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[35]), .ZN(n13) );
  OAI22D1BWP30P140 U40 ( .A1(n32), .A2(n61), .B1(n16), .B2(n13), .ZN(N290) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[0]), .ZN(n59) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[32]), .ZN(n14) );
  OAI22D1BWP30P140 U43 ( .A1(n32), .A2(n59), .B1(n16), .B2(n14), .ZN(N287) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[1]), .ZN(n60) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[33]), .ZN(n15) );
  OAI22D1BWP30P140 U46 ( .A1(n32), .A2(n60), .B1(n16), .B2(n15), .ZN(N288) );
  INVD1BWP30P140 U47 ( .I(n17), .ZN(n20) );
  INVD1BWP30P140 U48 ( .I(n49), .ZN(n18) );
  OAI21D1BWP30P140 U49 ( .A1(n20), .A2(i_cmd[1]), .B(n19), .ZN(N354) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[8]), .ZN(n91) );
  BUFFD4BWP30P140 U51 ( .I(n47), .Z(n44) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[40]), .ZN(n21) );
  OAI22D1BWP30P140 U53 ( .A1(n32), .A2(n91), .B1(n44), .B2(n21), .ZN(N295) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[9]), .ZN(n88) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[41]), .ZN(n22) );
  OAI22D1BWP30P140 U56 ( .A1(n32), .A2(n88), .B1(n44), .B2(n22), .ZN(N296) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[10]), .ZN(n87) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[42]), .ZN(n23) );
  OAI22D1BWP30P140 U59 ( .A1(n32), .A2(n87), .B1(n44), .B2(n23), .ZN(N297) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[11]), .ZN(n86) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[43]), .ZN(n24) );
  OAI22D1BWP30P140 U62 ( .A1(n32), .A2(n86), .B1(n44), .B2(n24), .ZN(N298) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[12]), .ZN(n85) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[44]), .ZN(n25) );
  OAI22D1BWP30P140 U65 ( .A1(n32), .A2(n85), .B1(n44), .B2(n25), .ZN(N299) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[13]), .ZN(n84) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[45]), .ZN(n26) );
  OAI22D1BWP30P140 U68 ( .A1(n32), .A2(n84), .B1(n44), .B2(n26), .ZN(N300) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[14]), .ZN(n83) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[46]), .ZN(n27) );
  OAI22D1BWP30P140 U71 ( .A1(n32), .A2(n83), .B1(n44), .B2(n27), .ZN(N301) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[15]), .ZN(n82) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[47]), .ZN(n28) );
  OAI22D1BWP30P140 U74 ( .A1(n32), .A2(n82), .B1(n44), .B2(n28), .ZN(N302) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[16]), .ZN(n81) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[48]), .ZN(n29) );
  OAI22D1BWP30P140 U77 ( .A1(n32), .A2(n81), .B1(n44), .B2(n29), .ZN(N303) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[17]), .ZN(n80) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[49]), .ZN(n30) );
  OAI22D1BWP30P140 U80 ( .A1(n32), .A2(n80), .B1(n44), .B2(n30), .ZN(N304) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[18]), .ZN(n79) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[50]), .ZN(n31) );
  OAI22D1BWP30P140 U83 ( .A1(n32), .A2(n79), .B1(n44), .B2(n31), .ZN(N305) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[51]), .ZN(n33) );
  OAI22D1BWP30P140 U86 ( .A1(n48), .A2(n78), .B1(n44), .B2(n33), .ZN(N306) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[20]), .ZN(n76) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[52]), .ZN(n34) );
  OAI22D1BWP30P140 U89 ( .A1(n48), .A2(n76), .B1(n44), .B2(n34), .ZN(N307) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[21]), .ZN(n74) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[53]), .ZN(n35) );
  OAI22D1BWP30P140 U92 ( .A1(n48), .A2(n74), .B1(n44), .B2(n35), .ZN(N308) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[22]), .ZN(n73) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[54]), .ZN(n36) );
  OAI22D1BWP30P140 U95 ( .A1(n48), .A2(n73), .B1(n44), .B2(n36), .ZN(N309) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[23]), .ZN(n72) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[55]), .ZN(n37) );
  OAI22D1BWP30P140 U98 ( .A1(n48), .A2(n72), .B1(n44), .B2(n37), .ZN(N310) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[24]), .ZN(n71) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[56]), .ZN(n38) );
  OAI22D1BWP30P140 U101 ( .A1(n48), .A2(n71), .B1(n44), .B2(n38), .ZN(N311) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[25]), .ZN(n70) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[57]), .ZN(n39) );
  OAI22D1BWP30P140 U104 ( .A1(n48), .A2(n70), .B1(n44), .B2(n39), .ZN(N312) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[26]), .ZN(n69) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[58]), .ZN(n40) );
  OAI22D1BWP30P140 U107 ( .A1(n48), .A2(n69), .B1(n44), .B2(n40), .ZN(N313) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[27]), .ZN(n68) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[59]), .ZN(n41) );
  OAI22D1BWP30P140 U110 ( .A1(n48), .A2(n68), .B1(n44), .B2(n41), .ZN(N314) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[28]), .ZN(n67) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[60]), .ZN(n42) );
  OAI22D1BWP30P140 U113 ( .A1(n48), .A2(n67), .B1(n44), .B2(n42), .ZN(N315) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[29]), .ZN(n66) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[61]), .ZN(n43) );
  OAI22D1BWP30P140 U116 ( .A1(n48), .A2(n66), .B1(n44), .B2(n43), .ZN(N316) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[30]), .ZN(n65) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[62]), .ZN(n45) );
  OAI22D1BWP30P140 U119 ( .A1(n48), .A2(n65), .B1(n47), .B2(n45), .ZN(N317) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[31]), .ZN(n64) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[63]), .ZN(n46) );
  OAI22D1BWP30P140 U122 ( .A1(n48), .A2(n64), .B1(n47), .B2(n46), .ZN(N318) );
  MUX2NUD1BWP30P140 U123 ( .I0(n51), .I1(n50), .S(i_cmd[0]), .ZN(n52) );
  ND2OPTIBD1BWP30P140 U124 ( .A1(n53), .A2(n52), .ZN(n54) );
  INVD2BWP30P140 U125 ( .I(n54), .ZN(n77) );
  MOAI22D1BWP30P140 U126 ( .A1(n55), .A2(n62), .B1(i_data_bus[37]), .B2(n89), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n62), .B1(i_data_bus[34]), .B2(n89), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n62), .B1(i_data_bus[39]), .B2(n89), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n62), .B1(i_data_bus[38]), .B2(n89), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n62), .B1(i_data_bus[32]), .B2(n89), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n62), .B1(i_data_bus[33]), .B2(n89), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n90), .B1(i_data_bus[35]), .B2(n89), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n75), .B1(i_data_bus[36]), .B2(n89), 
        .ZN(N323) );
  INVD2BWP30P140 U134 ( .I(n77), .ZN(n75) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n90), .B1(i_data_bus[63]), .B2(n89), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n75), .B1(i_data_bus[62]), .B2(n89), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n90), .B1(i_data_bus[61]), .B2(n89), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n75), .B1(i_data_bus[60]), .B2(n89), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n90), .B1(i_data_bus[59]), .B2(n89), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n75), .B1(i_data_bus[58]), .B2(n89), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n90), .B1(i_data_bus[57]), .B2(n89), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n75), .B1(i_data_bus[56]), .B2(n89), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n90), .B1(i_data_bus[55]), .B2(n89), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n75), .B1(i_data_bus[54]), .B2(n89), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n90), .B1(i_data_bus[53]), .B2(n89), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U146 ( .A1(n76), .A2(n75), .B1(i_data_bus[52]), .B2(n89), 
        .ZN(N339) );
  INVD2BWP30P140 U147 ( .I(n77), .ZN(n90) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n90), .B1(i_data_bus[51]), .B2(n89), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n75), .B1(i_data_bus[50]), .B2(n89), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n90), .B1(i_data_bus[49]), .B2(n89), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n75), .B1(i_data_bus[48]), .B2(n89), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n90), .B1(i_data_bus[47]), .B2(n89), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n75), .B1(i_data_bus[46]), .B2(n89), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n90), .B1(i_data_bus[45]), .B2(n89), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n75), .B1(i_data_bus[44]), .B2(n89), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n90), .B1(i_data_bus[43]), .B2(n89), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n75), .B1(i_data_bus[42]), .B2(n89), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n90), .B1(i_data_bus[41]), .B2(n89), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U159 ( .A1(n91), .A2(n75), .B1(i_data_bus[40]), .B2(n89), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_15 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n18), .Z(n89) );
  CKND2D3BWP30P140 U4 ( .A1(n5), .A2(n4), .ZN(n47) );
  NR2D1BWP30P140 U5 ( .A1(n49), .A2(i_cmd[1]), .ZN(n53) );
  INVD1BWP30P140 U6 ( .I(i_cmd[0]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U7 ( .A1(n17), .A2(n3), .ZN(n2) );
  ND2D1BWP30P140 U8 ( .A1(n1), .A2(i_en), .ZN(n49) );
  INVD1BWP30P140 U9 ( .I(n47), .ZN(n6) );
  INVD1BWP30P140 U10 ( .I(n77), .ZN(n62) );
  INVD1BWP30P140 U11 ( .I(n89), .ZN(n19) );
  INVD1BWP30P140 U12 ( .I(n2), .ZN(n9) );
  INVD1BWP30P140 U13 ( .I(rst), .ZN(n1) );
  INVD2BWP30P140 U14 ( .I(i_valid[1]), .ZN(n50) );
  INR2D2BWP30P140 U15 ( .A1(i_valid[0]), .B1(n49), .ZN(n17) );
  INVD2BWP30P140 U16 ( .I(n9), .ZN(n48) );
  OAI31D1BWP30P140 U17 ( .A1(n49), .A2(n50), .A3(n3), .B(n48), .ZN(N353) );
  INVD2BWP30P140 U18 ( .I(n9), .ZN(n32) );
  INVD1BWP30P140 U19 ( .I(i_data_bus[7]), .ZN(n63) );
  INVD1BWP30P140 U20 ( .I(i_valid[0]), .ZN(n51) );
  MUX2NOPTD2BWP30P140 U21 ( .I0(n51), .I1(n50), .S(i_cmd[1]), .ZN(n5) );
  NR2OPTPAD1BWP30P140 U22 ( .A1(n49), .A2(n3), .ZN(n4) );
  INVD2BWP30P140 U23 ( .I(n6), .ZN(n16) );
  INVD1BWP30P140 U24 ( .I(i_data_bus[39]), .ZN(n7) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n63), .B1(n16), .B2(n7), .ZN(N294) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[6]), .ZN(n61) );
  INVD1BWP30P140 U27 ( .I(i_data_bus[38]), .ZN(n8) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n61), .B1(n16), .B2(n8), .ZN(N293) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[0]), .ZN(n55) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[32]), .ZN(n10) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n55), .B1(n16), .B2(n10), .ZN(N287) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[2]), .ZN(n57) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[34]), .ZN(n11) );
  OAI22D1BWP30P140 U34 ( .A1(n32), .A2(n57), .B1(n16), .B2(n11), .ZN(N289) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[3]), .ZN(n58) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[35]), .ZN(n12) );
  OAI22D1BWP30P140 U37 ( .A1(n32), .A2(n58), .B1(n16), .B2(n12), .ZN(N290) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[36]), .ZN(n13) );
  OAI22D1BWP30P140 U40 ( .A1(n32), .A2(n59), .B1(n16), .B2(n13), .ZN(N291) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[5]), .ZN(n60) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[37]), .ZN(n14) );
  OAI22D1BWP30P140 U43 ( .A1(n32), .A2(n60), .B1(n16), .B2(n14), .ZN(N292) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[1]), .ZN(n56) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[33]), .ZN(n15) );
  OAI22D1BWP30P140 U46 ( .A1(n32), .A2(n56), .B1(n16), .B2(n15), .ZN(N288) );
  INVD1BWP30P140 U47 ( .I(n17), .ZN(n20) );
  INVD1BWP30P140 U48 ( .I(n49), .ZN(n18) );
  OAI21D1BWP30P140 U49 ( .A1(n20), .A2(i_cmd[1]), .B(n19), .ZN(N354) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[8]), .ZN(n91) );
  BUFFD4BWP30P140 U51 ( .I(n47), .Z(n44) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[40]), .ZN(n21) );
  OAI22D1BWP30P140 U53 ( .A1(n32), .A2(n91), .B1(n44), .B2(n21), .ZN(N295) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[9]), .ZN(n88) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[41]), .ZN(n22) );
  OAI22D1BWP30P140 U56 ( .A1(n32), .A2(n88), .B1(n44), .B2(n22), .ZN(N296) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[10]), .ZN(n87) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[42]), .ZN(n23) );
  OAI22D1BWP30P140 U59 ( .A1(n32), .A2(n87), .B1(n44), .B2(n23), .ZN(N297) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[11]), .ZN(n86) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[43]), .ZN(n24) );
  OAI22D1BWP30P140 U62 ( .A1(n32), .A2(n86), .B1(n44), .B2(n24), .ZN(N298) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[12]), .ZN(n85) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[44]), .ZN(n25) );
  OAI22D1BWP30P140 U65 ( .A1(n32), .A2(n85), .B1(n44), .B2(n25), .ZN(N299) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[13]), .ZN(n84) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[45]), .ZN(n26) );
  OAI22D1BWP30P140 U68 ( .A1(n32), .A2(n84), .B1(n44), .B2(n26), .ZN(N300) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[14]), .ZN(n83) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[46]), .ZN(n27) );
  OAI22D1BWP30P140 U71 ( .A1(n32), .A2(n83), .B1(n44), .B2(n27), .ZN(N301) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[15]), .ZN(n82) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[47]), .ZN(n28) );
  OAI22D1BWP30P140 U74 ( .A1(n32), .A2(n82), .B1(n44), .B2(n28), .ZN(N302) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[16]), .ZN(n81) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[48]), .ZN(n29) );
  OAI22D1BWP30P140 U77 ( .A1(n32), .A2(n81), .B1(n44), .B2(n29), .ZN(N303) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[17]), .ZN(n80) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[49]), .ZN(n30) );
  OAI22D1BWP30P140 U80 ( .A1(n32), .A2(n80), .B1(n44), .B2(n30), .ZN(N304) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[18]), .ZN(n79) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[50]), .ZN(n31) );
  OAI22D1BWP30P140 U83 ( .A1(n32), .A2(n79), .B1(n44), .B2(n31), .ZN(N305) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[51]), .ZN(n33) );
  OAI22D1BWP30P140 U86 ( .A1(n48), .A2(n78), .B1(n44), .B2(n33), .ZN(N306) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[20]), .ZN(n76) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[52]), .ZN(n34) );
  OAI22D1BWP30P140 U89 ( .A1(n48), .A2(n76), .B1(n44), .B2(n34), .ZN(N307) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[21]), .ZN(n74) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[53]), .ZN(n35) );
  OAI22D1BWP30P140 U92 ( .A1(n48), .A2(n74), .B1(n44), .B2(n35), .ZN(N308) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[22]), .ZN(n73) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[54]), .ZN(n36) );
  OAI22D1BWP30P140 U95 ( .A1(n48), .A2(n73), .B1(n44), .B2(n36), .ZN(N309) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[23]), .ZN(n72) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[55]), .ZN(n37) );
  OAI22D1BWP30P140 U98 ( .A1(n48), .A2(n72), .B1(n44), .B2(n37), .ZN(N310) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[24]), .ZN(n71) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[56]), .ZN(n38) );
  OAI22D1BWP30P140 U101 ( .A1(n48), .A2(n71), .B1(n44), .B2(n38), .ZN(N311) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[25]), .ZN(n70) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[57]), .ZN(n39) );
  OAI22D1BWP30P140 U104 ( .A1(n48), .A2(n70), .B1(n44), .B2(n39), .ZN(N312) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[26]), .ZN(n69) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[58]), .ZN(n40) );
  OAI22D1BWP30P140 U107 ( .A1(n48), .A2(n69), .B1(n44), .B2(n40), .ZN(N313) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[27]), .ZN(n68) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[59]), .ZN(n41) );
  OAI22D1BWP30P140 U110 ( .A1(n48), .A2(n68), .B1(n44), .B2(n41), .ZN(N314) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[28]), .ZN(n67) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[60]), .ZN(n42) );
  OAI22D1BWP30P140 U113 ( .A1(n48), .A2(n67), .B1(n44), .B2(n42), .ZN(N315) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[29]), .ZN(n66) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[61]), .ZN(n43) );
  OAI22D1BWP30P140 U116 ( .A1(n48), .A2(n66), .B1(n44), .B2(n43), .ZN(N316) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[30]), .ZN(n65) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[62]), .ZN(n45) );
  OAI22D1BWP30P140 U119 ( .A1(n48), .A2(n65), .B1(n47), .B2(n45), .ZN(N317) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[31]), .ZN(n64) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[63]), .ZN(n46) );
  OAI22D1BWP30P140 U122 ( .A1(n48), .A2(n64), .B1(n47), .B2(n46), .ZN(N318) );
  MUX2NUD1BWP30P140 U123 ( .I0(n51), .I1(n50), .S(i_cmd[0]), .ZN(n52) );
  ND2OPTIBD1BWP30P140 U124 ( .A1(n53), .A2(n52), .ZN(n54) );
  INVD2BWP30P140 U125 ( .I(n54), .ZN(n77) );
  MOAI22D1BWP30P140 U126 ( .A1(n55), .A2(n62), .B1(i_data_bus[32]), .B2(n89), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n62), .B1(i_data_bus[33]), .B2(n89), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n62), .B1(i_data_bus[34]), .B2(n89), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n62), .B1(i_data_bus[35]), .B2(n89), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n62), .B1(i_data_bus[36]), .B2(n89), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n62), .B1(i_data_bus[37]), .B2(n89), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n90), .B1(i_data_bus[38]), .B2(n89), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n75), .B1(i_data_bus[39]), .B2(n89), 
        .ZN(N326) );
  INVD2BWP30P140 U134 ( .I(n77), .ZN(n75) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n90), .B1(i_data_bus[63]), .B2(n89), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n75), .B1(i_data_bus[62]), .B2(n89), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n90), .B1(i_data_bus[61]), .B2(n89), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n75), .B1(i_data_bus[60]), .B2(n89), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n90), .B1(i_data_bus[59]), .B2(n89), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n75), .B1(i_data_bus[58]), .B2(n89), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n90), .B1(i_data_bus[57]), .B2(n89), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n75), .B1(i_data_bus[56]), .B2(n89), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n90), .B1(i_data_bus[55]), .B2(n89), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n75), .B1(i_data_bus[54]), .B2(n89), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n90), .B1(i_data_bus[53]), .B2(n89), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U146 ( .A1(n76), .A2(n75), .B1(i_data_bus[52]), .B2(n89), 
        .ZN(N339) );
  INVD2BWP30P140 U147 ( .I(n77), .ZN(n90) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n90), .B1(i_data_bus[51]), .B2(n89), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n75), .B1(i_data_bus[50]), .B2(n89), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n90), .B1(i_data_bus[49]), .B2(n89), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n75), .B1(i_data_bus[48]), .B2(n89), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n90), .B1(i_data_bus[47]), .B2(n89), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n75), .B1(i_data_bus[46]), .B2(n89), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n90), .B1(i_data_bus[45]), .B2(n89), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n75), .B1(i_data_bus[44]), .B2(n89), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n90), .B1(i_data_bus[43]), .B2(n89), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n75), .B1(i_data_bus[42]), .B2(n89), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n90), .B1(i_data_bus[41]), .B2(n89), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U159 ( .A1(n91), .A2(n75), .B1(i_data_bus[40]), .B2(n89), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_16 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n18), .Z(n89) );
  CKND2D3BWP30P140 U4 ( .A1(n5), .A2(n4), .ZN(n47) );
  NR2D1BWP30P140 U5 ( .A1(n49), .A2(i_cmd[1]), .ZN(n53) );
  INVD1BWP30P140 U6 ( .I(i_cmd[0]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U7 ( .A1(n17), .A2(n3), .ZN(n2) );
  ND2D1BWP30P140 U8 ( .A1(n1), .A2(i_en), .ZN(n49) );
  INVD1BWP30P140 U9 ( .I(n47), .ZN(n6) );
  INVD1BWP30P140 U10 ( .I(n69), .ZN(n62) );
  INVD1BWP30P140 U11 ( .I(n89), .ZN(n19) );
  INVD1BWP30P140 U12 ( .I(n2), .ZN(n11) );
  INVD1BWP30P140 U13 ( .I(rst), .ZN(n1) );
  INVD2BWP30P140 U14 ( .I(i_valid[1]), .ZN(n50) );
  INR2D2BWP30P140 U15 ( .A1(i_valid[0]), .B1(n49), .ZN(n17) );
  INVD2BWP30P140 U16 ( .I(n11), .ZN(n45) );
  OAI31D1BWP30P140 U17 ( .A1(n49), .A2(n50), .A3(n3), .B(n45), .ZN(N353) );
  INVD1BWP30P140 U18 ( .I(i_data_bus[0]), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(i_valid[0]), .ZN(n51) );
  MUX2NOPTD2BWP30P140 U20 ( .I0(n51), .I1(n50), .S(i_cmd[1]), .ZN(n5) );
  NR2OPTPAD1BWP30P140 U21 ( .A1(n49), .A2(n3), .ZN(n4) );
  INVD2BWP30P140 U22 ( .I(n6), .ZN(n16) );
  INVD1BWP30P140 U23 ( .I(i_data_bus[32]), .ZN(n7) );
  OAI22D1BWP30P140 U24 ( .A1(n48), .A2(n63), .B1(n16), .B2(n7), .ZN(N287) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[1]), .ZN(n61) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[33]), .ZN(n8) );
  OAI22D1BWP30P140 U27 ( .A1(n48), .A2(n61), .B1(n16), .B2(n8), .ZN(N288) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[34]), .ZN(n9) );
  OAI22D1BWP30P140 U30 ( .A1(n48), .A2(n60), .B1(n16), .B2(n9), .ZN(N289) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[3]), .ZN(n59) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[35]), .ZN(n10) );
  OAI22D1BWP30P140 U33 ( .A1(n48), .A2(n59), .B1(n16), .B2(n10), .ZN(N290) );
  INVD2BWP30P140 U34 ( .I(n11), .ZN(n48) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[4]), .ZN(n58) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[36]), .ZN(n12) );
  OAI22D1BWP30P140 U37 ( .A1(n48), .A2(n58), .B1(n16), .B2(n12), .ZN(N291) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[5]), .ZN(n57) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[37]), .ZN(n13) );
  OAI22D1BWP30P140 U40 ( .A1(n48), .A2(n57), .B1(n16), .B2(n13), .ZN(N292) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[6]), .ZN(n56) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[38]), .ZN(n14) );
  OAI22D1BWP30P140 U43 ( .A1(n48), .A2(n56), .B1(n16), .B2(n14), .ZN(N293) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[7]), .ZN(n55) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[39]), .ZN(n15) );
  OAI22D1BWP30P140 U46 ( .A1(n48), .A2(n55), .B1(n16), .B2(n15), .ZN(N294) );
  INVD1BWP30P140 U47 ( .I(n17), .ZN(n20) );
  INVD1BWP30P140 U48 ( .I(n49), .ZN(n18) );
  OAI21D1BWP30P140 U49 ( .A1(n20), .A2(i_cmd[1]), .B(n19), .ZN(N354) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n67) );
  BUFFD4BWP30P140 U51 ( .I(n47), .Z(n44) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[41]), .ZN(n21) );
  OAI22D1BWP30P140 U53 ( .A1(n48), .A2(n67), .B1(n44), .B2(n21), .ZN(N296) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[10]), .ZN(n66) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[42]), .ZN(n22) );
  OAI22D1BWP30P140 U56 ( .A1(n48), .A2(n66), .B1(n44), .B2(n22), .ZN(N297) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[11]), .ZN(n65) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[43]), .ZN(n23) );
  OAI22D1BWP30P140 U59 ( .A1(n48), .A2(n65), .B1(n44), .B2(n23), .ZN(N298) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[12]), .ZN(n64) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[44]), .ZN(n24) );
  OAI22D1BWP30P140 U62 ( .A1(n48), .A2(n64), .B1(n44), .B2(n24), .ZN(N299) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[13]), .ZN(n91) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[45]), .ZN(n25) );
  OAI22D1BWP30P140 U65 ( .A1(n48), .A2(n91), .B1(n44), .B2(n25), .ZN(N300) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[14]), .ZN(n88) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[46]), .ZN(n26) );
  OAI22D1BWP30P140 U68 ( .A1(n48), .A2(n88), .B1(n44), .B2(n26), .ZN(N301) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[15]), .ZN(n87) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[47]), .ZN(n27) );
  OAI22D1BWP30P140 U71 ( .A1(n48), .A2(n87), .B1(n44), .B2(n27), .ZN(N302) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[16]), .ZN(n86) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[48]), .ZN(n28) );
  OAI22D1BWP30P140 U74 ( .A1(n48), .A2(n86), .B1(n44), .B2(n28), .ZN(N303) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[17]), .ZN(n85) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[49]), .ZN(n29) );
  OAI22D1BWP30P140 U77 ( .A1(n48), .A2(n85), .B1(n44), .B2(n29), .ZN(N304) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[18]), .ZN(n84) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[50]), .ZN(n30) );
  OAI22D1BWP30P140 U80 ( .A1(n48), .A2(n84), .B1(n44), .B2(n30), .ZN(N305) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[19]), .ZN(n83) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[51]), .ZN(n31) );
  OAI22D1BWP30P140 U83 ( .A1(n45), .A2(n83), .B1(n47), .B2(n31), .ZN(N306) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[20]), .ZN(n82) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[52]), .ZN(n32) );
  OAI22D1BWP30P140 U86 ( .A1(n45), .A2(n82), .B1(n44), .B2(n32), .ZN(N307) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[53]), .ZN(n33) );
  OAI22D1BWP30P140 U89 ( .A1(n45), .A2(n80), .B1(n44), .B2(n33), .ZN(N308) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[22]), .ZN(n79) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[54]), .ZN(n34) );
  OAI22D1BWP30P140 U92 ( .A1(n45), .A2(n79), .B1(n44), .B2(n34), .ZN(N309) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[23]), .ZN(n78) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[55]), .ZN(n35) );
  OAI22D1BWP30P140 U95 ( .A1(n45), .A2(n78), .B1(n44), .B2(n35), .ZN(N310) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[24]), .ZN(n77) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[56]), .ZN(n36) );
  OAI22D1BWP30P140 U98 ( .A1(n45), .A2(n77), .B1(n44), .B2(n36), .ZN(N311) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[25]), .ZN(n76) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[57]), .ZN(n37) );
  OAI22D1BWP30P140 U101 ( .A1(n45), .A2(n76), .B1(n44), .B2(n37), .ZN(N312) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[26]), .ZN(n75) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[58]), .ZN(n38) );
  OAI22D1BWP30P140 U104 ( .A1(n45), .A2(n75), .B1(n44), .B2(n38), .ZN(N313) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[27]), .ZN(n74) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[59]), .ZN(n39) );
  OAI22D1BWP30P140 U107 ( .A1(n45), .A2(n74), .B1(n44), .B2(n39), .ZN(N314) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[28]), .ZN(n73) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[60]), .ZN(n40) );
  OAI22D1BWP30P140 U110 ( .A1(n45), .A2(n73), .B1(n44), .B2(n40), .ZN(N315) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[29]), .ZN(n72) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[61]), .ZN(n41) );
  OAI22D1BWP30P140 U113 ( .A1(n45), .A2(n72), .B1(n44), .B2(n41), .ZN(N316) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[30]), .ZN(n71) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[62]), .ZN(n42) );
  OAI22D1BWP30P140 U116 ( .A1(n45), .A2(n71), .B1(n44), .B2(n42), .ZN(N317) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[31]), .ZN(n70) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[63]), .ZN(n43) );
  OAI22D1BWP30P140 U119 ( .A1(n45), .A2(n70), .B1(n44), .B2(n43), .ZN(N318) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[8]), .ZN(n68) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[40]), .ZN(n46) );
  OAI22D1BWP30P140 U122 ( .A1(n48), .A2(n68), .B1(n47), .B2(n46), .ZN(N295) );
  MUX2NUD1BWP30P140 U123 ( .I0(n51), .I1(n50), .S(i_cmd[0]), .ZN(n52) );
  ND2OPTIBD1BWP30P140 U124 ( .A1(n53), .A2(n52), .ZN(n54) );
  INVD2BWP30P140 U125 ( .I(n54), .ZN(n69) );
  MOAI22D1BWP30P140 U126 ( .A1(n55), .A2(n62), .B1(i_data_bus[39]), .B2(n89), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n62), .B1(i_data_bus[38]), .B2(n89), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n62), .B1(i_data_bus[37]), .B2(n89), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n62), .B1(i_data_bus[36]), .B2(n89), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n62), .B1(i_data_bus[35]), .B2(n89), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n62), .B1(i_data_bus[34]), .B2(n89), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n81), .B1(i_data_bus[33]), .B2(n89), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n90), .B1(i_data_bus[32]), .B2(n89), 
        .ZN(N319) );
  INVD2BWP30P140 U134 ( .I(n69), .ZN(n90) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n81), .B1(i_data_bus[44]), .B2(n89), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n90), .B1(i_data_bus[43]), .B2(n89), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n81), .B1(i_data_bus[42]), .B2(n89), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n90), .B1(i_data_bus[41]), .B2(n89), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n81), .B1(i_data_bus[40]), .B2(n89), 
        .ZN(N327) );
  INVD2BWP30P140 U140 ( .I(n69), .ZN(n81) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n81), .B1(i_data_bus[63]), .B2(n89), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n90), .B1(i_data_bus[62]), .B2(n89), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n81), .B1(i_data_bus[61]), .B2(n89), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n90), .B1(i_data_bus[60]), .B2(n89), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n81), .B1(i_data_bus[59]), .B2(n89), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n90), .B1(i_data_bus[58]), .B2(n89), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n81), .B1(i_data_bus[57]), .B2(n89), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n90), .B1(i_data_bus[56]), .B2(n89), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n81), .B1(i_data_bus[55]), .B2(n89), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n90), .B1(i_data_bus[54]), .B2(n89), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n81), .B1(i_data_bus[53]), .B2(n89), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n90), .B1(i_data_bus[52]), .B2(n89), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n90), .B1(i_data_bus[51]), .B2(n89), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n81), .B1(i_data_bus[50]), .B2(n89), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n90), .B1(i_data_bus[49]), .B2(n89), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n81), .B1(i_data_bus[48]), .B2(n89), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n90), .B1(i_data_bus[47]), .B2(n89), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n81), .B1(i_data_bus[46]), .B2(n89), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U159 ( .A1(n91), .A2(n90), .B1(i_data_bus[45]), .B2(n89), 
        .ZN(N332) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_17 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n18), .Z(n89) );
  CKND2D3BWP30P140 U4 ( .A1(n5), .A2(n4), .ZN(n47) );
  INR2D1BWP30P140 U5 ( .A1(i_valid[0]), .B1(n49), .ZN(n17) );
  INVD1BWP30P140 U6 ( .I(i_cmd[0]), .ZN(n3) );
  NR2D1BWP30P140 U7 ( .A1(n49), .A2(i_cmd[1]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U8 ( .A1(n17), .A2(n3), .ZN(n2) );
  ND2D1BWP30P140 U9 ( .A1(n1), .A2(i_en), .ZN(n49) );
  INVD1BWP30P140 U10 ( .I(n47), .ZN(n6) );
  INVD1BWP30P140 U11 ( .I(n77), .ZN(n62) );
  INVD1BWP30P140 U12 ( .I(n89), .ZN(n19) );
  INVD1BWP30P140 U13 ( .I(n2), .ZN(n11) );
  INVD1BWP30P140 U14 ( .I(rst), .ZN(n1) );
  INVD2BWP30P140 U15 ( .I(i_valid[1]), .ZN(n50) );
  INVD2BWP30P140 U16 ( .I(n11), .ZN(n48) );
  OAI31D1BWP30P140 U17 ( .A1(n49), .A2(n50), .A3(n3), .B(n48), .ZN(N353) );
  INVD1BWP30P140 U18 ( .I(i_data_bus[0]), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(i_valid[0]), .ZN(n51) );
  MUX2NOPTD2BWP30P140 U20 ( .I0(n51), .I1(n50), .S(i_cmd[1]), .ZN(n5) );
  NR2OPTPAD1BWP30P140 U21 ( .A1(n49), .A2(n3), .ZN(n4) );
  INVD2BWP30P140 U22 ( .I(n6), .ZN(n16) );
  INVD1BWP30P140 U23 ( .I(i_data_bus[32]), .ZN(n7) );
  OAI22D1BWP30P140 U24 ( .A1(n45), .A2(n63), .B1(n16), .B2(n7), .ZN(N287) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[1]), .ZN(n61) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[33]), .ZN(n8) );
  OAI22D1BWP30P140 U27 ( .A1(n48), .A2(n61), .B1(n16), .B2(n8), .ZN(N288) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[34]), .ZN(n9) );
  OAI22D1BWP30P140 U30 ( .A1(n45), .A2(n60), .B1(n16), .B2(n9), .ZN(N289) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[3]), .ZN(n59) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[35]), .ZN(n10) );
  OAI22D1BWP30P140 U33 ( .A1(n48), .A2(n59), .B1(n16), .B2(n10), .ZN(N290) );
  INVD2BWP30P140 U34 ( .I(n11), .ZN(n45) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[4]), .ZN(n55) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[36]), .ZN(n12) );
  OAI22D1BWP30P140 U37 ( .A1(n45), .A2(n55), .B1(n16), .B2(n12), .ZN(N291) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[5]), .ZN(n56) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[37]), .ZN(n13) );
  OAI22D1BWP30P140 U40 ( .A1(n45), .A2(n56), .B1(n16), .B2(n13), .ZN(N292) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[6]), .ZN(n57) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[38]), .ZN(n14) );
  OAI22D1BWP30P140 U43 ( .A1(n45), .A2(n57), .B1(n16), .B2(n14), .ZN(N293) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[7]), .ZN(n58) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[39]), .ZN(n15) );
  OAI22D1BWP30P140 U46 ( .A1(n45), .A2(n58), .B1(n16), .B2(n15), .ZN(N294) );
  INVD1BWP30P140 U47 ( .I(n17), .ZN(n20) );
  INVD1BWP30P140 U48 ( .I(n49), .ZN(n18) );
  OAI21D1BWP30P140 U49 ( .A1(n20), .A2(i_cmd[1]), .B(n19), .ZN(N354) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[8]), .ZN(n91) );
  BUFFD4BWP30P140 U51 ( .I(n47), .Z(n44) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[40]), .ZN(n21) );
  OAI22D1BWP30P140 U53 ( .A1(n45), .A2(n91), .B1(n44), .B2(n21), .ZN(N295) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[10]), .ZN(n87) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[42]), .ZN(n22) );
  OAI22D1BWP30P140 U56 ( .A1(n45), .A2(n87), .B1(n44), .B2(n22), .ZN(N297) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[11]), .ZN(n86) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[43]), .ZN(n23) );
  OAI22D1BWP30P140 U59 ( .A1(n45), .A2(n86), .B1(n44), .B2(n23), .ZN(N298) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[13]), .ZN(n84) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[45]), .ZN(n24) );
  OAI22D1BWP30P140 U62 ( .A1(n45), .A2(n84), .B1(n44), .B2(n24), .ZN(N300) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[14]), .ZN(n83) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[46]), .ZN(n25) );
  OAI22D1BWP30P140 U65 ( .A1(n45), .A2(n83), .B1(n44), .B2(n25), .ZN(N301) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[15]), .ZN(n82) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[47]), .ZN(n26) );
  OAI22D1BWP30P140 U68 ( .A1(n45), .A2(n82), .B1(n44), .B2(n26), .ZN(N302) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[16]), .ZN(n81) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[48]), .ZN(n27) );
  OAI22D1BWP30P140 U71 ( .A1(n45), .A2(n81), .B1(n44), .B2(n27), .ZN(N303) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[51]), .ZN(n28) );
  OAI22D1BWP30P140 U74 ( .A1(n48), .A2(n78), .B1(n44), .B2(n28), .ZN(N306) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[20]), .ZN(n76) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[52]), .ZN(n29) );
  OAI22D1BWP30P140 U77 ( .A1(n48), .A2(n76), .B1(n44), .B2(n29), .ZN(N307) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[9]), .ZN(n88) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[41]), .ZN(n30) );
  OAI22D1BWP30P140 U80 ( .A1(n45), .A2(n88), .B1(n44), .B2(n30), .ZN(N296) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[22]), .ZN(n73) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[54]), .ZN(n31) );
  OAI22D1BWP30P140 U83 ( .A1(n48), .A2(n73), .B1(n44), .B2(n31), .ZN(N309) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[12]), .ZN(n85) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[44]), .ZN(n32) );
  OAI22D1BWP30P140 U86 ( .A1(n45), .A2(n85), .B1(n44), .B2(n32), .ZN(N299) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[24]), .ZN(n71) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[56]), .ZN(n33) );
  OAI22D1BWP30P140 U89 ( .A1(n48), .A2(n71), .B1(n44), .B2(n33), .ZN(N311) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[25]), .ZN(n70) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[57]), .ZN(n34) );
  OAI22D1BWP30P140 U92 ( .A1(n48), .A2(n70), .B1(n44), .B2(n34), .ZN(N312) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[26]), .ZN(n69) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[58]), .ZN(n35) );
  OAI22D1BWP30P140 U95 ( .A1(n48), .A2(n69), .B1(n44), .B2(n35), .ZN(N313) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[27]), .ZN(n68) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[59]), .ZN(n36) );
  OAI22D1BWP30P140 U98 ( .A1(n48), .A2(n68), .B1(n44), .B2(n36), .ZN(N314) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[28]), .ZN(n67) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[60]), .ZN(n37) );
  OAI22D1BWP30P140 U101 ( .A1(n48), .A2(n67), .B1(n44), .B2(n37), .ZN(N315) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[29]), .ZN(n66) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[61]), .ZN(n38) );
  OAI22D1BWP30P140 U104 ( .A1(n48), .A2(n66), .B1(n44), .B2(n38), .ZN(N316) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[30]), .ZN(n65) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[62]), .ZN(n39) );
  OAI22D1BWP30P140 U107 ( .A1(n48), .A2(n65), .B1(n44), .B2(n39), .ZN(N317) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[31]), .ZN(n64) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[63]), .ZN(n40) );
  OAI22D1BWP30P140 U110 ( .A1(n48), .A2(n64), .B1(n44), .B2(n40), .ZN(N318) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[23]), .ZN(n72) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[55]), .ZN(n41) );
  OAI22D1BWP30P140 U113 ( .A1(n48), .A2(n72), .B1(n47), .B2(n41), .ZN(N310) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[17]), .ZN(n80) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[49]), .ZN(n42) );
  OAI22D1BWP30P140 U116 ( .A1(n45), .A2(n80), .B1(n44), .B2(n42), .ZN(N304) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[18]), .ZN(n79) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[50]), .ZN(n43) );
  OAI22D1BWP30P140 U119 ( .A1(n45), .A2(n79), .B1(n44), .B2(n43), .ZN(N305) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[21]), .ZN(n74) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[53]), .ZN(n46) );
  OAI22D1BWP30P140 U122 ( .A1(n48), .A2(n74), .B1(n47), .B2(n46), .ZN(N308) );
  MUX2NUD1BWP30P140 U123 ( .I0(n51), .I1(n50), .S(i_cmd[0]), .ZN(n52) );
  ND2OPTIBD1BWP30P140 U124 ( .A1(n53), .A2(n52), .ZN(n54) );
  INVD2BWP30P140 U125 ( .I(n54), .ZN(n77) );
  MOAI22D1BWP30P140 U126 ( .A1(n55), .A2(n62), .B1(i_data_bus[36]), .B2(n89), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n62), .B1(i_data_bus[37]), .B2(n89), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n62), .B1(i_data_bus[38]), .B2(n89), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n62), .B1(i_data_bus[39]), .B2(n89), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n62), .B1(i_data_bus[35]), .B2(n89), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n62), .B1(i_data_bus[34]), .B2(n89), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n90), .B1(i_data_bus[33]), .B2(n89), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n75), .B1(i_data_bus[32]), .B2(n89), 
        .ZN(N319) );
  INVD2BWP30P140 U134 ( .I(n77), .ZN(n75) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n90), .B1(i_data_bus[63]), .B2(n89), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n75), .B1(i_data_bus[62]), .B2(n89), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n90), .B1(i_data_bus[61]), .B2(n89), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n75), .B1(i_data_bus[60]), .B2(n89), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n90), .B1(i_data_bus[59]), .B2(n89), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n75), .B1(i_data_bus[58]), .B2(n89), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n90), .B1(i_data_bus[57]), .B2(n89), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n75), .B1(i_data_bus[56]), .B2(n89), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n90), .B1(i_data_bus[55]), .B2(n89), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n75), .B1(i_data_bus[54]), .B2(n89), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n90), .B1(i_data_bus[53]), .B2(n89), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U146 ( .A1(n76), .A2(n75), .B1(i_data_bus[52]), .B2(n89), 
        .ZN(N339) );
  INVD2BWP30P140 U147 ( .I(n77), .ZN(n90) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n90), .B1(i_data_bus[51]), .B2(n89), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n75), .B1(i_data_bus[50]), .B2(n89), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n90), .B1(i_data_bus[49]), .B2(n89), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n75), .B1(i_data_bus[48]), .B2(n89), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n90), .B1(i_data_bus[47]), .B2(n89), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n75), .B1(i_data_bus[46]), .B2(n89), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n90), .B1(i_data_bus[45]), .B2(n89), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n75), .B1(i_data_bus[44]), .B2(n89), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n90), .B1(i_data_bus[43]), .B2(n89), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n75), .B1(i_data_bus[42]), .B2(n89), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n90), .B1(i_data_bus[41]), .B2(n89), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U159 ( .A1(n91), .A2(n75), .B1(i_data_bus[40]), .B2(n89), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_18 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n18), .Z(n89) );
  CKND2D3BWP30P140 U4 ( .A1(n5), .A2(n4), .ZN(n47) );
  NR2D1BWP30P140 U5 ( .A1(n49), .A2(i_cmd[1]), .ZN(n53) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n49), .ZN(n17) );
  INVD1BWP30P140 U7 ( .I(i_cmd[0]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U8 ( .A1(n17), .A2(n3), .ZN(n2) );
  ND2D1BWP30P140 U9 ( .A1(n1), .A2(i_en), .ZN(n49) );
  INVD1BWP30P140 U10 ( .I(n47), .ZN(n6) );
  INVD1BWP30P140 U11 ( .I(n77), .ZN(n62) );
  INVD1BWP30P140 U12 ( .I(n89), .ZN(n19) );
  INVD1BWP30P140 U13 ( .I(n2), .ZN(n11) );
  INVD1BWP30P140 U14 ( .I(rst), .ZN(n1) );
  INVD2BWP30P140 U15 ( .I(i_valid[1]), .ZN(n50) );
  INVD2BWP30P140 U16 ( .I(n11), .ZN(n48) );
  OAI31D1BWP30P140 U17 ( .A1(n49), .A2(n50), .A3(n3), .B(n48), .ZN(N353) );
  INVD1BWP30P140 U18 ( .I(i_data_bus[0]), .ZN(n55) );
  INVD1BWP30P140 U19 ( .I(i_valid[0]), .ZN(n51) );
  MUX2NOPTD2BWP30P140 U20 ( .I0(n51), .I1(n50), .S(i_cmd[1]), .ZN(n5) );
  NR2OPTPAD1BWP30P140 U21 ( .A1(n49), .A2(n3), .ZN(n4) );
  INVD2BWP30P140 U22 ( .I(n6), .ZN(n16) );
  INVD1BWP30P140 U23 ( .I(i_data_bus[32]), .ZN(n7) );
  OAI22D1BWP30P140 U24 ( .A1(n43), .A2(n55), .B1(n16), .B2(n7), .ZN(N287) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[1]), .ZN(n56) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[33]), .ZN(n8) );
  OAI22D1BWP30P140 U27 ( .A1(n48), .A2(n56), .B1(n16), .B2(n8), .ZN(N288) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[2]), .ZN(n57) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[34]), .ZN(n9) );
  OAI22D1BWP30P140 U30 ( .A1(n43), .A2(n57), .B1(n16), .B2(n9), .ZN(N289) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[3]), .ZN(n58) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[35]), .ZN(n10) );
  OAI22D1BWP30P140 U33 ( .A1(n48), .A2(n58), .B1(n16), .B2(n10), .ZN(N290) );
  INVD2BWP30P140 U34 ( .I(n11), .ZN(n43) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[36]), .ZN(n12) );
  OAI22D1BWP30P140 U37 ( .A1(n43), .A2(n59), .B1(n16), .B2(n12), .ZN(N291) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[5]), .ZN(n63) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[37]), .ZN(n13) );
  OAI22D1BWP30P140 U40 ( .A1(n43), .A2(n63), .B1(n16), .B2(n13), .ZN(N292) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[6]), .ZN(n60) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[38]), .ZN(n14) );
  OAI22D1BWP30P140 U43 ( .A1(n43), .A2(n60), .B1(n16), .B2(n14), .ZN(N293) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[7]), .ZN(n61) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[39]), .ZN(n15) );
  OAI22D1BWP30P140 U46 ( .A1(n43), .A2(n61), .B1(n16), .B2(n15), .ZN(N294) );
  INVD1BWP30P140 U47 ( .I(n17), .ZN(n20) );
  INVD1BWP30P140 U48 ( .I(n49), .ZN(n18) );
  OAI21D1BWP30P140 U49 ( .A1(n20), .A2(i_cmd[1]), .B(n19), .ZN(N354) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[24]), .ZN(n71) );
  BUFFD4BWP30P140 U51 ( .I(n47), .Z(n45) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[56]), .ZN(n21) );
  OAI22D1BWP30P140 U53 ( .A1(n48), .A2(n71), .B1(n45), .B2(n21), .ZN(N311) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[30]), .ZN(n65) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[62]), .ZN(n22) );
  OAI22D1BWP30P140 U56 ( .A1(n48), .A2(n65), .B1(n45), .B2(n22), .ZN(N317) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[28]), .ZN(n67) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[60]), .ZN(n23) );
  OAI22D1BWP30P140 U59 ( .A1(n48), .A2(n67), .B1(n45), .B2(n23), .ZN(N315) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[23]), .ZN(n72) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[55]), .ZN(n24) );
  OAI22D1BWP30P140 U62 ( .A1(n48), .A2(n72), .B1(n45), .B2(n24), .ZN(N310) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[25]), .ZN(n70) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[57]), .ZN(n25) );
  OAI22D1BWP30P140 U65 ( .A1(n48), .A2(n70), .B1(n45), .B2(n25), .ZN(N312) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[26]), .ZN(n69) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[58]), .ZN(n26) );
  OAI22D1BWP30P140 U68 ( .A1(n48), .A2(n69), .B1(n45), .B2(n26), .ZN(N313) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[27]), .ZN(n68) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[59]), .ZN(n27) );
  OAI22D1BWP30P140 U71 ( .A1(n48), .A2(n68), .B1(n45), .B2(n27), .ZN(N314) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[29]), .ZN(n66) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[61]), .ZN(n28) );
  OAI22D1BWP30P140 U74 ( .A1(n48), .A2(n66), .B1(n45), .B2(n28), .ZN(N316) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[31]), .ZN(n64) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[63]), .ZN(n29) );
  OAI22D1BWP30P140 U77 ( .A1(n48), .A2(n64), .B1(n45), .B2(n29), .ZN(N318) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n73) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[54]), .ZN(n30) );
  OAI22D1BWP30P140 U80 ( .A1(n48), .A2(n73), .B1(n45), .B2(n30), .ZN(N309) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[21]), .ZN(n74) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[53]), .ZN(n31) );
  OAI22D1BWP30P140 U83 ( .A1(n48), .A2(n74), .B1(n47), .B2(n31), .ZN(N308) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[8]), .ZN(n91) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[40]), .ZN(n32) );
  OAI22D1BWP30P140 U86 ( .A1(n43), .A2(n91), .B1(n45), .B2(n32), .ZN(N295) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[9]), .ZN(n88) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[41]), .ZN(n33) );
  OAI22D1BWP30P140 U89 ( .A1(n43), .A2(n88), .B1(n45), .B2(n33), .ZN(N296) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[10]), .ZN(n87) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[42]), .ZN(n34) );
  OAI22D1BWP30P140 U92 ( .A1(n43), .A2(n87), .B1(n45), .B2(n34), .ZN(N297) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[11]), .ZN(n86) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[43]), .ZN(n35) );
  OAI22D1BWP30P140 U95 ( .A1(n43), .A2(n86), .B1(n45), .B2(n35), .ZN(N298) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[12]), .ZN(n85) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[44]), .ZN(n36) );
  OAI22D1BWP30P140 U98 ( .A1(n43), .A2(n85), .B1(n45), .B2(n36), .ZN(N299) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[13]), .ZN(n84) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[45]), .ZN(n37) );
  OAI22D1BWP30P140 U101 ( .A1(n43), .A2(n84), .B1(n45), .B2(n37), .ZN(N300) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[14]), .ZN(n83) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[46]), .ZN(n38) );
  OAI22D1BWP30P140 U104 ( .A1(n43), .A2(n83), .B1(n45), .B2(n38), .ZN(N301) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[15]), .ZN(n82) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[47]), .ZN(n39) );
  OAI22D1BWP30P140 U107 ( .A1(n43), .A2(n82), .B1(n45), .B2(n39), .ZN(N302) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[16]), .ZN(n81) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[48]), .ZN(n40) );
  OAI22D1BWP30P140 U110 ( .A1(n43), .A2(n81), .B1(n45), .B2(n40), .ZN(N303) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[17]), .ZN(n80) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[49]), .ZN(n41) );
  OAI22D1BWP30P140 U113 ( .A1(n43), .A2(n80), .B1(n45), .B2(n41), .ZN(N304) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[18]), .ZN(n79) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[50]), .ZN(n42) );
  OAI22D1BWP30P140 U116 ( .A1(n43), .A2(n79), .B1(n45), .B2(n42), .ZN(N305) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[51]), .ZN(n44) );
  OAI22D1BWP30P140 U119 ( .A1(n48), .A2(n78), .B1(n45), .B2(n44), .ZN(N306) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[20]), .ZN(n76) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[52]), .ZN(n46) );
  OAI22D1BWP30P140 U122 ( .A1(n48), .A2(n76), .B1(n47), .B2(n46), .ZN(N307) );
  MUX2NUD1BWP30P140 U123 ( .I0(n51), .I1(n50), .S(i_cmd[0]), .ZN(n52) );
  ND2OPTIBD1BWP30P140 U124 ( .A1(n53), .A2(n52), .ZN(n54) );
  INVD2BWP30P140 U125 ( .I(n54), .ZN(n77) );
  MOAI22D1BWP30P140 U126 ( .A1(n55), .A2(n62), .B1(i_data_bus[32]), .B2(n89), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n62), .B1(i_data_bus[33]), .B2(n89), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n62), .B1(i_data_bus[34]), .B2(n89), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n62), .B1(i_data_bus[35]), .B2(n89), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n62), .B1(i_data_bus[36]), .B2(n89), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n62), .B1(i_data_bus[38]), .B2(n89), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n90), .B1(i_data_bus[39]), .B2(n89), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n75), .B1(i_data_bus[37]), .B2(n89), 
        .ZN(N324) );
  INVD2BWP30P140 U134 ( .I(n77), .ZN(n75) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n90), .B1(i_data_bus[63]), .B2(n89), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n75), .B1(i_data_bus[62]), .B2(n89), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n90), .B1(i_data_bus[61]), .B2(n89), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n75), .B1(i_data_bus[60]), .B2(n89), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n90), .B1(i_data_bus[59]), .B2(n89), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n75), .B1(i_data_bus[58]), .B2(n89), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n90), .B1(i_data_bus[57]), .B2(n89), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n75), .B1(i_data_bus[56]), .B2(n89), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n90), .B1(i_data_bus[55]), .B2(n89), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n75), .B1(i_data_bus[54]), .B2(n89), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n90), .B1(i_data_bus[53]), .B2(n89), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U146 ( .A1(n76), .A2(n75), .B1(i_data_bus[52]), .B2(n89), 
        .ZN(N339) );
  INVD2BWP30P140 U147 ( .I(n77), .ZN(n90) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n90), .B1(i_data_bus[51]), .B2(n89), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n75), .B1(i_data_bus[50]), .B2(n89), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n90), .B1(i_data_bus[49]), .B2(n89), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n75), .B1(i_data_bus[48]), .B2(n89), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n90), .B1(i_data_bus[47]), .B2(n89), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n75), .B1(i_data_bus[46]), .B2(n89), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n90), .B1(i_data_bus[45]), .B2(n89), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n75), .B1(i_data_bus[44]), .B2(n89), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n90), .B1(i_data_bus[43]), .B2(n89), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n75), .B1(i_data_bus[42]), .B2(n89), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n90), .B1(i_data_bus[41]), .B2(n89), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U159 ( .A1(n91), .A2(n75), .B1(i_data_bus[40]), .B2(n89), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_19 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  INVD1BWP30P140 U4 ( .I(n4), .ZN(n13) );
  NR2D1BWP30P140 U5 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  INVD1BWP30P140 U7 ( .I(n13), .ZN(n1) );
  INVD1BWP30P140 U8 ( .I(n13), .ZN(n2) );
  BUFFD12BWP30P140 U9 ( .I(n46), .Z(n48) );
  CKND2D3BWP30P140 U10 ( .A1(n7), .A2(n6), .ZN(n46) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U14 ( .I(n13), .ZN(n33) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n13), .ZN(n49) );
  INVD1BWP30P140 U18 ( .I(n67), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n49), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n13), .ZN(n12) );
  INVD1BWP30P140 U24 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U25 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[32]), .ZN(n8) );
  OAI22D1BWP30P140 U27 ( .A1(n2), .A2(n64), .B1(n48), .B2(n8), .ZN(N287) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[1]), .ZN(n57) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[33]), .ZN(n9) );
  OAI22D1BWP30P140 U30 ( .A1(n1), .A2(n57), .B1(n48), .B2(n9), .ZN(N288) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[2]), .ZN(n56) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[34]), .ZN(n10) );
  OAI22D1BWP30P140 U33 ( .A1(n33), .A2(n56), .B1(n48), .B2(n10), .ZN(N289) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[3]), .ZN(n62) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[35]), .ZN(n11) );
  OAI22D1BWP30P140 U36 ( .A1(n12), .A2(n62), .B1(n48), .B2(n11), .ZN(N290) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[36]), .ZN(n14) );
  OAI22D1BWP30P140 U39 ( .A1(n49), .A2(n59), .B1(n48), .B2(n14), .ZN(N291) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[5]), .ZN(n58) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[37]), .ZN(n15) );
  OAI22D1BWP30P140 U42 ( .A1(n49), .A2(n58), .B1(n48), .B2(n15), .ZN(N292) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[6]), .ZN(n61) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[38]), .ZN(n16) );
  OAI22D1BWP30P140 U45 ( .A1(n49), .A2(n61), .B1(n48), .B2(n16), .ZN(N293) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[7]), .ZN(n60) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[39]), .ZN(n17) );
  OAI22D1BWP30P140 U48 ( .A1(n49), .A2(n60), .B1(n46), .B2(n17), .ZN(N294) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[40]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n49), .A2(n65), .B1(n48), .B2(n22), .ZN(N295) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[41]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n1), .A2(n66), .B1(n48), .B2(n23), .ZN(N296) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[10]), .ZN(n81) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[42]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n33), .A2(n81), .B1(n48), .B2(n24), .ZN(N297) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[11]), .ZN(n79) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[43]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n12), .A2(n79), .B1(n48), .B2(n25), .ZN(N298) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[12]), .ZN(n78) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[44]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n2), .A2(n78), .B1(n48), .B2(n26), .ZN(N299) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[13]), .ZN(n77) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[45]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n1), .A2(n77), .B1(n48), .B2(n27), .ZN(N300) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[14]), .ZN(n76) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[46]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n33), .A2(n76), .B1(n48), .B2(n28), .ZN(N301) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[15]), .ZN(n75) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[47]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n12), .A2(n75), .B1(n48), .B2(n29), .ZN(N302) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[16]), .ZN(n74) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[48]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n2), .A2(n74), .B1(n46), .B2(n30), .ZN(N303) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[17]), .ZN(n73) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[49]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n1), .A2(n73), .B1(n48), .B2(n31), .ZN(N304) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[18]), .ZN(n72) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[50]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n33), .A2(n72), .B1(n48), .B2(n32), .ZN(N305) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[19]), .ZN(n71) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[51]), .ZN(n34) );
  OAI22D1BWP30P140 U87 ( .A1(n12), .A2(n71), .B1(n48), .B2(n34), .ZN(N306) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[20]), .ZN(n70) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[52]), .ZN(n35) );
  OAI22D1BWP30P140 U90 ( .A1(n2), .A2(n70), .B1(n48), .B2(n35), .ZN(N307) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[21]), .ZN(n69) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[53]), .ZN(n36) );
  OAI22D1BWP30P140 U93 ( .A1(n1), .A2(n69), .B1(n48), .B2(n36), .ZN(N308) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[22]), .ZN(n68) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[54]), .ZN(n37) );
  OAI22D1BWP30P140 U96 ( .A1(n33), .A2(n68), .B1(n48), .B2(n37), .ZN(N309) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[23]), .ZN(n92) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[55]), .ZN(n38) );
  OAI22D1BWP30P140 U99 ( .A1(n12), .A2(n92), .B1(n48), .B2(n38), .ZN(N310) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[24]), .ZN(n89) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[56]), .ZN(n39) );
  OAI22D1BWP30P140 U102 ( .A1(n2), .A2(n89), .B1(n48), .B2(n39), .ZN(N311) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[25]), .ZN(n88) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[57]), .ZN(n40) );
  OAI22D1BWP30P140 U105 ( .A1(n1), .A2(n88), .B1(n48), .B2(n40), .ZN(N312) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[26]), .ZN(n87) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[58]), .ZN(n41) );
  OAI22D1BWP30P140 U108 ( .A1(n33), .A2(n87), .B1(n48), .B2(n41), .ZN(N313) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[59]), .ZN(n42) );
  OAI22D1BWP30P140 U111 ( .A1(n12), .A2(n86), .B1(n48), .B2(n42), .ZN(N314) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[28]), .ZN(n85) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[60]), .ZN(n43) );
  OAI22D1BWP30P140 U114 ( .A1(n2), .A2(n85), .B1(n48), .B2(n43), .ZN(N315) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[29]), .ZN(n84) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[61]), .ZN(n44) );
  OAI22D1BWP30P140 U117 ( .A1(n1), .A2(n84), .B1(n48), .B2(n44), .ZN(N316) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[30]), .ZN(n83) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[62]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n33), .A2(n83), .B1(n48), .B2(n45), .ZN(N317) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[31]), .ZN(n82) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[63]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n12), .A2(n82), .B1(n48), .B2(n47), .ZN(N318) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n67) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n91), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  INVD2BWP30P140 U135 ( .I(n67), .ZN(n80) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n80), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n80), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  INVD2BWP30P140 U138 ( .I(n67), .ZN(n91) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n80), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n80), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n80), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n80), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n80), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n80), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n80), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n80), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n80), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n80), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_20 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  INVD1BWP30P140 U4 ( .I(n4), .ZN(n13) );
  NR2D1BWP30P140 U5 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  INVD1BWP30P140 U7 ( .I(n13), .ZN(n1) );
  INVD1BWP30P140 U8 ( .I(n13), .ZN(n2) );
  BUFFD12BWP30P140 U9 ( .I(n46), .Z(n48) );
  CKND2D3BWP30P140 U10 ( .A1(n7), .A2(n6), .ZN(n46) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U14 ( .I(n13), .ZN(n33) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n13), .ZN(n49) );
  INVD1BWP30P140 U18 ( .I(n78), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n49), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n13), .ZN(n12) );
  INVD1BWP30P140 U24 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U25 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[32]), .ZN(n8) );
  OAI22D1BWP30P140 U27 ( .A1(n2), .A2(n64), .B1(n48), .B2(n8), .ZN(N287) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[1]), .ZN(n62) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[33]), .ZN(n9) );
  OAI22D1BWP30P140 U30 ( .A1(n1), .A2(n62), .B1(n48), .B2(n9), .ZN(N288) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[2]), .ZN(n61) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[34]), .ZN(n10) );
  OAI22D1BWP30P140 U33 ( .A1(n33), .A2(n61), .B1(n48), .B2(n10), .ZN(N289) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[35]), .ZN(n11) );
  OAI22D1BWP30P140 U36 ( .A1(n12), .A2(n60), .B1(n48), .B2(n11), .ZN(N290) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[36]), .ZN(n14) );
  OAI22D1BWP30P140 U39 ( .A1(n49), .A2(n59), .B1(n48), .B2(n14), .ZN(N291) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[5]), .ZN(n58) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[37]), .ZN(n15) );
  OAI22D1BWP30P140 U42 ( .A1(n49), .A2(n58), .B1(n48), .B2(n15), .ZN(N292) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[39]), .ZN(n16) );
  OAI22D1BWP30P140 U45 ( .A1(n49), .A2(n56), .B1(n48), .B2(n16), .ZN(N294) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[6]), .ZN(n57) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[38]), .ZN(n17) );
  OAI22D1BWP30P140 U48 ( .A1(n49), .A2(n57), .B1(n46), .B2(n17), .ZN(N293) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[8]), .ZN(n92) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[40]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n49), .A2(n92), .B1(n48), .B2(n22), .ZN(N295) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[9]), .ZN(n89) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[41]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n1), .A2(n89), .B1(n48), .B2(n23), .ZN(N296) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[42]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n33), .A2(n88), .B1(n48), .B2(n24), .ZN(N297) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[11]), .ZN(n87) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[43]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n12), .A2(n87), .B1(n48), .B2(n25), .ZN(N298) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[44]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n2), .A2(n86), .B1(n48), .B2(n26), .ZN(N299) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[13]), .ZN(n85) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[45]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n1), .A2(n85), .B1(n48), .B2(n27), .ZN(N300) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[14]), .ZN(n84) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[46]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n33), .A2(n84), .B1(n48), .B2(n28), .ZN(N301) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[15]), .ZN(n83) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[47]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n12), .A2(n83), .B1(n48), .B2(n29), .ZN(N302) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[16]), .ZN(n82) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[48]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n2), .A2(n82), .B1(n46), .B2(n30), .ZN(N303) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[17]), .ZN(n81) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[49]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n1), .A2(n81), .B1(n48), .B2(n31), .ZN(N304) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[18]), .ZN(n80) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[50]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n33), .A2(n80), .B1(n48), .B2(n32), .ZN(N305) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[19]), .ZN(n79) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[51]), .ZN(n34) );
  OAI22D1BWP30P140 U87 ( .A1(n12), .A2(n79), .B1(n48), .B2(n34), .ZN(N306) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[52]), .ZN(n35) );
  OAI22D1BWP30P140 U90 ( .A1(n2), .A2(n77), .B1(n48), .B2(n35), .ZN(N307) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[21]), .ZN(n75) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[53]), .ZN(n36) );
  OAI22D1BWP30P140 U93 ( .A1(n1), .A2(n75), .B1(n48), .B2(n36), .ZN(N308) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[54]), .ZN(n37) );
  OAI22D1BWP30P140 U96 ( .A1(n33), .A2(n74), .B1(n48), .B2(n37), .ZN(N309) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[23]), .ZN(n73) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[55]), .ZN(n38) );
  OAI22D1BWP30P140 U99 ( .A1(n12), .A2(n73), .B1(n48), .B2(n38), .ZN(N310) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[24]), .ZN(n72) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[56]), .ZN(n39) );
  OAI22D1BWP30P140 U102 ( .A1(n2), .A2(n72), .B1(n48), .B2(n39), .ZN(N311) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[25]), .ZN(n71) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[57]), .ZN(n40) );
  OAI22D1BWP30P140 U105 ( .A1(n1), .A2(n71), .B1(n48), .B2(n40), .ZN(N312) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[26]), .ZN(n70) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[58]), .ZN(n41) );
  OAI22D1BWP30P140 U108 ( .A1(n33), .A2(n70), .B1(n48), .B2(n41), .ZN(N313) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[59]), .ZN(n42) );
  OAI22D1BWP30P140 U111 ( .A1(n12), .A2(n69), .B1(n48), .B2(n42), .ZN(N314) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[28]), .ZN(n68) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[60]), .ZN(n43) );
  OAI22D1BWP30P140 U114 ( .A1(n2), .A2(n68), .B1(n48), .B2(n43), .ZN(N315) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[29]), .ZN(n67) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[61]), .ZN(n44) );
  OAI22D1BWP30P140 U117 ( .A1(n1), .A2(n67), .B1(n48), .B2(n44), .ZN(N316) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[30]), .ZN(n66) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[62]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n33), .A2(n66), .B1(n48), .B2(n45), .ZN(N317) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[31]), .ZN(n65) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[63]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n12), .A2(n65), .B1(n48), .B2(n47), .ZN(N318) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n78) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  INVD2BWP30P140 U135 ( .I(n78), .ZN(n76) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_21 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  INVD1BWP30P140 U4 ( .I(n4), .ZN(n10) );
  NR2D1BWP30P140 U5 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  INVD1BWP30P140 U7 ( .I(n10), .ZN(n1) );
  INVD1BWP30P140 U8 ( .I(n10), .ZN(n2) );
  BUFFD12BWP30P140 U9 ( .I(n46), .Z(n48) );
  CKND2D3BWP30P140 U10 ( .A1(n7), .A2(n6), .ZN(n46) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U14 ( .I(n10), .ZN(n33) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n10), .ZN(n49) );
  INVD1BWP30P140 U18 ( .I(n71), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n49), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(i_data_bus[5]), .ZN(n58) );
  INVD1BWP30P140 U24 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[37]), .ZN(n8) );
  OAI22D1BWP30P140 U26 ( .A1(n49), .A2(n58), .B1(n48), .B2(n8), .ZN(N292) );
  INVD1BWP30P140 U27 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[36]), .ZN(n9) );
  OAI22D1BWP30P140 U29 ( .A1(n49), .A2(n59), .B1(n48), .B2(n9), .ZN(N291) );
  INVD1BWP30P140 U30 ( .I(n10), .ZN(n15) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[35]), .ZN(n11) );
  OAI22D1BWP30P140 U33 ( .A1(n2), .A2(n60), .B1(n48), .B2(n11), .ZN(N290) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[2]), .ZN(n61) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[34]), .ZN(n12) );
  OAI22D1BWP30P140 U36 ( .A1(n1), .A2(n61), .B1(n48), .B2(n12), .ZN(N289) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[1]), .ZN(n62) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[33]), .ZN(n13) );
  OAI22D1BWP30P140 U39 ( .A1(n33), .A2(n62), .B1(n48), .B2(n13), .ZN(N288) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[32]), .ZN(n14) );
  OAI22D1BWP30P140 U42 ( .A1(n15), .A2(n64), .B1(n48), .B2(n14), .ZN(N287) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[39]), .ZN(n16) );
  OAI22D1BWP30P140 U45 ( .A1(n49), .A2(n56), .B1(n48), .B2(n16), .ZN(N294) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[6]), .ZN(n57) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[38]), .ZN(n17) );
  OAI22D1BWP30P140 U48 ( .A1(n49), .A2(n57), .B1(n46), .B2(n17), .ZN(N293) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[8]), .ZN(n84) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[40]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n49), .A2(n84), .B1(n48), .B2(n22), .ZN(N295) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[9]), .ZN(n82) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[41]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n1), .A2(n82), .B1(n48), .B2(n23), .ZN(N296) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[10]), .ZN(n81) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[42]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n33), .A2(n81), .B1(n48), .B2(n24), .ZN(N297) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[11]), .ZN(n80) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[43]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n15), .A2(n80), .B1(n48), .B2(n25), .ZN(N298) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[12]), .ZN(n79) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[44]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n2), .A2(n79), .B1(n48), .B2(n26), .ZN(N299) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[13]), .ZN(n78) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[45]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n1), .A2(n78), .B1(n48), .B2(n27), .ZN(N300) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[14]), .ZN(n77) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[46]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n33), .A2(n77), .B1(n48), .B2(n28), .ZN(N301) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[15]), .ZN(n76) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[47]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n15), .A2(n76), .B1(n48), .B2(n29), .ZN(N302) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[16]), .ZN(n75) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[48]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n2), .A2(n75), .B1(n46), .B2(n30), .ZN(N303) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[49]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n1), .A2(n74), .B1(n48), .B2(n31), .ZN(N304) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[18]), .ZN(n73) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[50]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n33), .A2(n73), .B1(n48), .B2(n32), .ZN(N305) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[19]), .ZN(n72) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[51]), .ZN(n34) );
  OAI22D1BWP30P140 U87 ( .A1(n15), .A2(n72), .B1(n48), .B2(n34), .ZN(N306) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[20]), .ZN(n70) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[52]), .ZN(n35) );
  OAI22D1BWP30P140 U90 ( .A1(n2), .A2(n70), .B1(n48), .B2(n35), .ZN(N307) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[21]), .ZN(n69) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[53]), .ZN(n36) );
  OAI22D1BWP30P140 U93 ( .A1(n1), .A2(n69), .B1(n48), .B2(n36), .ZN(N308) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[22]), .ZN(n68) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[54]), .ZN(n37) );
  OAI22D1BWP30P140 U96 ( .A1(n33), .A2(n68), .B1(n48), .B2(n37), .ZN(N309) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[23]), .ZN(n67) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[55]), .ZN(n38) );
  OAI22D1BWP30P140 U99 ( .A1(n15), .A2(n67), .B1(n48), .B2(n38), .ZN(N310) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[24]), .ZN(n66) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[56]), .ZN(n39) );
  OAI22D1BWP30P140 U102 ( .A1(n2), .A2(n66), .B1(n48), .B2(n39), .ZN(N311) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[25]), .ZN(n65) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[57]), .ZN(n40) );
  OAI22D1BWP30P140 U105 ( .A1(n1), .A2(n65), .B1(n48), .B2(n40), .ZN(N312) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[26]), .ZN(n92) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[58]), .ZN(n41) );
  OAI22D1BWP30P140 U108 ( .A1(n33), .A2(n92), .B1(n48), .B2(n41), .ZN(N313) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[27]), .ZN(n89) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[59]), .ZN(n42) );
  OAI22D1BWP30P140 U111 ( .A1(n15), .A2(n89), .B1(n48), .B2(n42), .ZN(N314) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[28]), .ZN(n88) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[60]), .ZN(n43) );
  OAI22D1BWP30P140 U114 ( .A1(n2), .A2(n88), .B1(n48), .B2(n43), .ZN(N315) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[29]), .ZN(n87) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[61]), .ZN(n44) );
  OAI22D1BWP30P140 U117 ( .A1(n1), .A2(n87), .B1(n48), .B2(n44), .ZN(N316) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[30]), .ZN(n86) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[62]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n33), .A2(n86), .B1(n48), .B2(n45), .ZN(N317) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[31]), .ZN(n85) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[63]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n15), .A2(n85), .B1(n48), .B2(n47), .ZN(N318) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n71) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n83), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  INVD2BWP30P140 U135 ( .I(n71), .ZN(n91) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  INVD2BWP30P140 U142 ( .I(n71), .ZN(n83) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n83), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n83), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n83), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n83), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n83), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n83), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n83), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n83), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n83), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n83), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n83), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n83), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_22 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  NR2D1BWP30P140 U4 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INR2D1BWP30P140 U5 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  INVD1BWP30P140 U6 ( .I(n4), .ZN(n12) );
  INVD1BWP30P140 U7 ( .I(n12), .ZN(n1) );
  INVD1BWP30P140 U8 ( .I(n12), .ZN(n2) );
  BUFFD12BWP30P140 U9 ( .I(n46), .Z(n48) );
  CKND2D3BWP30P140 U10 ( .A1(n7), .A2(n6), .ZN(n46) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U14 ( .I(n12), .ZN(n49) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n12), .ZN(n35) );
  INVD1BWP30P140 U18 ( .I(n76), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n35), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD1BWP30P140 U24 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[39]), .ZN(n8) );
  OAI22D1BWP30P140 U26 ( .A1(n35), .A2(n64), .B1(n48), .B2(n8), .ZN(N294) );
  INVD1BWP30P140 U27 ( .I(i_data_bus[6]), .ZN(n62) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[38]), .ZN(n9) );
  OAI22D1BWP30P140 U29 ( .A1(n35), .A2(n62), .B1(n48), .B2(n9), .ZN(N293) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[5]), .ZN(n61) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[37]), .ZN(n10) );
  OAI22D1BWP30P140 U32 ( .A1(n35), .A2(n61), .B1(n48), .B2(n10), .ZN(N292) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[36]), .ZN(n11) );
  OAI22D1BWP30P140 U35 ( .A1(n35), .A2(n60), .B1(n48), .B2(n11), .ZN(N291) );
  INVD1BWP30P140 U36 ( .I(n12), .ZN(n17) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[3]), .ZN(n59) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[35]), .ZN(n13) );
  OAI22D1BWP30P140 U39 ( .A1(n1), .A2(n59), .B1(n48), .B2(n13), .ZN(N290) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[2]), .ZN(n58) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[34]), .ZN(n14) );
  OAI22D1BWP30P140 U42 ( .A1(n49), .A2(n58), .B1(n48), .B2(n14), .ZN(N289) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[1]), .ZN(n57) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[33]), .ZN(n15) );
  OAI22D1BWP30P140 U45 ( .A1(n17), .A2(n57), .B1(n48), .B2(n15), .ZN(N288) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[0]), .ZN(n56) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[32]), .ZN(n16) );
  OAI22D1BWP30P140 U48 ( .A1(n2), .A2(n56), .B1(n46), .B2(n16), .ZN(N287) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[63]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n17), .A2(n92), .B1(n48), .B2(n22), .ZN(N318) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[30]), .ZN(n87) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[62]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n2), .A2(n87), .B1(n48), .B2(n23), .ZN(N317) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[29]), .ZN(n86) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[61]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n1), .A2(n86), .B1(n48), .B2(n24), .ZN(N316) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[28]), .ZN(n85) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[60]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n49), .A2(n85), .B1(n48), .B2(n25), .ZN(N315) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[27]), .ZN(n84) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[59]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n17), .A2(n84), .B1(n48), .B2(n26), .ZN(N314) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[26]), .ZN(n83) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[58]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n2), .A2(n83), .B1(n48), .B2(n27), .ZN(N313) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[25]), .ZN(n82) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[57]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n1), .A2(n82), .B1(n48), .B2(n28), .ZN(N312) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[24]), .ZN(n81) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[56]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n49), .A2(n81), .B1(n48), .B2(n29), .ZN(N311) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[23]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[55]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n17), .A2(n80), .B1(n46), .B2(n30), .ZN(N310) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[22]), .ZN(n79) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[54]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n2), .A2(n79), .B1(n48), .B2(n31), .ZN(N309) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[21]), .ZN(n78) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[53]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n1), .A2(n78), .B1(n48), .B2(n32), .ZN(N308) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[52]), .ZN(n33) );
  OAI22D1BWP30P140 U87 ( .A1(n49), .A2(n77), .B1(n48), .B2(n33), .ZN(N307) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[19]), .ZN(n75) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[51]), .ZN(n34) );
  OAI22D1BWP30P140 U90 ( .A1(n17), .A2(n75), .B1(n48), .B2(n34), .ZN(N306) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[18]), .ZN(n74) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[50]), .ZN(n36) );
  OAI22D1BWP30P140 U93 ( .A1(n35), .A2(n74), .B1(n48), .B2(n36), .ZN(N305) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[17]), .ZN(n73) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[49]), .ZN(n37) );
  OAI22D1BWP30P140 U96 ( .A1(n1), .A2(n73), .B1(n48), .B2(n37), .ZN(N304) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[16]), .ZN(n72) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[48]), .ZN(n38) );
  OAI22D1BWP30P140 U99 ( .A1(n49), .A2(n72), .B1(n48), .B2(n38), .ZN(N303) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[15]), .ZN(n71) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[47]), .ZN(n39) );
  OAI22D1BWP30P140 U102 ( .A1(n17), .A2(n71), .B1(n48), .B2(n39), .ZN(N302) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[14]), .ZN(n70) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[46]), .ZN(n40) );
  OAI22D1BWP30P140 U105 ( .A1(n2), .A2(n70), .B1(n48), .B2(n40), .ZN(N301) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[13]), .ZN(n69) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[45]), .ZN(n41) );
  OAI22D1BWP30P140 U108 ( .A1(n1), .A2(n69), .B1(n48), .B2(n41), .ZN(N300) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[12]), .ZN(n68) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[44]), .ZN(n42) );
  OAI22D1BWP30P140 U111 ( .A1(n49), .A2(n68), .B1(n48), .B2(n42), .ZN(N299) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[11]), .ZN(n67) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[43]), .ZN(n43) );
  OAI22D1BWP30P140 U114 ( .A1(n17), .A2(n67), .B1(n48), .B2(n43), .ZN(N298) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[10]), .ZN(n66) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[42]), .ZN(n44) );
  OAI22D1BWP30P140 U117 ( .A1(n2), .A2(n66), .B1(n48), .B2(n44), .ZN(N297) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[9]), .ZN(n65) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[41]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n1), .A2(n65), .B1(n48), .B2(n45), .ZN(N296) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[8]), .ZN(n89) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[40]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n49), .A2(n89), .B1(n48), .B2(n47), .ZN(N295) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n76) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n91), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  INVD2BWP30P140 U135 ( .I(n76), .ZN(n88) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n88), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n88), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n88), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n88), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n88), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n88), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n88), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n88), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n88), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n88), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n88), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U147 ( .I(n76), .ZN(n91) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U156 ( .A1(n85), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U157 ( .A1(n86), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U158 ( .A1(n87), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n88), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_23 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  INVD1BWP30P140 U4 ( .I(n4), .ZN(n12) );
  NR2D1BWP30P140 U5 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  INVD1BWP30P140 U7 ( .I(n12), .ZN(n1) );
  INVD1BWP30P140 U8 ( .I(n12), .ZN(n2) );
  BUFFD12BWP30P140 U9 ( .I(n46), .Z(n48) );
  CKND2D3BWP30P140 U10 ( .A1(n7), .A2(n6), .ZN(n46) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U14 ( .I(n12), .ZN(n44) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n12), .ZN(n49) );
  INVD1BWP30P140 U18 ( .I(n78), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n49), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(i_data_bus[7]), .ZN(n61) );
  INVD1BWP30P140 U24 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[39]), .ZN(n8) );
  OAI22D1BWP30P140 U26 ( .A1(n49), .A2(n61), .B1(n48), .B2(n8), .ZN(N294) );
  INVD1BWP30P140 U27 ( .I(i_data_bus[6]), .ZN(n62) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[38]), .ZN(n9) );
  OAI22D1BWP30P140 U29 ( .A1(n49), .A2(n62), .B1(n48), .B2(n9), .ZN(N293) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[5]), .ZN(n64) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[37]), .ZN(n10) );
  OAI22D1BWP30P140 U32 ( .A1(n49), .A2(n64), .B1(n48), .B2(n10), .ZN(N292) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[36]), .ZN(n11) );
  OAI22D1BWP30P140 U35 ( .A1(n49), .A2(n60), .B1(n48), .B2(n11), .ZN(N291) );
  INVD1BWP30P140 U36 ( .I(n12), .ZN(n17) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[3]), .ZN(n59) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[35]), .ZN(n13) );
  OAI22D1BWP30P140 U39 ( .A1(n1), .A2(n59), .B1(n48), .B2(n13), .ZN(N290) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[2]), .ZN(n58) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[34]), .ZN(n14) );
  OAI22D1BWP30P140 U42 ( .A1(n44), .A2(n58), .B1(n48), .B2(n14), .ZN(N289) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[1]), .ZN(n57) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[33]), .ZN(n15) );
  OAI22D1BWP30P140 U45 ( .A1(n17), .A2(n57), .B1(n48), .B2(n15), .ZN(N288) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[0]), .ZN(n56) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[32]), .ZN(n16) );
  OAI22D1BWP30P140 U48 ( .A1(n2), .A2(n56), .B1(n46), .B2(n16), .ZN(N287) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[61]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n17), .A2(n88), .B1(n48), .B2(n22), .ZN(N316) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[60]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n2), .A2(n87), .B1(n48), .B2(n23), .ZN(N315) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[59]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n1), .A2(n86), .B1(n48), .B2(n24), .ZN(N314) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[58]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n44), .A2(n85), .B1(n48), .B2(n25), .ZN(N313) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[57]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n17), .A2(n84), .B1(n48), .B2(n26), .ZN(N312) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[56]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n2), .A2(n83), .B1(n48), .B2(n27), .ZN(N311) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[55]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n1), .A2(n82), .B1(n48), .B2(n28), .ZN(N310) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[54]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n44), .A2(n81), .B1(n48), .B2(n29), .ZN(N309) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[53]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n17), .A2(n80), .B1(n48), .B2(n30), .ZN(N308) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[52]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n2), .A2(n79), .B1(n48), .B2(n31), .ZN(N307) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[19]), .ZN(n77) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[51]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n1), .A2(n77), .B1(n48), .B2(n32), .ZN(N306) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[50]), .ZN(n33) );
  OAI22D1BWP30P140 U87 ( .A1(n49), .A2(n75), .B1(n48), .B2(n33), .ZN(N305) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[49]), .ZN(n34) );
  OAI22D1BWP30P140 U90 ( .A1(n1), .A2(n74), .B1(n48), .B2(n34), .ZN(N304) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[48]), .ZN(n35) );
  OAI22D1BWP30P140 U93 ( .A1(n44), .A2(n73), .B1(n48), .B2(n35), .ZN(N303) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[47]), .ZN(n36) );
  OAI22D1BWP30P140 U96 ( .A1(n17), .A2(n72), .B1(n48), .B2(n36), .ZN(N302) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[46]), .ZN(n37) );
  OAI22D1BWP30P140 U99 ( .A1(n2), .A2(n71), .B1(n48), .B2(n37), .ZN(N301) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[45]), .ZN(n38) );
  OAI22D1BWP30P140 U102 ( .A1(n1), .A2(n70), .B1(n48), .B2(n38), .ZN(N300) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[44]), .ZN(n39) );
  OAI22D1BWP30P140 U105 ( .A1(n44), .A2(n69), .B1(n48), .B2(n39), .ZN(N299) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[43]), .ZN(n40) );
  OAI22D1BWP30P140 U108 ( .A1(n17), .A2(n68), .B1(n46), .B2(n40), .ZN(N298) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[42]), .ZN(n41) );
  OAI22D1BWP30P140 U111 ( .A1(n2), .A2(n67), .B1(n48), .B2(n41), .ZN(N297) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[41]), .ZN(n42) );
  OAI22D1BWP30P140 U114 ( .A1(n1), .A2(n66), .B1(n48), .B2(n42), .ZN(N296) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[40]), .ZN(n43) );
  OAI22D1BWP30P140 U117 ( .A1(n44), .A2(n65), .B1(n48), .B2(n43), .ZN(N295) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[62]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n44), .A2(n89), .B1(n48), .B2(n45), .ZN(N317) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[63]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n17), .A2(n92), .B1(n48), .B2(n47), .ZN(N318) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n78) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n91), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  INVD2BWP30P140 U135 ( .I(n78), .ZN(n76) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_24 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  INVD1BWP30P140 U4 ( .I(n4), .ZN(n10) );
  NR2D1BWP30P140 U5 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  INVD1BWP30P140 U7 ( .I(n10), .ZN(n1) );
  INVD1BWP30P140 U8 ( .I(n10), .ZN(n2) );
  BUFFD12BWP30P140 U9 ( .I(n46), .Z(n48) );
  CKND2D3BWP30P140 U10 ( .A1(n7), .A2(n6), .ZN(n46) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U14 ( .I(n10), .ZN(n49) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n10), .ZN(n35) );
  INVD1BWP30P140 U18 ( .I(n78), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n35), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n10), .ZN(n17) );
  INVD1BWP30P140 U24 ( .I(i_data_bus[1]), .ZN(n64) );
  INVD1BWP30P140 U25 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[33]), .ZN(n8) );
  OAI22D1BWP30P140 U27 ( .A1(n1), .A2(n64), .B1(n48), .B2(n8), .ZN(N288) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[0]), .ZN(n62) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[32]), .ZN(n9) );
  OAI22D1BWP30P140 U30 ( .A1(n49), .A2(n62), .B1(n48), .B2(n9), .ZN(N287) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[7]), .ZN(n61) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[39]), .ZN(n11) );
  OAI22D1BWP30P140 U33 ( .A1(n35), .A2(n61), .B1(n48), .B2(n11), .ZN(N294) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[6]), .ZN(n60) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[38]), .ZN(n12) );
  OAI22D1BWP30P140 U36 ( .A1(n35), .A2(n60), .B1(n48), .B2(n12), .ZN(N293) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[37]), .ZN(n13) );
  OAI22D1BWP30P140 U39 ( .A1(n35), .A2(n59), .B1(n48), .B2(n13), .ZN(N292) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[4]), .ZN(n58) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[36]), .ZN(n14) );
  OAI22D1BWP30P140 U42 ( .A1(n35), .A2(n58), .B1(n48), .B2(n14), .ZN(N291) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[3]), .ZN(n57) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[35]), .ZN(n15) );
  OAI22D1BWP30P140 U45 ( .A1(n17), .A2(n57), .B1(n48), .B2(n15), .ZN(N290) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[2]), .ZN(n56) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[34]), .ZN(n16) );
  OAI22D1BWP30P140 U48 ( .A1(n2), .A2(n56), .B1(n46), .B2(n16), .ZN(N289) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[63]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n17), .A2(n92), .B1(n48), .B2(n22), .ZN(N318) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[62]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n2), .A2(n89), .B1(n48), .B2(n23), .ZN(N317) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[61]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n1), .A2(n88), .B1(n48), .B2(n24), .ZN(N316) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[60]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n49), .A2(n87), .B1(n48), .B2(n25), .ZN(N315) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[59]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n17), .A2(n86), .B1(n48), .B2(n26), .ZN(N314) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[58]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n2), .A2(n85), .B1(n48), .B2(n27), .ZN(N313) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[57]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n1), .A2(n84), .B1(n48), .B2(n28), .ZN(N312) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[56]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n49), .A2(n83), .B1(n48), .B2(n29), .ZN(N311) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[55]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n17), .A2(n82), .B1(n46), .B2(n30), .ZN(N310) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[54]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n2), .A2(n81), .B1(n48), .B2(n31), .ZN(N309) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[53]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n1), .A2(n80), .B1(n48), .B2(n32), .ZN(N308) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[52]), .ZN(n33) );
  OAI22D1BWP30P140 U87 ( .A1(n49), .A2(n79), .B1(n48), .B2(n33), .ZN(N307) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[19]), .ZN(n77) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[51]), .ZN(n34) );
  OAI22D1BWP30P140 U90 ( .A1(n17), .A2(n77), .B1(n48), .B2(n34), .ZN(N306) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[50]), .ZN(n36) );
  OAI22D1BWP30P140 U93 ( .A1(n35), .A2(n75), .B1(n48), .B2(n36), .ZN(N305) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[49]), .ZN(n37) );
  OAI22D1BWP30P140 U96 ( .A1(n1), .A2(n74), .B1(n48), .B2(n37), .ZN(N304) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[48]), .ZN(n38) );
  OAI22D1BWP30P140 U99 ( .A1(n49), .A2(n73), .B1(n48), .B2(n38), .ZN(N303) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[47]), .ZN(n39) );
  OAI22D1BWP30P140 U102 ( .A1(n17), .A2(n72), .B1(n48), .B2(n39), .ZN(N302) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[46]), .ZN(n40) );
  OAI22D1BWP30P140 U105 ( .A1(n2), .A2(n71), .B1(n48), .B2(n40), .ZN(N301) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[45]), .ZN(n41) );
  OAI22D1BWP30P140 U108 ( .A1(n1), .A2(n70), .B1(n48), .B2(n41), .ZN(N300) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[44]), .ZN(n42) );
  OAI22D1BWP30P140 U111 ( .A1(n49), .A2(n69), .B1(n48), .B2(n42), .ZN(N299) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[43]), .ZN(n43) );
  OAI22D1BWP30P140 U114 ( .A1(n17), .A2(n68), .B1(n48), .B2(n43), .ZN(N298) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[42]), .ZN(n44) );
  OAI22D1BWP30P140 U117 ( .A1(n2), .A2(n67), .B1(n48), .B2(n44), .ZN(N297) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[41]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n1), .A2(n66), .B1(n48), .B2(n45), .ZN(N296) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[40]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n49), .A2(n65), .B1(n48), .B2(n47), .ZN(N295) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n78) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n91), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  INVD2BWP30P140 U135 ( .I(n78), .ZN(n76) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_25 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  BUFFD6BWP30P140 U3 ( .I(n46), .Z(n48) );
  AN3D4BWP30P140 U4 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  INVD1BWP30P140 U5 ( .I(n4), .ZN(n9) );
  NR2D1BWP30P140 U6 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INR2D1BWP30P140 U7 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  INVD1BWP30P140 U8 ( .I(n9), .ZN(n1) );
  INVD1BWP30P140 U9 ( .I(n9), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U10 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U11 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U12 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U13 ( .I(n9), .ZN(n34) );
  CKND2D2BWP30P140 U14 ( .A1(n7), .A2(n6), .ZN(n46) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n9), .ZN(n49) );
  INVD1BWP30P140 U18 ( .I(n75), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n49), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD1BWP30P140 U24 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[39]), .ZN(n8) );
  OAI22D1BWP30P140 U26 ( .A1(n49), .A2(n56), .B1(n48), .B2(n8), .ZN(N294) );
  INVD1BWP30P140 U27 ( .I(n9), .ZN(n15) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[2]), .ZN(n61) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[34]), .ZN(n10) );
  OAI22D1BWP30P140 U30 ( .A1(n2), .A2(n61), .B1(n48), .B2(n10), .ZN(N289) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[1]), .ZN(n62) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[33]), .ZN(n11) );
  OAI22D1BWP30P140 U33 ( .A1(n1), .A2(n62), .B1(n48), .B2(n11), .ZN(N288) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[32]), .ZN(n12) );
  OAI22D1BWP30P140 U36 ( .A1(n34), .A2(n64), .B1(n48), .B2(n12), .ZN(N287) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[6]), .ZN(n57) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[38]), .ZN(n13) );
  OAI22D1BWP30P140 U39 ( .A1(n49), .A2(n57), .B1(n48), .B2(n13), .ZN(N293) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[35]), .ZN(n14) );
  OAI22D1BWP30P140 U42 ( .A1(n15), .A2(n60), .B1(n48), .B2(n14), .ZN(N290) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[5]), .ZN(n58) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[37]), .ZN(n16) );
  OAI22D1BWP30P140 U45 ( .A1(n49), .A2(n58), .B1(n48), .B2(n16), .ZN(N292) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[36]), .ZN(n17) );
  OAI22D1BWP30P140 U48 ( .A1(n49), .A2(n59), .B1(n48), .B2(n17), .ZN(N291) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[29]), .ZN(n85) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[61]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n15), .A2(n85), .B1(n48), .B2(n22), .ZN(N316) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[8]), .ZN(n89) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[40]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n49), .A2(n89), .B1(n48), .B2(n23), .ZN(N295) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[9]), .ZN(n92) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[41]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n1), .A2(n92), .B1(n48), .B2(n24), .ZN(N296) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[10]), .ZN(n65) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[42]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n34), .A2(n65), .B1(n48), .B2(n25), .ZN(N297) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[11]), .ZN(n66) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[43]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n15), .A2(n66), .B1(n48), .B2(n26), .ZN(N298) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[12]), .ZN(n67) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[44]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n2), .A2(n67), .B1(n48), .B2(n27), .ZN(N299) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[13]), .ZN(n68) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[45]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n1), .A2(n68), .B1(n48), .B2(n28), .ZN(N300) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[14]), .ZN(n69) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[46]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n34), .A2(n69), .B1(n48), .B2(n29), .ZN(N301) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[15]), .ZN(n70) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[47]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n15), .A2(n70), .B1(n48), .B2(n30), .ZN(N302) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[16]), .ZN(n71) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[48]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n2), .A2(n71), .B1(n48), .B2(n31), .ZN(N303) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[17]), .ZN(n72) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[49]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n1), .A2(n72), .B1(n48), .B2(n32), .ZN(N304) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[18]), .ZN(n73) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[50]), .ZN(n33) );
  OAI22D1BWP30P140 U87 ( .A1(n34), .A2(n73), .B1(n48), .B2(n33), .ZN(N305) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[19]), .ZN(n74) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[51]), .ZN(n35) );
  OAI22D1BWP30P140 U90 ( .A1(n2), .A2(n74), .B1(n48), .B2(n35), .ZN(N306) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[20]), .ZN(n76) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[52]), .ZN(n36) );
  OAI22D1BWP30P140 U93 ( .A1(n1), .A2(n76), .B1(n48), .B2(n36), .ZN(N307) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[21]), .ZN(n77) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[53]), .ZN(n37) );
  OAI22D1BWP30P140 U96 ( .A1(n34), .A2(n77), .B1(n48), .B2(n37), .ZN(N308) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[22]), .ZN(n78) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[54]), .ZN(n38) );
  OAI22D1BWP30P140 U99 ( .A1(n15), .A2(n78), .B1(n48), .B2(n38), .ZN(N309) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[23]), .ZN(n79) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[55]), .ZN(n39) );
  OAI22D1BWP30P140 U102 ( .A1(n2), .A2(n79), .B1(n48), .B2(n39), .ZN(N310) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[24]), .ZN(n80) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[56]), .ZN(n40) );
  OAI22D1BWP30P140 U105 ( .A1(n1), .A2(n80), .B1(n48), .B2(n40), .ZN(N311) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[25]), .ZN(n81) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[57]), .ZN(n41) );
  OAI22D1BWP30P140 U108 ( .A1(n34), .A2(n81), .B1(n48), .B2(n41), .ZN(N312) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[26]), .ZN(n82) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[58]), .ZN(n42) );
  OAI22D1BWP30P140 U111 ( .A1(n15), .A2(n82), .B1(n48), .B2(n42), .ZN(N313) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[27]), .ZN(n83) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[59]), .ZN(n43) );
  OAI22D1BWP30P140 U114 ( .A1(n2), .A2(n83), .B1(n48), .B2(n43), .ZN(N314) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[28]), .ZN(n84) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[60]), .ZN(n44) );
  OAI22D1BWP30P140 U117 ( .A1(n1), .A2(n84), .B1(n48), .B2(n44), .ZN(N315) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[31]), .ZN(n88) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[63]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n34), .A2(n88), .B1(n48), .B2(n45), .ZN(N318) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[30]), .ZN(n86) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[62]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n15), .A2(n86), .B1(n48), .B2(n47), .ZN(N317) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n75) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n87), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  INVD2BWP30P140 U135 ( .I(n75), .ZN(n91) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U146 ( .I(n75), .ZN(n87) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n87), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n87), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n87), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n87), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n87), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n87), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n87), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n87), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n87), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U156 ( .A1(n85), .A2(n87), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U157 ( .A1(n86), .A2(n87), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n87), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_26 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  INVD1BWP30P140 U4 ( .I(n4), .ZN(n12) );
  NR2D1BWP30P140 U5 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  INVD1BWP30P140 U7 ( .I(n12), .ZN(n1) );
  INVD1BWP30P140 U8 ( .I(n12), .ZN(n2) );
  BUFFD12BWP30P140 U9 ( .I(n46), .Z(n48) );
  CKND2D3BWP30P140 U10 ( .A1(n7), .A2(n6), .ZN(n46) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U14 ( .I(n12), .ZN(n33) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n12), .ZN(n49) );
  INVD1BWP30P140 U18 ( .I(n78), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n49), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(i_data_bus[7]), .ZN(n59) );
  INVD1BWP30P140 U24 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[39]), .ZN(n8) );
  OAI22D1BWP30P140 U26 ( .A1(n49), .A2(n59), .B1(n48), .B2(n8), .ZN(N294) );
  INVD1BWP30P140 U27 ( .I(i_data_bus[6]), .ZN(n56) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[38]), .ZN(n9) );
  OAI22D1BWP30P140 U29 ( .A1(n49), .A2(n56), .B1(n48), .B2(n9), .ZN(N293) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[5]), .ZN(n57) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[37]), .ZN(n10) );
  OAI22D1BWP30P140 U32 ( .A1(n49), .A2(n57), .B1(n48), .B2(n10), .ZN(N292) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[36]), .ZN(n11) );
  OAI22D1BWP30P140 U35 ( .A1(n49), .A2(n62), .B1(n48), .B2(n11), .ZN(N291) );
  INVD1BWP30P140 U36 ( .I(n12), .ZN(n17) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[3]), .ZN(n58) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[35]), .ZN(n13) );
  OAI22D1BWP30P140 U39 ( .A1(n1), .A2(n58), .B1(n48), .B2(n13), .ZN(N290) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[34]), .ZN(n14) );
  OAI22D1BWP30P140 U42 ( .A1(n33), .A2(n60), .B1(n48), .B2(n14), .ZN(N289) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[1]), .ZN(n61) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[33]), .ZN(n15) );
  OAI22D1BWP30P140 U45 ( .A1(n17), .A2(n61), .B1(n48), .B2(n15), .ZN(N288) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[32]), .ZN(n16) );
  OAI22D1BWP30P140 U48 ( .A1(n2), .A2(n64), .B1(n46), .B2(n16), .ZN(N287) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[40]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n49), .A2(n65), .B1(n48), .B2(n22), .ZN(N295) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[41]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n1), .A2(n66), .B1(n48), .B2(n23), .ZN(N296) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[42]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n33), .A2(n67), .B1(n48), .B2(n24), .ZN(N297) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[43]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n17), .A2(n68), .B1(n48), .B2(n25), .ZN(N298) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[44]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n2), .A2(n69), .B1(n48), .B2(n26), .ZN(N299) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[45]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n1), .A2(n70), .B1(n48), .B2(n27), .ZN(N300) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[46]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n33), .A2(n71), .B1(n48), .B2(n28), .ZN(N301) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[47]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n17), .A2(n72), .B1(n48), .B2(n29), .ZN(N302) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[48]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n2), .A2(n73), .B1(n46), .B2(n30), .ZN(N303) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[49]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n1), .A2(n74), .B1(n48), .B2(n31), .ZN(N304) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[50]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n33), .A2(n75), .B1(n48), .B2(n32), .ZN(N305) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[19]), .ZN(n77) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[51]), .ZN(n34) );
  OAI22D1BWP30P140 U87 ( .A1(n17), .A2(n77), .B1(n48), .B2(n34), .ZN(N306) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[52]), .ZN(n35) );
  OAI22D1BWP30P140 U90 ( .A1(n2), .A2(n79), .B1(n48), .B2(n35), .ZN(N307) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[53]), .ZN(n36) );
  OAI22D1BWP30P140 U93 ( .A1(n1), .A2(n80), .B1(n48), .B2(n36), .ZN(N308) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[54]), .ZN(n37) );
  OAI22D1BWP30P140 U96 ( .A1(n33), .A2(n81), .B1(n48), .B2(n37), .ZN(N309) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[55]), .ZN(n38) );
  OAI22D1BWP30P140 U99 ( .A1(n17), .A2(n82), .B1(n48), .B2(n38), .ZN(N310) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[56]), .ZN(n39) );
  OAI22D1BWP30P140 U102 ( .A1(n2), .A2(n83), .B1(n48), .B2(n39), .ZN(N311) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[57]), .ZN(n40) );
  OAI22D1BWP30P140 U105 ( .A1(n1), .A2(n84), .B1(n48), .B2(n40), .ZN(N312) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[58]), .ZN(n41) );
  OAI22D1BWP30P140 U108 ( .A1(n33), .A2(n85), .B1(n48), .B2(n41), .ZN(N313) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[59]), .ZN(n42) );
  OAI22D1BWP30P140 U111 ( .A1(n17), .A2(n86), .B1(n48), .B2(n42), .ZN(N314) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[60]), .ZN(n43) );
  OAI22D1BWP30P140 U114 ( .A1(n2), .A2(n87), .B1(n48), .B2(n43), .ZN(N315) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[61]), .ZN(n44) );
  OAI22D1BWP30P140 U117 ( .A1(n1), .A2(n88), .B1(n48), .B2(n44), .ZN(N316) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[62]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n33), .A2(n89), .B1(n48), .B2(n45), .ZN(N317) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[63]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n17), .A2(n92), .B1(n48), .B2(n47), .ZN(N318) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n78) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n91), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  INVD2BWP30P140 U135 ( .I(n78), .ZN(n76) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_27 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  INVD1BWP30P140 U4 ( .I(n4), .ZN(n12) );
  NR2D1BWP30P140 U5 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  INVD1BWP30P140 U7 ( .I(n12), .ZN(n1) );
  INVD1BWP30P140 U8 ( .I(n12), .ZN(n2) );
  BUFFD12BWP30P140 U9 ( .I(n46), .Z(n48) );
  CKND2D3BWP30P140 U10 ( .A1(n7), .A2(n6), .ZN(n46) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U14 ( .I(n12), .ZN(n49) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n12), .ZN(n40) );
  INVD1BWP30P140 U18 ( .I(n78), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n40), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD1BWP30P140 U24 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[39]), .ZN(n8) );
  OAI22D1BWP30P140 U26 ( .A1(n40), .A2(n56), .B1(n48), .B2(n8), .ZN(N294) );
  INVD1BWP30P140 U27 ( .I(i_data_bus[6]), .ZN(n57) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[38]), .ZN(n9) );
  OAI22D1BWP30P140 U29 ( .A1(n40), .A2(n57), .B1(n48), .B2(n9), .ZN(N293) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[5]), .ZN(n58) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[37]), .ZN(n10) );
  OAI22D1BWP30P140 U32 ( .A1(n40), .A2(n58), .B1(n48), .B2(n10), .ZN(N292) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[36]), .ZN(n11) );
  OAI22D1BWP30P140 U35 ( .A1(n40), .A2(n59), .B1(n48), .B2(n11), .ZN(N291) );
  INVD1BWP30P140 U36 ( .I(n12), .ZN(n17) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[35]), .ZN(n13) );
  OAI22D1BWP30P140 U39 ( .A1(n1), .A2(n60), .B1(n48), .B2(n13), .ZN(N290) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[2]), .ZN(n61) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[34]), .ZN(n14) );
  OAI22D1BWP30P140 U42 ( .A1(n49), .A2(n61), .B1(n48), .B2(n14), .ZN(N289) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[1]), .ZN(n62) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[33]), .ZN(n15) );
  OAI22D1BWP30P140 U45 ( .A1(n17), .A2(n62), .B1(n48), .B2(n15), .ZN(N288) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[32]), .ZN(n16) );
  OAI22D1BWP30P140 U48 ( .A1(n2), .A2(n64), .B1(n46), .B2(n16), .ZN(N287) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[46]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n40), .A2(n71), .B1(n48), .B2(n22), .ZN(N301) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[47]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n1), .A2(n72), .B1(n48), .B2(n23), .ZN(N302) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[48]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n49), .A2(n73), .B1(n48), .B2(n24), .ZN(N303) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[49]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n17), .A2(n74), .B1(n48), .B2(n25), .ZN(N304) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[50]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n2), .A2(n75), .B1(n48), .B2(n26), .ZN(N305) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[19]), .ZN(n77) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n17), .A2(n77), .B1(n48), .B2(n27), .ZN(N306) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[52]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n2), .A2(n79), .B1(n48), .B2(n28), .ZN(N307) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[53]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n1), .A2(n80), .B1(n48), .B2(n29), .ZN(N308) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n49), .A2(n81), .B1(n48), .B2(n30), .ZN(N309) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[55]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n17), .A2(n82), .B1(n48), .B2(n31), .ZN(N310) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[56]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n2), .A2(n83), .B1(n48), .B2(n32), .ZN(N311) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[57]), .ZN(n33) );
  OAI22D1BWP30P140 U87 ( .A1(n1), .A2(n84), .B1(n48), .B2(n33), .ZN(N312) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[58]), .ZN(n34) );
  OAI22D1BWP30P140 U90 ( .A1(n49), .A2(n85), .B1(n48), .B2(n34), .ZN(N313) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[59]), .ZN(n35) );
  OAI22D1BWP30P140 U93 ( .A1(n17), .A2(n86), .B1(n48), .B2(n35), .ZN(N314) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[60]), .ZN(n36) );
  OAI22D1BWP30P140 U96 ( .A1(n2), .A2(n87), .B1(n46), .B2(n36), .ZN(N315) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[61]), .ZN(n37) );
  OAI22D1BWP30P140 U99 ( .A1(n1), .A2(n88), .B1(n48), .B2(n37), .ZN(N316) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[62]), .ZN(n38) );
  OAI22D1BWP30P140 U102 ( .A1(n49), .A2(n89), .B1(n48), .B2(n38), .ZN(N317) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[63]), .ZN(n39) );
  OAI22D1BWP30P140 U105 ( .A1(n17), .A2(n92), .B1(n48), .B2(n39), .ZN(N318) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[45]), .ZN(n41) );
  OAI22D1BWP30P140 U108 ( .A1(n1), .A2(n70), .B1(n48), .B2(n41), .ZN(N300) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[43]), .ZN(n42) );
  OAI22D1BWP30P140 U111 ( .A1(n49), .A2(n68), .B1(n48), .B2(n42), .ZN(N298) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[42]), .ZN(n43) );
  OAI22D1BWP30P140 U114 ( .A1(n17), .A2(n67), .B1(n48), .B2(n43), .ZN(N297) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[44]), .ZN(n44) );
  OAI22D1BWP30P140 U117 ( .A1(n2), .A2(n69), .B1(n48), .B2(n44), .ZN(N299) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[41]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n1), .A2(n66), .B1(n48), .B2(n45), .ZN(N296) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[40]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n49), .A2(n65), .B1(n48), .B2(n47), .ZN(N295) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n78) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  INVD2BWP30P140 U135 ( .I(n78), .ZN(n76) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_28 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  INVD1BWP30P140 U4 ( .I(n4), .ZN(n12) );
  NR2D1BWP30P140 U5 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  INVD1BWP30P140 U7 ( .I(n12), .ZN(n1) );
  INVD1BWP30P140 U8 ( .I(n12), .ZN(n2) );
  BUFFD12BWP30P140 U9 ( .I(n46), .Z(n48) );
  CKND2D3BWP30P140 U10 ( .A1(n7), .A2(n6), .ZN(n46) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U14 ( .I(n12), .ZN(n33) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n12), .ZN(n49) );
  INVD1BWP30P140 U18 ( .I(n78), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n49), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD1BWP30P140 U24 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[39]), .ZN(n8) );
  OAI22D1BWP30P140 U26 ( .A1(n49), .A2(n56), .B1(n48), .B2(n8), .ZN(N294) );
  INVD1BWP30P140 U27 ( .I(i_data_bus[6]), .ZN(n57) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[38]), .ZN(n9) );
  OAI22D1BWP30P140 U29 ( .A1(n49), .A2(n57), .B1(n48), .B2(n9), .ZN(N293) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[5]), .ZN(n58) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[37]), .ZN(n10) );
  OAI22D1BWP30P140 U32 ( .A1(n49), .A2(n58), .B1(n48), .B2(n10), .ZN(N292) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[36]), .ZN(n11) );
  OAI22D1BWP30P140 U35 ( .A1(n49), .A2(n59), .B1(n48), .B2(n11), .ZN(N291) );
  INVD1BWP30P140 U36 ( .I(n12), .ZN(n17) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[35]), .ZN(n13) );
  OAI22D1BWP30P140 U39 ( .A1(n1), .A2(n60), .B1(n48), .B2(n13), .ZN(N290) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[2]), .ZN(n61) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[34]), .ZN(n14) );
  OAI22D1BWP30P140 U42 ( .A1(n33), .A2(n61), .B1(n48), .B2(n14), .ZN(N289) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[1]), .ZN(n62) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[33]), .ZN(n15) );
  OAI22D1BWP30P140 U45 ( .A1(n17), .A2(n62), .B1(n48), .B2(n15), .ZN(N288) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[32]), .ZN(n16) );
  OAI22D1BWP30P140 U48 ( .A1(n2), .A2(n64), .B1(n46), .B2(n16), .ZN(N287) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[40]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n49), .A2(n65), .B1(n48), .B2(n22), .ZN(N295) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[41]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n1), .A2(n66), .B1(n48), .B2(n23), .ZN(N296) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[42]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n33), .A2(n67), .B1(n48), .B2(n24), .ZN(N297) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[43]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n17), .A2(n68), .B1(n48), .B2(n25), .ZN(N298) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[44]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n2), .A2(n69), .B1(n48), .B2(n26), .ZN(N299) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[45]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n1), .A2(n70), .B1(n48), .B2(n27), .ZN(N300) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[46]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n33), .A2(n71), .B1(n48), .B2(n28), .ZN(N301) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[47]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n17), .A2(n72), .B1(n48), .B2(n29), .ZN(N302) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[48]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n2), .A2(n73), .B1(n46), .B2(n30), .ZN(N303) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[49]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n1), .A2(n74), .B1(n48), .B2(n31), .ZN(N304) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[50]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n33), .A2(n75), .B1(n48), .B2(n32), .ZN(N305) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[19]), .ZN(n77) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[51]), .ZN(n34) );
  OAI22D1BWP30P140 U87 ( .A1(n17), .A2(n77), .B1(n48), .B2(n34), .ZN(N306) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[52]), .ZN(n35) );
  OAI22D1BWP30P140 U90 ( .A1(n2), .A2(n79), .B1(n48), .B2(n35), .ZN(N307) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[53]), .ZN(n36) );
  OAI22D1BWP30P140 U93 ( .A1(n1), .A2(n80), .B1(n48), .B2(n36), .ZN(N308) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[54]), .ZN(n37) );
  OAI22D1BWP30P140 U96 ( .A1(n33), .A2(n81), .B1(n48), .B2(n37), .ZN(N309) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[55]), .ZN(n38) );
  OAI22D1BWP30P140 U99 ( .A1(n17), .A2(n82), .B1(n48), .B2(n38), .ZN(N310) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[56]), .ZN(n39) );
  OAI22D1BWP30P140 U102 ( .A1(n2), .A2(n83), .B1(n48), .B2(n39), .ZN(N311) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[57]), .ZN(n40) );
  OAI22D1BWP30P140 U105 ( .A1(n1), .A2(n84), .B1(n48), .B2(n40), .ZN(N312) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[58]), .ZN(n41) );
  OAI22D1BWP30P140 U108 ( .A1(n33), .A2(n85), .B1(n48), .B2(n41), .ZN(N313) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[59]), .ZN(n42) );
  OAI22D1BWP30P140 U111 ( .A1(n17), .A2(n86), .B1(n48), .B2(n42), .ZN(N314) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[60]), .ZN(n43) );
  OAI22D1BWP30P140 U114 ( .A1(n2), .A2(n87), .B1(n48), .B2(n43), .ZN(N315) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[61]), .ZN(n44) );
  OAI22D1BWP30P140 U117 ( .A1(n1), .A2(n88), .B1(n48), .B2(n44), .ZN(N316) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[62]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n33), .A2(n89), .B1(n48), .B2(n45), .ZN(N317) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[63]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n17), .A2(n92), .B1(n48), .B2(n47), .ZN(N318) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n78) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  INVD2BWP30P140 U135 ( .I(n78), .ZN(n76) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_29 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  INVD1BWP30P140 U4 ( .I(n4), .ZN(n12) );
  NR2D1BWP30P140 U5 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  INVD1BWP30P140 U7 ( .I(n12), .ZN(n1) );
  INVD1BWP30P140 U8 ( .I(n12), .ZN(n2) );
  BUFFD12BWP30P140 U9 ( .I(n46), .Z(n48) );
  CKND2D3BWP30P140 U10 ( .A1(n7), .A2(n6), .ZN(n46) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U14 ( .I(n12), .ZN(n34) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n12), .ZN(n49) );
  INVD1BWP30P140 U18 ( .I(n75), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n49), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(i_data_bus[7]), .ZN(n58) );
  INVD1BWP30P140 U24 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[39]), .ZN(n8) );
  OAI22D1BWP30P140 U26 ( .A1(n49), .A2(n58), .B1(n48), .B2(n8), .ZN(N294) );
  INVD1BWP30P140 U27 ( .I(i_data_bus[6]), .ZN(n56) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[38]), .ZN(n9) );
  OAI22D1BWP30P140 U29 ( .A1(n49), .A2(n56), .B1(n48), .B2(n9), .ZN(N293) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[5]), .ZN(n57) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[37]), .ZN(n10) );
  OAI22D1BWP30P140 U32 ( .A1(n49), .A2(n57), .B1(n48), .B2(n10), .ZN(N292) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[36]), .ZN(n11) );
  OAI22D1BWP30P140 U35 ( .A1(n49), .A2(n59), .B1(n48), .B2(n11), .ZN(N291) );
  INVD1BWP30P140 U36 ( .I(n12), .ZN(n17) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[35]), .ZN(n13) );
  OAI22D1BWP30P140 U39 ( .A1(n1), .A2(n60), .B1(n48), .B2(n13), .ZN(N290) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[2]), .ZN(n61) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[34]), .ZN(n14) );
  OAI22D1BWP30P140 U42 ( .A1(n34), .A2(n61), .B1(n48), .B2(n14), .ZN(N289) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[1]), .ZN(n62) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[33]), .ZN(n15) );
  OAI22D1BWP30P140 U45 ( .A1(n17), .A2(n62), .B1(n48), .B2(n15), .ZN(N288) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[32]), .ZN(n16) );
  OAI22D1BWP30P140 U48 ( .A1(n2), .A2(n64), .B1(n46), .B2(n16), .ZN(N287) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[19]), .ZN(n76) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[51]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n17), .A2(n76), .B1(n48), .B2(n22), .ZN(N306) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[18]), .ZN(n77) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[50]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n49), .A2(n77), .B1(n48), .B2(n23), .ZN(N305) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[17]), .ZN(n78) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[49]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n1), .A2(n78), .B1(n48), .B2(n24), .ZN(N304) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[16]), .ZN(n79) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[48]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n34), .A2(n79), .B1(n48), .B2(n25), .ZN(N303) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[15]), .ZN(n80) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[47]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n17), .A2(n80), .B1(n48), .B2(n26), .ZN(N302) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[14]), .ZN(n81) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[46]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n2), .A2(n81), .B1(n48), .B2(n27), .ZN(N301) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[8]), .ZN(n88) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[40]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n1), .A2(n88), .B1(n48), .B2(n28), .ZN(N295) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[9]), .ZN(n86) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[41]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n34), .A2(n86), .B1(n48), .B2(n29), .ZN(N296) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[13]), .ZN(n82) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[45]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n17), .A2(n82), .B1(n46), .B2(n30), .ZN(N300) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[12]), .ZN(n83) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[44]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n2), .A2(n83), .B1(n48), .B2(n31), .ZN(N299) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[10]), .ZN(n85) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[42]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n1), .A2(n85), .B1(n48), .B2(n32), .ZN(N297) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[11]), .ZN(n84) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[43]), .ZN(n33) );
  OAI22D1BWP30P140 U87 ( .A1(n34), .A2(n84), .B1(n48), .B2(n33), .ZN(N298) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[25]), .ZN(n69) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[57]), .ZN(n35) );
  OAI22D1BWP30P140 U90 ( .A1(n2), .A2(n69), .B1(n48), .B2(n35), .ZN(N312) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[26]), .ZN(n68) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[58]), .ZN(n36) );
  OAI22D1BWP30P140 U93 ( .A1(n1), .A2(n68), .B1(n48), .B2(n36), .ZN(N313) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[27]), .ZN(n67) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[59]), .ZN(n37) );
  OAI22D1BWP30P140 U96 ( .A1(n34), .A2(n67), .B1(n48), .B2(n37), .ZN(N314) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[24]), .ZN(n70) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[56]), .ZN(n38) );
  OAI22D1BWP30P140 U99 ( .A1(n17), .A2(n70), .B1(n48), .B2(n38), .ZN(N311) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[28]), .ZN(n66) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[60]), .ZN(n39) );
  OAI22D1BWP30P140 U102 ( .A1(n2), .A2(n66), .B1(n48), .B2(n39), .ZN(N315) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[29]), .ZN(n89) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[61]), .ZN(n40) );
  OAI22D1BWP30P140 U105 ( .A1(n1), .A2(n89), .B1(n48), .B2(n40), .ZN(N316) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[31]), .ZN(n65) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[63]), .ZN(n41) );
  OAI22D1BWP30P140 U108 ( .A1(n34), .A2(n65), .B1(n48), .B2(n41), .ZN(N318) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[20]), .ZN(n74) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[52]), .ZN(n42) );
  OAI22D1BWP30P140 U111 ( .A1(n17), .A2(n74), .B1(n48), .B2(n42), .ZN(N307) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[21]), .ZN(n73) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[53]), .ZN(n43) );
  OAI22D1BWP30P140 U114 ( .A1(n2), .A2(n73), .B1(n48), .B2(n43), .ZN(N308) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[22]), .ZN(n72) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[54]), .ZN(n44) );
  OAI22D1BWP30P140 U117 ( .A1(n1), .A2(n72), .B1(n48), .B2(n44), .ZN(N309) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[23]), .ZN(n71) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[55]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n34), .A2(n71), .B1(n48), .B2(n45), .ZN(N310) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[30]), .ZN(n92) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[62]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n17), .A2(n92), .B1(n48), .B2(n47), .ZN(N317) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n75) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n87), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  INVD2BWP30P140 U135 ( .I(n75), .ZN(n91) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  INVD2BWP30P140 U146 ( .I(n75), .ZN(n87) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n87), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n87), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n87), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n87), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n87), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n87), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n87), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n87), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n87), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U156 ( .A1(n85), .A2(n87), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U157 ( .A1(n86), .A2(n87), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n87), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_30 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  INVD1BWP30P140 U4 ( .I(n4), .ZN(n13) );
  NR2D1BWP30P140 U5 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  INVD1BWP30P140 U7 ( .I(n13), .ZN(n1) );
  INVD1BWP30P140 U8 ( .I(n13), .ZN(n2) );
  BUFFD12BWP30P140 U9 ( .I(n46), .Z(n48) );
  CKND2D3BWP30P140 U10 ( .A1(n7), .A2(n6), .ZN(n46) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U14 ( .I(n13), .ZN(n33) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n13), .ZN(n49) );
  INVD1BWP30P140 U18 ( .I(n72), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n49), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n13), .ZN(n12) );
  INVD1BWP30P140 U24 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U25 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[32]), .ZN(n8) );
  OAI22D1BWP30P140 U27 ( .A1(n2), .A2(n64), .B1(n48), .B2(n8), .ZN(N287) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[1]), .ZN(n62) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[33]), .ZN(n9) );
  OAI22D1BWP30P140 U30 ( .A1(n1), .A2(n62), .B1(n48), .B2(n9), .ZN(N288) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[2]), .ZN(n61) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[34]), .ZN(n10) );
  OAI22D1BWP30P140 U33 ( .A1(n33), .A2(n61), .B1(n48), .B2(n10), .ZN(N289) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[35]), .ZN(n11) );
  OAI22D1BWP30P140 U36 ( .A1(n12), .A2(n60), .B1(n48), .B2(n11), .ZN(N290) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[36]), .ZN(n14) );
  OAI22D1BWP30P140 U39 ( .A1(n49), .A2(n59), .B1(n48), .B2(n14), .ZN(N291) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[5]), .ZN(n58) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[37]), .ZN(n15) );
  OAI22D1BWP30P140 U42 ( .A1(n49), .A2(n58), .B1(n48), .B2(n15), .ZN(N292) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[6]), .ZN(n57) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[38]), .ZN(n16) );
  OAI22D1BWP30P140 U45 ( .A1(n49), .A2(n57), .B1(n48), .B2(n16), .ZN(N293) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[39]), .ZN(n17) );
  OAI22D1BWP30P140 U48 ( .A1(n49), .A2(n56), .B1(n46), .B2(n17), .ZN(N294) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[8]), .ZN(n69) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[40]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n49), .A2(n69), .B1(n48), .B2(n22), .ZN(N295) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[9]), .ZN(n68) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[41]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n1), .A2(n68), .B1(n48), .B2(n23), .ZN(N296) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[42]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n33), .A2(n67), .B1(n48), .B2(n24), .ZN(N297) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[11]), .ZN(n66) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[43]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n12), .A2(n66), .B1(n48), .B2(n25), .ZN(N298) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[12]), .ZN(n65) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[44]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n2), .A2(n65), .B1(n48), .B2(n26), .ZN(N299) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[45]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n1), .A2(n70), .B1(n48), .B2(n27), .ZN(N300) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[46]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n33), .A2(n71), .B1(n48), .B2(n28), .ZN(N301) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[15]), .ZN(n92) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[47]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n12), .A2(n92), .B1(n48), .B2(n29), .ZN(N302) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[16]), .ZN(n89) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[48]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n2), .A2(n89), .B1(n46), .B2(n30), .ZN(N303) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[17]), .ZN(n88) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[49]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n1), .A2(n88), .B1(n48), .B2(n31), .ZN(N304) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[18]), .ZN(n87) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[50]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n33), .A2(n87), .B1(n48), .B2(n32), .ZN(N305) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[19]), .ZN(n86) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[51]), .ZN(n34) );
  OAI22D1BWP30P140 U87 ( .A1(n12), .A2(n86), .B1(n48), .B2(n34), .ZN(N306) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[20]), .ZN(n85) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[52]), .ZN(n35) );
  OAI22D1BWP30P140 U90 ( .A1(n2), .A2(n85), .B1(n48), .B2(n35), .ZN(N307) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[21]), .ZN(n83) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[53]), .ZN(n36) );
  OAI22D1BWP30P140 U93 ( .A1(n1), .A2(n83), .B1(n48), .B2(n36), .ZN(N308) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[22]), .ZN(n82) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[54]), .ZN(n37) );
  OAI22D1BWP30P140 U96 ( .A1(n33), .A2(n82), .B1(n48), .B2(n37), .ZN(N309) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[23]), .ZN(n81) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[55]), .ZN(n38) );
  OAI22D1BWP30P140 U99 ( .A1(n12), .A2(n81), .B1(n48), .B2(n38), .ZN(N310) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[24]), .ZN(n80) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[56]), .ZN(n39) );
  OAI22D1BWP30P140 U102 ( .A1(n2), .A2(n80), .B1(n48), .B2(n39), .ZN(N311) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[25]), .ZN(n79) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[57]), .ZN(n40) );
  OAI22D1BWP30P140 U105 ( .A1(n1), .A2(n79), .B1(n48), .B2(n40), .ZN(N312) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[26]), .ZN(n78) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[58]), .ZN(n41) );
  OAI22D1BWP30P140 U108 ( .A1(n33), .A2(n78), .B1(n48), .B2(n41), .ZN(N313) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[27]), .ZN(n77) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[59]), .ZN(n42) );
  OAI22D1BWP30P140 U111 ( .A1(n12), .A2(n77), .B1(n48), .B2(n42), .ZN(N314) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[28]), .ZN(n76) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[60]), .ZN(n43) );
  OAI22D1BWP30P140 U114 ( .A1(n2), .A2(n76), .B1(n48), .B2(n43), .ZN(N315) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[29]), .ZN(n75) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[61]), .ZN(n44) );
  OAI22D1BWP30P140 U117 ( .A1(n1), .A2(n75), .B1(n48), .B2(n44), .ZN(N316) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[30]), .ZN(n74) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[62]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n33), .A2(n74), .B1(n48), .B2(n45), .ZN(N317) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[31]), .ZN(n73) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[63]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n12), .A2(n73), .B1(n48), .B2(n47), .ZN(N318) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n72) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n84), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  INVD2BWP30P140 U135 ( .I(n72), .ZN(n91) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  INVD2BWP30P140 U143 ( .I(n72), .ZN(n84) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n84), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n84), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n84), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n84), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n84), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n84), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n84), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n84), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n84), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n84), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n84), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n84), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_31 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  INVD1BWP30P140 U4 ( .I(n4), .ZN(n13) );
  NR2D1BWP30P140 U5 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  INVD1BWP30P140 U7 ( .I(n13), .ZN(n1) );
  INVD1BWP30P140 U8 ( .I(n13), .ZN(n2) );
  BUFFD12BWP30P140 U9 ( .I(n46), .Z(n48) );
  CKND2D3BWP30P140 U10 ( .A1(n7), .A2(n6), .ZN(n46) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U14 ( .I(n13), .ZN(n49) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n13), .ZN(n42) );
  INVD1BWP30P140 U18 ( .I(n78), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n42), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n13), .ZN(n12) );
  INVD1BWP30P140 U24 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U25 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[32]), .ZN(n8) );
  OAI22D1BWP30P140 U27 ( .A1(n2), .A2(n64), .B1(n48), .B2(n8), .ZN(N287) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[1]), .ZN(n62) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[33]), .ZN(n9) );
  OAI22D1BWP30P140 U30 ( .A1(n1), .A2(n62), .B1(n48), .B2(n9), .ZN(N288) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[2]), .ZN(n61) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[34]), .ZN(n10) );
  OAI22D1BWP30P140 U33 ( .A1(n49), .A2(n61), .B1(n48), .B2(n10), .ZN(N289) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[35]), .ZN(n11) );
  OAI22D1BWP30P140 U36 ( .A1(n12), .A2(n60), .B1(n48), .B2(n11), .ZN(N290) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[36]), .ZN(n14) );
  OAI22D1BWP30P140 U39 ( .A1(n42), .A2(n59), .B1(n48), .B2(n14), .ZN(N291) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[5]), .ZN(n58) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[37]), .ZN(n15) );
  OAI22D1BWP30P140 U42 ( .A1(n42), .A2(n58), .B1(n48), .B2(n15), .ZN(N292) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[6]), .ZN(n57) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[38]), .ZN(n16) );
  OAI22D1BWP30P140 U45 ( .A1(n42), .A2(n57), .B1(n48), .B2(n16), .ZN(N293) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[39]), .ZN(n17) );
  OAI22D1BWP30P140 U48 ( .A1(n42), .A2(n56), .B1(n46), .B2(n17), .ZN(N294) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[44]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n42), .A2(n86), .B1(n48), .B2(n22), .ZN(N299) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[13]), .ZN(n85) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n1), .A2(n85), .B1(n48), .B2(n23), .ZN(N300) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[14]), .ZN(n84) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n49), .A2(n84), .B1(n48), .B2(n24), .ZN(N301) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n83) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[47]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n12), .A2(n83), .B1(n48), .B2(n25), .ZN(N302) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n82) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[48]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n2), .A2(n82), .B1(n48), .B2(n26), .ZN(N303) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[17]), .ZN(n81) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[49]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n1), .A2(n81), .B1(n48), .B2(n27), .ZN(N304) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[18]), .ZN(n80) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[50]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n49), .A2(n80), .B1(n48), .B2(n28), .ZN(N305) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[19]), .ZN(n79) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[51]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n12), .A2(n79), .B1(n48), .B2(n29), .ZN(N306) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[52]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n2), .A2(n77), .B1(n48), .B2(n30), .ZN(N307) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[21]), .ZN(n75) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[53]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n1), .A2(n75), .B1(n48), .B2(n31), .ZN(N308) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[54]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n49), .A2(n74), .B1(n48), .B2(n32), .ZN(N309) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[23]), .ZN(n73) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[55]), .ZN(n33) );
  OAI22D1BWP30P140 U87 ( .A1(n12), .A2(n73), .B1(n48), .B2(n33), .ZN(N310) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[24]), .ZN(n72) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[56]), .ZN(n34) );
  OAI22D1BWP30P140 U90 ( .A1(n2), .A2(n72), .B1(n48), .B2(n34), .ZN(N311) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[25]), .ZN(n71) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[57]), .ZN(n35) );
  OAI22D1BWP30P140 U93 ( .A1(n1), .A2(n71), .B1(n48), .B2(n35), .ZN(N312) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[26]), .ZN(n70) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[58]), .ZN(n36) );
  OAI22D1BWP30P140 U96 ( .A1(n49), .A2(n70), .B1(n48), .B2(n36), .ZN(N313) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[59]), .ZN(n37) );
  OAI22D1BWP30P140 U99 ( .A1(n12), .A2(n69), .B1(n48), .B2(n37), .ZN(N314) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[28]), .ZN(n68) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[60]), .ZN(n38) );
  OAI22D1BWP30P140 U102 ( .A1(n2), .A2(n68), .B1(n46), .B2(n38), .ZN(N315) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[29]), .ZN(n67) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[61]), .ZN(n39) );
  OAI22D1BWP30P140 U105 ( .A1(n1), .A2(n67), .B1(n48), .B2(n39), .ZN(N316) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[30]), .ZN(n66) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[62]), .ZN(n40) );
  OAI22D1BWP30P140 U108 ( .A1(n49), .A2(n66), .B1(n48), .B2(n40), .ZN(N317) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[31]), .ZN(n65) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[63]), .ZN(n41) );
  OAI22D1BWP30P140 U111 ( .A1(n12), .A2(n65), .B1(n48), .B2(n41), .ZN(N318) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[11]), .ZN(n87) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[43]), .ZN(n43) );
  OAI22D1BWP30P140 U114 ( .A1(n12), .A2(n87), .B1(n48), .B2(n43), .ZN(N298) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[42]), .ZN(n44) );
  OAI22D1BWP30P140 U117 ( .A1(n2), .A2(n88), .B1(n48), .B2(n44), .ZN(N297) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[9]), .ZN(n89) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[41]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n1), .A2(n89), .B1(n48), .B2(n45), .ZN(N296) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[8]), .ZN(n92) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[40]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n49), .A2(n92), .B1(n48), .B2(n47), .ZN(N295) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n78) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  INVD2BWP30P140 U135 ( .I(n78), .ZN(n76) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_32 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  INVD1BWP30P140 U4 ( .I(n4), .ZN(n13) );
  NR2D1BWP30P140 U5 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  INVD1BWP30P140 U7 ( .I(n13), .ZN(n1) );
  INVD1BWP30P140 U8 ( .I(n13), .ZN(n2) );
  BUFFD12BWP30P140 U9 ( .I(n46), .Z(n48) );
  CKND2D3BWP30P140 U10 ( .A1(n7), .A2(n6), .ZN(n46) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U14 ( .I(n13), .ZN(n49) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n13), .ZN(n38) );
  INVD1BWP30P140 U18 ( .I(n68), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n38), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n13), .ZN(n12) );
  INVD1BWP30P140 U24 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD1BWP30P140 U25 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[32]), .ZN(n8) );
  OAI22D1BWP30P140 U27 ( .A1(n2), .A2(n57), .B1(n48), .B2(n8), .ZN(N287) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[1]), .ZN(n56) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[33]), .ZN(n9) );
  OAI22D1BWP30P140 U30 ( .A1(n1), .A2(n56), .B1(n48), .B2(n9), .ZN(N288) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[34]), .ZN(n10) );
  OAI22D1BWP30P140 U33 ( .A1(n49), .A2(n59), .B1(n48), .B2(n10), .ZN(N289) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[3]), .ZN(n58) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[35]), .ZN(n11) );
  OAI22D1BWP30P140 U36 ( .A1(n12), .A2(n58), .B1(n48), .B2(n11), .ZN(N290) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[4]), .ZN(n64) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[36]), .ZN(n14) );
  OAI22D1BWP30P140 U39 ( .A1(n38), .A2(n64), .B1(n48), .B2(n14), .ZN(N291) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[37]), .ZN(n15) );
  OAI22D1BWP30P140 U42 ( .A1(n38), .A2(n62), .B1(n48), .B2(n15), .ZN(N292) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[6]), .ZN(n61) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[38]), .ZN(n16) );
  OAI22D1BWP30P140 U45 ( .A1(n38), .A2(n61), .B1(n48), .B2(n16), .ZN(N293) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[7]), .ZN(n60) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[39]), .ZN(n17) );
  OAI22D1BWP30P140 U48 ( .A1(n38), .A2(n60), .B1(n46), .B2(n17), .ZN(N294) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[31]), .ZN(n69) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[63]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n12), .A2(n69), .B1(n48), .B2(n22), .ZN(N318) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[13]), .ZN(n88) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n38), .A2(n88), .B1(n48), .B2(n23), .ZN(N300) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[14]), .ZN(n87) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n1), .A2(n87), .B1(n48), .B2(n24), .ZN(N301) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[18]), .ZN(n83) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[50]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n49), .A2(n83), .B1(n48), .B2(n25), .ZN(N305) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[19]), .ZN(n82) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[51]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n2), .A2(n82), .B1(n48), .B2(n26), .ZN(N306) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[20]), .ZN(n81) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[52]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n1), .A2(n81), .B1(n48), .B2(n27), .ZN(N307) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[21]), .ZN(n79) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[53]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n49), .A2(n79), .B1(n48), .B2(n28), .ZN(N308) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[22]), .ZN(n78) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[54]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n12), .A2(n78), .B1(n48), .B2(n29), .ZN(N309) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[30]), .ZN(n70) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[62]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n2), .A2(n70), .B1(n48), .B2(n30), .ZN(N317) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[29]), .ZN(n71) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[61]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n1), .A2(n71), .B1(n48), .B2(n31), .ZN(N316) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[28]), .ZN(n72) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[60]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n49), .A2(n72), .B1(n48), .B2(n32), .ZN(N315) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[27]), .ZN(n73) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[59]), .ZN(n33) );
  OAI22D1BWP30P140 U87 ( .A1(n12), .A2(n73), .B1(n48), .B2(n33), .ZN(N314) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[26]), .ZN(n74) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[58]), .ZN(n34) );
  OAI22D1BWP30P140 U90 ( .A1(n2), .A2(n74), .B1(n46), .B2(n34), .ZN(N313) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[25]), .ZN(n75) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[57]), .ZN(n35) );
  OAI22D1BWP30P140 U93 ( .A1(n1), .A2(n75), .B1(n48), .B2(n35), .ZN(N312) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[24]), .ZN(n76) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[56]), .ZN(n36) );
  OAI22D1BWP30P140 U96 ( .A1(n49), .A2(n76), .B1(n48), .B2(n36), .ZN(N311) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[23]), .ZN(n77) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[55]), .ZN(n37) );
  OAI22D1BWP30P140 U99 ( .A1(n12), .A2(n77), .B1(n48), .B2(n37), .ZN(N310) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[40]), .ZN(n39) );
  OAI22D1BWP30P140 U102 ( .A1(n12), .A2(n66), .B1(n48), .B2(n39), .ZN(N295) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[9]), .ZN(n67) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[41]), .ZN(n40) );
  OAI22D1BWP30P140 U105 ( .A1(n2), .A2(n67), .B1(n48), .B2(n40), .ZN(N296) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[10]), .ZN(n65) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[42]), .ZN(n41) );
  OAI22D1BWP30P140 U108 ( .A1(n1), .A2(n65), .B1(n48), .B2(n41), .ZN(N297) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[11]), .ZN(n92) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[43]), .ZN(n42) );
  OAI22D1BWP30P140 U111 ( .A1(n49), .A2(n92), .B1(n48), .B2(n42), .ZN(N298) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[12]), .ZN(n89) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[44]), .ZN(n43) );
  OAI22D1BWP30P140 U114 ( .A1(n12), .A2(n89), .B1(n48), .B2(n43), .ZN(N299) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[15]), .ZN(n86) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[47]), .ZN(n44) );
  OAI22D1BWP30P140 U117 ( .A1(n2), .A2(n86), .B1(n48), .B2(n44), .ZN(N302) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[16]), .ZN(n85) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[48]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n1), .A2(n85), .B1(n48), .B2(n45), .ZN(N303) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[17]), .ZN(n84) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[49]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n49), .A2(n84), .B1(n48), .B2(n47), .ZN(N304) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n68) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n80), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  INVD2BWP30P140 U135 ( .I(n68), .ZN(n91) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  INVD2BWP30P140 U139 ( .I(n68), .ZN(n80) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n80), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n80), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n80), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n80), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n80), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n80), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n80), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n80), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n80), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n80), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n80), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n80), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_33 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  INVD1BWP30P140 U4 ( .I(n4), .ZN(n13) );
  NR2D1BWP30P140 U5 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  INVD1BWP30P140 U7 ( .I(n13), .ZN(n1) );
  INVD1BWP30P140 U8 ( .I(n13), .ZN(n2) );
  BUFFD12BWP30P140 U9 ( .I(n46), .Z(n48) );
  CKND2D3BWP30P140 U10 ( .A1(n7), .A2(n6), .ZN(n46) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U14 ( .I(n13), .ZN(n33) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n13), .ZN(n49) );
  INVD1BWP30P140 U18 ( .I(n78), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n49), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n13), .ZN(n12) );
  INVD1BWP30P140 U24 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U25 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[32]), .ZN(n8) );
  OAI22D1BWP30P140 U27 ( .A1(n2), .A2(n64), .B1(n48), .B2(n8), .ZN(N287) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[1]), .ZN(n62) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[33]), .ZN(n9) );
  OAI22D1BWP30P140 U30 ( .A1(n1), .A2(n62), .B1(n48), .B2(n9), .ZN(N288) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[2]), .ZN(n61) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[34]), .ZN(n10) );
  OAI22D1BWP30P140 U33 ( .A1(n33), .A2(n61), .B1(n48), .B2(n10), .ZN(N289) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[35]), .ZN(n11) );
  OAI22D1BWP30P140 U36 ( .A1(n12), .A2(n60), .B1(n48), .B2(n11), .ZN(N290) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[36]), .ZN(n14) );
  OAI22D1BWP30P140 U39 ( .A1(n49), .A2(n59), .B1(n48), .B2(n14), .ZN(N291) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[5]), .ZN(n58) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[37]), .ZN(n15) );
  OAI22D1BWP30P140 U42 ( .A1(n49), .A2(n58), .B1(n48), .B2(n15), .ZN(N292) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[6]), .ZN(n57) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[38]), .ZN(n16) );
  OAI22D1BWP30P140 U45 ( .A1(n49), .A2(n57), .B1(n48), .B2(n16), .ZN(N293) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[39]), .ZN(n17) );
  OAI22D1BWP30P140 U48 ( .A1(n49), .A2(n56), .B1(n46), .B2(n17), .ZN(N294) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[8]), .ZN(n92) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[40]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n49), .A2(n92), .B1(n48), .B2(n22), .ZN(N295) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[9]), .ZN(n89) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[41]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n1), .A2(n89), .B1(n48), .B2(n23), .ZN(N296) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[42]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n33), .A2(n88), .B1(n48), .B2(n24), .ZN(N297) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[11]), .ZN(n87) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[43]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n12), .A2(n87), .B1(n48), .B2(n25), .ZN(N298) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[44]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n2), .A2(n86), .B1(n48), .B2(n26), .ZN(N299) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[13]), .ZN(n85) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[45]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n1), .A2(n85), .B1(n48), .B2(n27), .ZN(N300) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[14]), .ZN(n84) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[46]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n33), .A2(n84), .B1(n48), .B2(n28), .ZN(N301) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[15]), .ZN(n83) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[47]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n12), .A2(n83), .B1(n48), .B2(n29), .ZN(N302) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[16]), .ZN(n82) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[48]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n2), .A2(n82), .B1(n46), .B2(n30), .ZN(N303) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[17]), .ZN(n81) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[49]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n1), .A2(n81), .B1(n48), .B2(n31), .ZN(N304) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[18]), .ZN(n80) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[50]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n33), .A2(n80), .B1(n48), .B2(n32), .ZN(N305) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[19]), .ZN(n79) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[51]), .ZN(n34) );
  OAI22D1BWP30P140 U87 ( .A1(n12), .A2(n79), .B1(n48), .B2(n34), .ZN(N306) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[52]), .ZN(n35) );
  OAI22D1BWP30P140 U90 ( .A1(n2), .A2(n77), .B1(n48), .B2(n35), .ZN(N307) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[21]), .ZN(n75) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[53]), .ZN(n36) );
  OAI22D1BWP30P140 U93 ( .A1(n1), .A2(n75), .B1(n48), .B2(n36), .ZN(N308) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[54]), .ZN(n37) );
  OAI22D1BWP30P140 U96 ( .A1(n33), .A2(n74), .B1(n48), .B2(n37), .ZN(N309) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[23]), .ZN(n73) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[55]), .ZN(n38) );
  OAI22D1BWP30P140 U99 ( .A1(n12), .A2(n73), .B1(n48), .B2(n38), .ZN(N310) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[24]), .ZN(n72) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[56]), .ZN(n39) );
  OAI22D1BWP30P140 U102 ( .A1(n2), .A2(n72), .B1(n48), .B2(n39), .ZN(N311) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[25]), .ZN(n71) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[57]), .ZN(n40) );
  OAI22D1BWP30P140 U105 ( .A1(n1), .A2(n71), .B1(n48), .B2(n40), .ZN(N312) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[26]), .ZN(n70) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[58]), .ZN(n41) );
  OAI22D1BWP30P140 U108 ( .A1(n33), .A2(n70), .B1(n48), .B2(n41), .ZN(N313) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[59]), .ZN(n42) );
  OAI22D1BWP30P140 U111 ( .A1(n12), .A2(n69), .B1(n48), .B2(n42), .ZN(N314) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[28]), .ZN(n68) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[60]), .ZN(n43) );
  OAI22D1BWP30P140 U114 ( .A1(n2), .A2(n68), .B1(n48), .B2(n43), .ZN(N315) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[29]), .ZN(n67) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[61]), .ZN(n44) );
  OAI22D1BWP30P140 U117 ( .A1(n1), .A2(n67), .B1(n48), .B2(n44), .ZN(N316) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[30]), .ZN(n66) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[62]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n33), .A2(n66), .B1(n48), .B2(n45), .ZN(N317) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[31]), .ZN(n65) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[63]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n12), .A2(n65), .B1(n48), .B2(n47), .ZN(N318) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n78) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  INVD2BWP30P140 U135 ( .I(n78), .ZN(n76) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_34 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  INVD1BWP30P140 U4 ( .I(n4), .ZN(n13) );
  NR2D1BWP30P140 U5 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  INVD1BWP30P140 U7 ( .I(n13), .ZN(n1) );
  INVD1BWP30P140 U8 ( .I(n13), .ZN(n2) );
  BUFFD12BWP30P140 U9 ( .I(n46), .Z(n48) );
  CKND2D3BWP30P140 U10 ( .A1(n7), .A2(n6), .ZN(n46) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U14 ( .I(n13), .ZN(n33) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n13), .ZN(n49) );
  INVD1BWP30P140 U18 ( .I(n76), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n49), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n13), .ZN(n12) );
  INVD1BWP30P140 U24 ( .I(i_data_bus[0]), .ZN(n56) );
  INVD1BWP30P140 U25 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[32]), .ZN(n8) );
  OAI22D1BWP30P140 U27 ( .A1(n2), .A2(n56), .B1(n48), .B2(n8), .ZN(N287) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[1]), .ZN(n57) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[33]), .ZN(n9) );
  OAI22D1BWP30P140 U30 ( .A1(n1), .A2(n57), .B1(n48), .B2(n9), .ZN(N288) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[2]), .ZN(n58) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[34]), .ZN(n10) );
  OAI22D1BWP30P140 U33 ( .A1(n33), .A2(n58), .B1(n48), .B2(n10), .ZN(N289) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[3]), .ZN(n59) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[35]), .ZN(n11) );
  OAI22D1BWP30P140 U36 ( .A1(n12), .A2(n59), .B1(n48), .B2(n11), .ZN(N290) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[36]), .ZN(n14) );
  OAI22D1BWP30P140 U39 ( .A1(n49), .A2(n60), .B1(n48), .B2(n14), .ZN(N291) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[5]), .ZN(n61) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[37]), .ZN(n15) );
  OAI22D1BWP30P140 U42 ( .A1(n49), .A2(n61), .B1(n48), .B2(n15), .ZN(N292) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[6]), .ZN(n62) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[38]), .ZN(n16) );
  OAI22D1BWP30P140 U45 ( .A1(n49), .A2(n62), .B1(n48), .B2(n16), .ZN(N293) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[39]), .ZN(n17) );
  OAI22D1BWP30P140 U48 ( .A1(n49), .A2(n64), .B1(n46), .B2(n17), .ZN(N294) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[8]), .ZN(n89) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[40]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n49), .A2(n89), .B1(n48), .B2(n22), .ZN(N295) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[9]), .ZN(n87) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[41]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n1), .A2(n87), .B1(n48), .B2(n23), .ZN(N296) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[10]), .ZN(n86) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[42]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n33), .A2(n86), .B1(n48), .B2(n24), .ZN(N297) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[11]), .ZN(n85) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[43]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n12), .A2(n85), .B1(n48), .B2(n25), .ZN(N298) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[12]), .ZN(n84) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[44]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n2), .A2(n84), .B1(n48), .B2(n26), .ZN(N299) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[13]), .ZN(n83) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[45]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n1), .A2(n83), .B1(n48), .B2(n27), .ZN(N300) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[14]), .ZN(n82) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[46]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n33), .A2(n82), .B1(n48), .B2(n28), .ZN(N301) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[15]), .ZN(n81) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[47]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n12), .A2(n81), .B1(n48), .B2(n29), .ZN(N302) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[16]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[48]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n2), .A2(n80), .B1(n46), .B2(n30), .ZN(N303) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[17]), .ZN(n79) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[49]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n1), .A2(n79), .B1(n48), .B2(n31), .ZN(N304) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[18]), .ZN(n78) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[50]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n33), .A2(n78), .B1(n48), .B2(n32), .ZN(N305) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[19]), .ZN(n77) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[51]), .ZN(n34) );
  OAI22D1BWP30P140 U87 ( .A1(n12), .A2(n77), .B1(n48), .B2(n34), .ZN(N306) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[20]), .ZN(n75) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[52]), .ZN(n35) );
  OAI22D1BWP30P140 U90 ( .A1(n2), .A2(n75), .B1(n48), .B2(n35), .ZN(N307) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[21]), .ZN(n74) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[53]), .ZN(n36) );
  OAI22D1BWP30P140 U93 ( .A1(n1), .A2(n74), .B1(n48), .B2(n36), .ZN(N308) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[22]), .ZN(n73) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[54]), .ZN(n37) );
  OAI22D1BWP30P140 U96 ( .A1(n33), .A2(n73), .B1(n48), .B2(n37), .ZN(N309) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[23]), .ZN(n72) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[55]), .ZN(n38) );
  OAI22D1BWP30P140 U99 ( .A1(n12), .A2(n72), .B1(n48), .B2(n38), .ZN(N310) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[24]), .ZN(n71) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[56]), .ZN(n39) );
  OAI22D1BWP30P140 U102 ( .A1(n2), .A2(n71), .B1(n48), .B2(n39), .ZN(N311) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[25]), .ZN(n70) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[57]), .ZN(n40) );
  OAI22D1BWP30P140 U105 ( .A1(n1), .A2(n70), .B1(n48), .B2(n40), .ZN(N312) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[26]), .ZN(n69) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[58]), .ZN(n41) );
  OAI22D1BWP30P140 U108 ( .A1(n33), .A2(n69), .B1(n48), .B2(n41), .ZN(N313) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[27]), .ZN(n68) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[59]), .ZN(n42) );
  OAI22D1BWP30P140 U111 ( .A1(n12), .A2(n68), .B1(n48), .B2(n42), .ZN(N314) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[28]), .ZN(n67) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[60]), .ZN(n43) );
  OAI22D1BWP30P140 U114 ( .A1(n2), .A2(n67), .B1(n48), .B2(n43), .ZN(N315) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[29]), .ZN(n66) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[61]), .ZN(n44) );
  OAI22D1BWP30P140 U117 ( .A1(n1), .A2(n66), .B1(n48), .B2(n44), .ZN(N316) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[30]), .ZN(n65) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[62]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n33), .A2(n65), .B1(n48), .B2(n45), .ZN(N317) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[63]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n12), .A2(n92), .B1(n48), .B2(n47), .ZN(N318) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n76) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n88), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  INVD2BWP30P140 U135 ( .I(n76), .ZN(n91) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  INVD2BWP30P140 U147 ( .I(n76), .ZN(n88) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n88), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n88), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n88), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n88), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n88), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n88), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n88), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n88), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U156 ( .A1(n85), .A2(n88), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U157 ( .A1(n86), .A2(n88), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U158 ( .A1(n87), .A2(n88), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n88), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_35 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  NR2D1BWP30P140 U4 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INR2D1BWP30P140 U5 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  INVD1BWP30P140 U6 ( .I(n4), .ZN(n12) );
  INVD1BWP30P140 U7 ( .I(n12), .ZN(n1) );
  INVD1BWP30P140 U8 ( .I(n12), .ZN(n2) );
  BUFFD12BWP30P140 U9 ( .I(n46), .Z(n48) );
  CKND2D3BWP30P140 U10 ( .A1(n7), .A2(n6), .ZN(n46) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U14 ( .I(n12), .ZN(n42) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n12), .ZN(n49) );
  INVD1BWP30P140 U18 ( .I(n66), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n49), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD1BWP30P140 U24 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[39]), .ZN(n8) );
  OAI22D1BWP30P140 U26 ( .A1(n49), .A2(n57), .B1(n48), .B2(n8), .ZN(N294) );
  INVD1BWP30P140 U27 ( .I(i_data_bus[6]), .ZN(n60) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[38]), .ZN(n9) );
  OAI22D1BWP30P140 U29 ( .A1(n49), .A2(n60), .B1(n48), .B2(n9), .ZN(N293) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[37]), .ZN(n10) );
  OAI22D1BWP30P140 U32 ( .A1(n49), .A2(n59), .B1(n48), .B2(n10), .ZN(N292) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[4]), .ZN(n58) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[36]), .ZN(n11) );
  OAI22D1BWP30P140 U35 ( .A1(n49), .A2(n58), .B1(n48), .B2(n11), .ZN(N291) );
  INVD1BWP30P140 U36 ( .I(n12), .ZN(n17) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[3]), .ZN(n56) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[35]), .ZN(n13) );
  OAI22D1BWP30P140 U39 ( .A1(n1), .A2(n56), .B1(n48), .B2(n13), .ZN(N290) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[2]), .ZN(n61) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[34]), .ZN(n14) );
  OAI22D1BWP30P140 U42 ( .A1(n42), .A2(n61), .B1(n48), .B2(n14), .ZN(N289) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[1]), .ZN(n62) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[33]), .ZN(n15) );
  OAI22D1BWP30P140 U45 ( .A1(n17), .A2(n62), .B1(n48), .B2(n15), .ZN(N288) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[32]), .ZN(n16) );
  OAI22D1BWP30P140 U48 ( .A1(n2), .A2(n64), .B1(n46), .B2(n16), .ZN(N287) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[24]), .ZN(n74) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[56]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n17), .A2(n74), .B1(n48), .B2(n22), .ZN(N311) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[23]), .ZN(n75) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[55]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n2), .A2(n75), .B1(n48), .B2(n23), .ZN(N310) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[22]), .ZN(n76) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[54]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n1), .A2(n76), .B1(n48), .B2(n24), .ZN(N309) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[21]), .ZN(n77) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[53]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n42), .A2(n77), .B1(n48), .B2(n25), .ZN(N308) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[27]), .ZN(n71) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[59]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n17), .A2(n71), .B1(n48), .B2(n26), .ZN(N314) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[26]), .ZN(n72) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[58]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n2), .A2(n72), .B1(n48), .B2(n27), .ZN(N313) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[25]), .ZN(n73) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[57]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n1), .A2(n73), .B1(n48), .B2(n28), .ZN(N312) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[17]), .ZN(n82) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[49]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n49), .A2(n82), .B1(n48), .B2(n29), .ZN(N304) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[16]), .ZN(n83) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[48]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n1), .A2(n83), .B1(n48), .B2(n30), .ZN(N303) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[15]), .ZN(n84) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[47]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n42), .A2(n84), .B1(n48), .B2(n31), .ZN(N302) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[14]), .ZN(n85) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[46]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n17), .A2(n85), .B1(n48), .B2(n32), .ZN(N301) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[13]), .ZN(n86) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[45]), .ZN(n33) );
  OAI22D1BWP30P140 U87 ( .A1(n2), .A2(n86), .B1(n48), .B2(n33), .ZN(N300) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[12]), .ZN(n87) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[44]), .ZN(n34) );
  OAI22D1BWP30P140 U90 ( .A1(n1), .A2(n87), .B1(n48), .B2(n34), .ZN(N299) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[11]), .ZN(n89) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[43]), .ZN(n35) );
  OAI22D1BWP30P140 U93 ( .A1(n42), .A2(n89), .B1(n48), .B2(n35), .ZN(N298) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[10]), .ZN(n92) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[42]), .ZN(n36) );
  OAI22D1BWP30P140 U96 ( .A1(n17), .A2(n92), .B1(n48), .B2(n36), .ZN(N297) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[9]), .ZN(n65) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[41]), .ZN(n37) );
  OAI22D1BWP30P140 U99 ( .A1(n2), .A2(n65), .B1(n46), .B2(n37), .ZN(N296) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[8]), .ZN(n88) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[40]), .ZN(n38) );
  OAI22D1BWP30P140 U102 ( .A1(n1), .A2(n88), .B1(n48), .B2(n38), .ZN(N295) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[52]), .ZN(n39) );
  OAI22D1BWP30P140 U105 ( .A1(n42), .A2(n79), .B1(n48), .B2(n39), .ZN(N307) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[19]), .ZN(n80) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[51]), .ZN(n40) );
  OAI22D1BWP30P140 U108 ( .A1(n17), .A2(n80), .B1(n48), .B2(n40), .ZN(N306) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[18]), .ZN(n81) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[50]), .ZN(n41) );
  OAI22D1BWP30P140 U111 ( .A1(n42), .A2(n81), .B1(n48), .B2(n41), .ZN(N305) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[30]), .ZN(n68) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[62]), .ZN(n43) );
  OAI22D1BWP30P140 U114 ( .A1(n2), .A2(n68), .B1(n48), .B2(n43), .ZN(N317) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[31]), .ZN(n67) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[63]), .ZN(n44) );
  OAI22D1BWP30P140 U117 ( .A1(n1), .A2(n67), .B1(n48), .B2(n44), .ZN(N318) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[29]), .ZN(n69) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[61]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n42), .A2(n69), .B1(n48), .B2(n45), .ZN(N316) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[28]), .ZN(n70) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[60]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n17), .A2(n70), .B1(n48), .B2(n47), .ZN(N315) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n66) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n78), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  INVD2BWP30P140 U135 ( .I(n66), .ZN(n91) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  INVD2BWP30P140 U137 ( .I(n66), .ZN(n78) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n78), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n78), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n78), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n78), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n78), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n78), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n78), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n78), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n78), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n78), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n78), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n78), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_36 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  INVD1BWP30P140 U4 ( .I(n4), .ZN(n13) );
  NR2D1BWP30P140 U5 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  INVD1BWP30P140 U7 ( .I(n13), .ZN(n1) );
  INVD1BWP30P140 U8 ( .I(n13), .ZN(n2) );
  BUFFD12BWP30P140 U9 ( .I(n46), .Z(n48) );
  CKND2D3BWP30P140 U10 ( .A1(n7), .A2(n6), .ZN(n46) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U14 ( .I(n13), .ZN(n49) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n13), .ZN(n40) );
  INVD1BWP30P140 U18 ( .I(n78), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n40), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n13), .ZN(n12) );
  INVD1BWP30P140 U24 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U25 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[32]), .ZN(n8) );
  OAI22D1BWP30P140 U27 ( .A1(n2), .A2(n64), .B1(n48), .B2(n8), .ZN(N287) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[1]), .ZN(n62) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[33]), .ZN(n9) );
  OAI22D1BWP30P140 U30 ( .A1(n1), .A2(n62), .B1(n48), .B2(n9), .ZN(N288) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[2]), .ZN(n61) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[34]), .ZN(n10) );
  OAI22D1BWP30P140 U33 ( .A1(n49), .A2(n61), .B1(n48), .B2(n10), .ZN(N289) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[35]), .ZN(n11) );
  OAI22D1BWP30P140 U36 ( .A1(n12), .A2(n60), .B1(n48), .B2(n11), .ZN(N290) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[36]), .ZN(n14) );
  OAI22D1BWP30P140 U39 ( .A1(n40), .A2(n59), .B1(n48), .B2(n14), .ZN(N291) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[5]), .ZN(n58) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[37]), .ZN(n15) );
  OAI22D1BWP30P140 U42 ( .A1(n40), .A2(n58), .B1(n48), .B2(n15), .ZN(N292) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[6]), .ZN(n57) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[38]), .ZN(n16) );
  OAI22D1BWP30P140 U45 ( .A1(n40), .A2(n57), .B1(n48), .B2(n16), .ZN(N293) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[39]), .ZN(n17) );
  OAI22D1BWP30P140 U48 ( .A1(n40), .A2(n56), .B1(n46), .B2(n17), .ZN(N294) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[44]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n40), .A2(n86), .B1(n48), .B2(n22), .ZN(N299) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[8]), .ZN(n92) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[40]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n1), .A2(n92), .B1(n48), .B2(n23), .ZN(N295) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[9]), .ZN(n89) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[41]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n49), .A2(n89), .B1(n48), .B2(n24), .ZN(N296) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[42]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n12), .A2(n88), .B1(n48), .B2(n25), .ZN(N297) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[11]), .ZN(n87) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[43]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n2), .A2(n87), .B1(n48), .B2(n26), .ZN(N298) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[31]), .ZN(n65) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[63]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n12), .A2(n65), .B1(n48), .B2(n27), .ZN(N318) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[30]), .ZN(n66) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[62]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n2), .A2(n66), .B1(n48), .B2(n28), .ZN(N317) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[29]), .ZN(n67) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[61]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n1), .A2(n67), .B1(n48), .B2(n29), .ZN(N316) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[28]), .ZN(n68) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[60]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n49), .A2(n68), .B1(n48), .B2(n30), .ZN(N315) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[59]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n12), .A2(n69), .B1(n48), .B2(n31), .ZN(N314) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[26]), .ZN(n70) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[58]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n2), .A2(n70), .B1(n48), .B2(n32), .ZN(N313) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[25]), .ZN(n71) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[57]), .ZN(n33) );
  OAI22D1BWP30P140 U87 ( .A1(n1), .A2(n71), .B1(n48), .B2(n33), .ZN(N312) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[24]), .ZN(n72) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[56]), .ZN(n34) );
  OAI22D1BWP30P140 U90 ( .A1(n49), .A2(n72), .B1(n48), .B2(n34), .ZN(N311) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[23]), .ZN(n73) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[55]), .ZN(n35) );
  OAI22D1BWP30P140 U93 ( .A1(n12), .A2(n73), .B1(n46), .B2(n35), .ZN(N310) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[54]), .ZN(n36) );
  OAI22D1BWP30P140 U96 ( .A1(n2), .A2(n74), .B1(n48), .B2(n36), .ZN(N309) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[21]), .ZN(n75) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[53]), .ZN(n37) );
  OAI22D1BWP30P140 U99 ( .A1(n1), .A2(n75), .B1(n48), .B2(n37), .ZN(N308) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[52]), .ZN(n38) );
  OAI22D1BWP30P140 U102 ( .A1(n49), .A2(n77), .B1(n48), .B2(n38), .ZN(N307) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[19]), .ZN(n79) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[51]), .ZN(n39) );
  OAI22D1BWP30P140 U105 ( .A1(n12), .A2(n79), .B1(n48), .B2(n39), .ZN(N306) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[18]), .ZN(n80) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[50]), .ZN(n41) );
  OAI22D1BWP30P140 U108 ( .A1(n1), .A2(n80), .B1(n48), .B2(n41), .ZN(N305) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[17]), .ZN(n81) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[49]), .ZN(n42) );
  OAI22D1BWP30P140 U111 ( .A1(n49), .A2(n81), .B1(n48), .B2(n42), .ZN(N304) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[16]), .ZN(n82) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[48]), .ZN(n43) );
  OAI22D1BWP30P140 U114 ( .A1(n12), .A2(n82), .B1(n48), .B2(n43), .ZN(N303) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[15]), .ZN(n83) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[47]), .ZN(n44) );
  OAI22D1BWP30P140 U117 ( .A1(n2), .A2(n83), .B1(n48), .B2(n44), .ZN(N302) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[14]), .ZN(n84) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[46]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n1), .A2(n84), .B1(n48), .B2(n45), .ZN(N301) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[13]), .ZN(n85) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[45]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n49), .A2(n85), .B1(n48), .B2(n47), .ZN(N300) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n78) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  INVD2BWP30P140 U135 ( .I(n78), .ZN(n76) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_37 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  INVD1BWP30P140 U4 ( .I(n4), .ZN(n13) );
  NR2D1BWP30P140 U5 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  INVD1BWP30P140 U7 ( .I(n13), .ZN(n1) );
  INVD1BWP30P140 U8 ( .I(n13), .ZN(n2) );
  BUFFD12BWP30P140 U9 ( .I(n46), .Z(n48) );
  CKND2D3BWP30P140 U10 ( .A1(n7), .A2(n6), .ZN(n46) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U14 ( .I(n13), .ZN(n33) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n13), .ZN(n49) );
  INVD1BWP30P140 U18 ( .I(n78), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n49), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n13), .ZN(n12) );
  INVD1BWP30P140 U24 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U25 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[32]), .ZN(n8) );
  OAI22D1BWP30P140 U27 ( .A1(n2), .A2(n64), .B1(n48), .B2(n8), .ZN(N287) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[1]), .ZN(n62) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[33]), .ZN(n9) );
  OAI22D1BWP30P140 U30 ( .A1(n1), .A2(n62), .B1(n48), .B2(n9), .ZN(N288) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[2]), .ZN(n61) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[34]), .ZN(n10) );
  OAI22D1BWP30P140 U33 ( .A1(n33), .A2(n61), .B1(n48), .B2(n10), .ZN(N289) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[35]), .ZN(n11) );
  OAI22D1BWP30P140 U36 ( .A1(n12), .A2(n60), .B1(n48), .B2(n11), .ZN(N290) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[36]), .ZN(n14) );
  OAI22D1BWP30P140 U39 ( .A1(n49), .A2(n59), .B1(n48), .B2(n14), .ZN(N291) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[5]), .ZN(n58) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[37]), .ZN(n15) );
  OAI22D1BWP30P140 U42 ( .A1(n49), .A2(n58), .B1(n48), .B2(n15), .ZN(N292) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[6]), .ZN(n57) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[38]), .ZN(n16) );
  OAI22D1BWP30P140 U45 ( .A1(n49), .A2(n57), .B1(n48), .B2(n16), .ZN(N293) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[39]), .ZN(n17) );
  OAI22D1BWP30P140 U48 ( .A1(n49), .A2(n56), .B1(n46), .B2(n17), .ZN(N294) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[8]), .ZN(n92) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[40]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n49), .A2(n92), .B1(n48), .B2(n22), .ZN(N295) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[9]), .ZN(n89) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[41]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n1), .A2(n89), .B1(n48), .B2(n23), .ZN(N296) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[42]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n33), .A2(n88), .B1(n48), .B2(n24), .ZN(N297) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[11]), .ZN(n87) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[43]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n12), .A2(n87), .B1(n48), .B2(n25), .ZN(N298) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[44]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n2), .A2(n86), .B1(n48), .B2(n26), .ZN(N299) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[13]), .ZN(n85) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[45]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n1), .A2(n85), .B1(n48), .B2(n27), .ZN(N300) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[14]), .ZN(n84) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[46]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n33), .A2(n84), .B1(n48), .B2(n28), .ZN(N301) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[15]), .ZN(n83) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[47]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n12), .A2(n83), .B1(n48), .B2(n29), .ZN(N302) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[16]), .ZN(n82) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[48]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n2), .A2(n82), .B1(n46), .B2(n30), .ZN(N303) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[17]), .ZN(n81) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[49]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n1), .A2(n81), .B1(n48), .B2(n31), .ZN(N304) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[18]), .ZN(n80) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[50]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n33), .A2(n80), .B1(n48), .B2(n32), .ZN(N305) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[19]), .ZN(n79) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[51]), .ZN(n34) );
  OAI22D1BWP30P140 U87 ( .A1(n12), .A2(n79), .B1(n48), .B2(n34), .ZN(N306) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[52]), .ZN(n35) );
  OAI22D1BWP30P140 U90 ( .A1(n2), .A2(n77), .B1(n48), .B2(n35), .ZN(N307) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[21]), .ZN(n75) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[53]), .ZN(n36) );
  OAI22D1BWP30P140 U93 ( .A1(n1), .A2(n75), .B1(n48), .B2(n36), .ZN(N308) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[54]), .ZN(n37) );
  OAI22D1BWP30P140 U96 ( .A1(n33), .A2(n74), .B1(n48), .B2(n37), .ZN(N309) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[23]), .ZN(n73) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[55]), .ZN(n38) );
  OAI22D1BWP30P140 U99 ( .A1(n12), .A2(n73), .B1(n48), .B2(n38), .ZN(N310) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[24]), .ZN(n72) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[56]), .ZN(n39) );
  OAI22D1BWP30P140 U102 ( .A1(n2), .A2(n72), .B1(n48), .B2(n39), .ZN(N311) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[25]), .ZN(n71) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[57]), .ZN(n40) );
  OAI22D1BWP30P140 U105 ( .A1(n1), .A2(n71), .B1(n48), .B2(n40), .ZN(N312) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[26]), .ZN(n70) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[58]), .ZN(n41) );
  OAI22D1BWP30P140 U108 ( .A1(n33), .A2(n70), .B1(n48), .B2(n41), .ZN(N313) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[59]), .ZN(n42) );
  OAI22D1BWP30P140 U111 ( .A1(n12), .A2(n69), .B1(n48), .B2(n42), .ZN(N314) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[28]), .ZN(n68) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[60]), .ZN(n43) );
  OAI22D1BWP30P140 U114 ( .A1(n2), .A2(n68), .B1(n48), .B2(n43), .ZN(N315) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[29]), .ZN(n67) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[61]), .ZN(n44) );
  OAI22D1BWP30P140 U117 ( .A1(n1), .A2(n67), .B1(n48), .B2(n44), .ZN(N316) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[30]), .ZN(n66) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[62]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n33), .A2(n66), .B1(n48), .B2(n45), .ZN(N317) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[31]), .ZN(n65) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[63]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n12), .A2(n65), .B1(n48), .B2(n47), .ZN(N318) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n78) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  INVD2BWP30P140 U135 ( .I(n78), .ZN(n76) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_38 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  INVD1BWP30P140 U4 ( .I(n4), .ZN(n13) );
  NR2D1BWP30P140 U5 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  INVD1BWP30P140 U7 ( .I(n13), .ZN(n1) );
  INVD1BWP30P140 U8 ( .I(n13), .ZN(n2) );
  BUFFD12BWP30P140 U9 ( .I(n46), .Z(n48) );
  CKND2D3BWP30P140 U10 ( .A1(n7), .A2(n6), .ZN(n46) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U14 ( .I(n13), .ZN(n33) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n13), .ZN(n49) );
  INVD1BWP30P140 U18 ( .I(n78), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n49), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n13), .ZN(n12) );
  INVD1BWP30P140 U24 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U25 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[32]), .ZN(n8) );
  OAI22D1BWP30P140 U27 ( .A1(n2), .A2(n64), .B1(n48), .B2(n8), .ZN(N287) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[1]), .ZN(n62) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[33]), .ZN(n9) );
  OAI22D1BWP30P140 U30 ( .A1(n1), .A2(n62), .B1(n48), .B2(n9), .ZN(N288) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[2]), .ZN(n61) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[34]), .ZN(n10) );
  OAI22D1BWP30P140 U33 ( .A1(n33), .A2(n61), .B1(n48), .B2(n10), .ZN(N289) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[35]), .ZN(n11) );
  OAI22D1BWP30P140 U36 ( .A1(n12), .A2(n60), .B1(n48), .B2(n11), .ZN(N290) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[36]), .ZN(n14) );
  OAI22D1BWP30P140 U39 ( .A1(n49), .A2(n59), .B1(n48), .B2(n14), .ZN(N291) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[5]), .ZN(n58) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[37]), .ZN(n15) );
  OAI22D1BWP30P140 U42 ( .A1(n49), .A2(n58), .B1(n48), .B2(n15), .ZN(N292) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[6]), .ZN(n57) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[38]), .ZN(n16) );
  OAI22D1BWP30P140 U45 ( .A1(n49), .A2(n57), .B1(n48), .B2(n16), .ZN(N293) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[39]), .ZN(n17) );
  OAI22D1BWP30P140 U48 ( .A1(n49), .A2(n56), .B1(n46), .B2(n17), .ZN(N294) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[8]), .ZN(n92) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[40]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n49), .A2(n92), .B1(n48), .B2(n22), .ZN(N295) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[9]), .ZN(n89) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[41]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n1), .A2(n89), .B1(n48), .B2(n23), .ZN(N296) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[42]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n33), .A2(n88), .B1(n48), .B2(n24), .ZN(N297) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[11]), .ZN(n87) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[43]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n12), .A2(n87), .B1(n48), .B2(n25), .ZN(N298) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[44]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n2), .A2(n86), .B1(n48), .B2(n26), .ZN(N299) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[13]), .ZN(n85) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[45]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n1), .A2(n85), .B1(n48), .B2(n27), .ZN(N300) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[14]), .ZN(n84) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[46]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n33), .A2(n84), .B1(n48), .B2(n28), .ZN(N301) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[15]), .ZN(n83) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[47]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n12), .A2(n83), .B1(n48), .B2(n29), .ZN(N302) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[16]), .ZN(n82) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[48]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n2), .A2(n82), .B1(n46), .B2(n30), .ZN(N303) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[17]), .ZN(n81) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[49]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n1), .A2(n81), .B1(n48), .B2(n31), .ZN(N304) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[18]), .ZN(n80) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[50]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n33), .A2(n80), .B1(n48), .B2(n32), .ZN(N305) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[19]), .ZN(n79) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[51]), .ZN(n34) );
  OAI22D1BWP30P140 U87 ( .A1(n12), .A2(n79), .B1(n48), .B2(n34), .ZN(N306) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[52]), .ZN(n35) );
  OAI22D1BWP30P140 U90 ( .A1(n2), .A2(n77), .B1(n48), .B2(n35), .ZN(N307) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[21]), .ZN(n75) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[53]), .ZN(n36) );
  OAI22D1BWP30P140 U93 ( .A1(n1), .A2(n75), .B1(n48), .B2(n36), .ZN(N308) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[54]), .ZN(n37) );
  OAI22D1BWP30P140 U96 ( .A1(n33), .A2(n74), .B1(n48), .B2(n37), .ZN(N309) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[23]), .ZN(n73) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[55]), .ZN(n38) );
  OAI22D1BWP30P140 U99 ( .A1(n12), .A2(n73), .B1(n48), .B2(n38), .ZN(N310) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[24]), .ZN(n72) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[56]), .ZN(n39) );
  OAI22D1BWP30P140 U102 ( .A1(n2), .A2(n72), .B1(n48), .B2(n39), .ZN(N311) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[25]), .ZN(n71) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[57]), .ZN(n40) );
  OAI22D1BWP30P140 U105 ( .A1(n1), .A2(n71), .B1(n48), .B2(n40), .ZN(N312) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[26]), .ZN(n70) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[58]), .ZN(n41) );
  OAI22D1BWP30P140 U108 ( .A1(n33), .A2(n70), .B1(n48), .B2(n41), .ZN(N313) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[59]), .ZN(n42) );
  OAI22D1BWP30P140 U111 ( .A1(n12), .A2(n69), .B1(n48), .B2(n42), .ZN(N314) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[28]), .ZN(n68) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[60]), .ZN(n43) );
  OAI22D1BWP30P140 U114 ( .A1(n2), .A2(n68), .B1(n48), .B2(n43), .ZN(N315) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[29]), .ZN(n67) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[61]), .ZN(n44) );
  OAI22D1BWP30P140 U117 ( .A1(n1), .A2(n67), .B1(n48), .B2(n44), .ZN(N316) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[30]), .ZN(n66) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[62]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n33), .A2(n66), .B1(n48), .B2(n45), .ZN(N317) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[31]), .ZN(n65) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[63]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n12), .A2(n65), .B1(n48), .B2(n47), .ZN(N318) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n78) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  INVD2BWP30P140 U135 ( .I(n78), .ZN(n76) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_39 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  INVD1BWP30P140 U4 ( .I(n4), .ZN(n13) );
  INR2D1BWP30P140 U5 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  NR2D1BWP30P140 U6 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INVD1BWP30P140 U7 ( .I(n13), .ZN(n1) );
  INVD1BWP30P140 U8 ( .I(n13), .ZN(n2) );
  BUFFD12BWP30P140 U9 ( .I(n46), .Z(n48) );
  CKND2D3BWP30P140 U10 ( .A1(n7), .A2(n6), .ZN(n46) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U14 ( .I(n13), .ZN(n33) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n13), .ZN(n49) );
  INVD1BWP30P140 U18 ( .I(n76), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n49), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n13), .ZN(n12) );
  INVD1BWP30P140 U24 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U25 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[32]), .ZN(n8) );
  OAI22D1BWP30P140 U27 ( .A1(n2), .A2(n64), .B1(n48), .B2(n8), .ZN(N287) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[1]), .ZN(n62) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[33]), .ZN(n9) );
  OAI22D1BWP30P140 U30 ( .A1(n1), .A2(n62), .B1(n48), .B2(n9), .ZN(N288) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[2]), .ZN(n61) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[34]), .ZN(n10) );
  OAI22D1BWP30P140 U33 ( .A1(n33), .A2(n61), .B1(n48), .B2(n10), .ZN(N289) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[35]), .ZN(n11) );
  OAI22D1BWP30P140 U36 ( .A1(n12), .A2(n60), .B1(n48), .B2(n11), .ZN(N290) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[36]), .ZN(n14) );
  OAI22D1BWP30P140 U39 ( .A1(n49), .A2(n59), .B1(n48), .B2(n14), .ZN(N291) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[5]), .ZN(n58) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[37]), .ZN(n15) );
  OAI22D1BWP30P140 U42 ( .A1(n49), .A2(n58), .B1(n48), .B2(n15), .ZN(N292) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[6]), .ZN(n57) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[38]), .ZN(n16) );
  OAI22D1BWP30P140 U45 ( .A1(n49), .A2(n57), .B1(n48), .B2(n16), .ZN(N293) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[39]), .ZN(n17) );
  OAI22D1BWP30P140 U48 ( .A1(n49), .A2(n56), .B1(n46), .B2(n17), .ZN(N294) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[8]), .ZN(n89) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[40]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n49), .A2(n89), .B1(n48), .B2(n22), .ZN(N295) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[9]), .ZN(n87) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[41]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n1), .A2(n87), .B1(n48), .B2(n23), .ZN(N296) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[10]), .ZN(n86) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[42]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n33), .A2(n86), .B1(n48), .B2(n24), .ZN(N297) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[11]), .ZN(n85) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[43]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n12), .A2(n85), .B1(n48), .B2(n25), .ZN(N298) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[12]), .ZN(n84) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[44]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n2), .A2(n84), .B1(n48), .B2(n26), .ZN(N299) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[13]), .ZN(n83) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[45]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n1), .A2(n83), .B1(n48), .B2(n27), .ZN(N300) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[14]), .ZN(n82) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[46]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n33), .A2(n82), .B1(n48), .B2(n28), .ZN(N301) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[15]), .ZN(n81) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[47]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n12), .A2(n81), .B1(n48), .B2(n29), .ZN(N302) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[16]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[48]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n2), .A2(n80), .B1(n46), .B2(n30), .ZN(N303) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[17]), .ZN(n79) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[49]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n1), .A2(n79), .B1(n48), .B2(n31), .ZN(N304) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[18]), .ZN(n78) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[50]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n33), .A2(n78), .B1(n48), .B2(n32), .ZN(N305) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[19]), .ZN(n77) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[51]), .ZN(n34) );
  OAI22D1BWP30P140 U87 ( .A1(n12), .A2(n77), .B1(n48), .B2(n34), .ZN(N306) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[20]), .ZN(n72) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[52]), .ZN(n35) );
  OAI22D1BWP30P140 U90 ( .A1(n2), .A2(n72), .B1(n48), .B2(n35), .ZN(N307) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[21]), .ZN(n71) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[53]), .ZN(n36) );
  OAI22D1BWP30P140 U93 ( .A1(n1), .A2(n71), .B1(n48), .B2(n36), .ZN(N308) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[22]), .ZN(n70) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[54]), .ZN(n37) );
  OAI22D1BWP30P140 U96 ( .A1(n33), .A2(n70), .B1(n48), .B2(n37), .ZN(N309) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[23]), .ZN(n69) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[55]), .ZN(n38) );
  OAI22D1BWP30P140 U99 ( .A1(n12), .A2(n69), .B1(n48), .B2(n38), .ZN(N310) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[24]), .ZN(n68) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[56]), .ZN(n39) );
  OAI22D1BWP30P140 U102 ( .A1(n2), .A2(n68), .B1(n48), .B2(n39), .ZN(N311) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[25]), .ZN(n67) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[57]), .ZN(n40) );
  OAI22D1BWP30P140 U105 ( .A1(n1), .A2(n67), .B1(n48), .B2(n40), .ZN(N312) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[26]), .ZN(n66) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[58]), .ZN(n41) );
  OAI22D1BWP30P140 U108 ( .A1(n33), .A2(n66), .B1(n48), .B2(n41), .ZN(N313) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[27]), .ZN(n65) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[59]), .ZN(n42) );
  OAI22D1BWP30P140 U111 ( .A1(n12), .A2(n65), .B1(n48), .B2(n42), .ZN(N314) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[28]), .ZN(n75) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[60]), .ZN(n43) );
  OAI22D1BWP30P140 U114 ( .A1(n2), .A2(n75), .B1(n48), .B2(n43), .ZN(N315) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[29]), .ZN(n74) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[61]), .ZN(n44) );
  OAI22D1BWP30P140 U117 ( .A1(n1), .A2(n74), .B1(n48), .B2(n44), .ZN(N316) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[30]), .ZN(n73) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[62]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n33), .A2(n73), .B1(n48), .B2(n45), .ZN(N317) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[63]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n12), .A2(n92), .B1(n48), .B2(n47), .ZN(N318) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n76) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n88), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  INVD2BWP30P140 U135 ( .I(n76), .ZN(n91) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  INVD2BWP30P140 U147 ( .I(n76), .ZN(n88) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n88), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n88), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n88), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n88), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n88), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n88), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n88), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n88), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U156 ( .A1(n85), .A2(n88), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U157 ( .A1(n86), .A2(n88), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U158 ( .A1(n87), .A2(n88), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n88), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_40 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  INVD1BWP30P140 U4 ( .I(n4), .ZN(n10) );
  NR2D1BWP30P140 U5 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  INVD1BWP30P140 U7 ( .I(n10), .ZN(n1) );
  INVD1BWP30P140 U8 ( .I(n10), .ZN(n2) );
  BUFFD12BWP30P140 U9 ( .I(n46), .Z(n48) );
  CKND2D3BWP30P140 U10 ( .A1(n7), .A2(n6), .ZN(n46) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U14 ( .I(n10), .ZN(n44) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n10), .ZN(n49) );
  INVD1BWP30P140 U18 ( .I(n70), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n49), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n10), .ZN(n17) );
  INVD1BWP30P140 U24 ( .I(i_data_bus[3]), .ZN(n59) );
  INVD1BWP30P140 U25 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[35]), .ZN(n8) );
  OAI22D1BWP30P140 U27 ( .A1(n1), .A2(n59), .B1(n48), .B2(n8), .ZN(N290) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[34]), .ZN(n9) );
  OAI22D1BWP30P140 U30 ( .A1(n44), .A2(n60), .B1(n48), .B2(n9), .ZN(N289) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[5]), .ZN(n57) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[37]), .ZN(n11) );
  OAI22D1BWP30P140 U33 ( .A1(n49), .A2(n57), .B1(n48), .B2(n11), .ZN(N292) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[6]), .ZN(n56) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[38]), .ZN(n12) );
  OAI22D1BWP30P140 U36 ( .A1(n49), .A2(n56), .B1(n48), .B2(n12), .ZN(N293) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[39]), .ZN(n13) );
  OAI22D1BWP30P140 U39 ( .A1(n49), .A2(n64), .B1(n48), .B2(n13), .ZN(N294) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[4]), .ZN(n58) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[36]), .ZN(n14) );
  OAI22D1BWP30P140 U42 ( .A1(n49), .A2(n58), .B1(n48), .B2(n14), .ZN(N291) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[1]), .ZN(n61) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[33]), .ZN(n15) );
  OAI22D1BWP30P140 U45 ( .A1(n17), .A2(n61), .B1(n48), .B2(n15), .ZN(N288) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[0]), .ZN(n62) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[32]), .ZN(n16) );
  OAI22D1BWP30P140 U48 ( .A1(n2), .A2(n62), .B1(n46), .B2(n16), .ZN(N287) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[9]), .ZN(n89) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[41]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n49), .A2(n89), .B1(n48), .B2(n22), .ZN(N296) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[42]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n1), .A2(n88), .B1(n48), .B2(n23), .ZN(N297) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[11]), .ZN(n87) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[43]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n44), .A2(n87), .B1(n48), .B2(n24), .ZN(N298) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[44]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n17), .A2(n86), .B1(n48), .B2(n25), .ZN(N299) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[13]), .ZN(n85) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[45]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n2), .A2(n85), .B1(n48), .B2(n26), .ZN(N300) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[14]), .ZN(n84) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[46]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n1), .A2(n84), .B1(n48), .B2(n27), .ZN(N301) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[15]), .ZN(n67) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[47]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n44), .A2(n67), .B1(n48), .B2(n28), .ZN(N302) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[16]), .ZN(n68) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[48]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n17), .A2(n68), .B1(n48), .B2(n29), .ZN(N303) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[17]), .ZN(n66) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[49]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n2), .A2(n66), .B1(n46), .B2(n30), .ZN(N304) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[18]), .ZN(n65) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[50]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n1), .A2(n65), .B1(n48), .B2(n31), .ZN(N305) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[19]), .ZN(n69) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[51]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n17), .A2(n69), .B1(n48), .B2(n32), .ZN(N306) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[20]), .ZN(n71) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[52]), .ZN(n33) );
  OAI22D1BWP30P140 U87 ( .A1(n2), .A2(n71), .B1(n48), .B2(n33), .ZN(N307) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[21]), .ZN(n72) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[53]), .ZN(n34) );
  OAI22D1BWP30P140 U90 ( .A1(n1), .A2(n72), .B1(n48), .B2(n34), .ZN(N308) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[22]), .ZN(n73) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[54]), .ZN(n35) );
  OAI22D1BWP30P140 U93 ( .A1(n44), .A2(n73), .B1(n48), .B2(n35), .ZN(N309) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[23]), .ZN(n74) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[55]), .ZN(n36) );
  OAI22D1BWP30P140 U96 ( .A1(n17), .A2(n74), .B1(n48), .B2(n36), .ZN(N310) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[24]), .ZN(n75) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[56]), .ZN(n37) );
  OAI22D1BWP30P140 U99 ( .A1(n2), .A2(n75), .B1(n48), .B2(n37), .ZN(N311) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[25]), .ZN(n76) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[57]), .ZN(n38) );
  OAI22D1BWP30P140 U102 ( .A1(n1), .A2(n76), .B1(n48), .B2(n38), .ZN(N312) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[26]), .ZN(n77) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[58]), .ZN(n39) );
  OAI22D1BWP30P140 U105 ( .A1(n44), .A2(n77), .B1(n48), .B2(n39), .ZN(N313) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[27]), .ZN(n78) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[59]), .ZN(n40) );
  OAI22D1BWP30P140 U108 ( .A1(n17), .A2(n78), .B1(n48), .B2(n40), .ZN(N314) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[28]), .ZN(n79) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[60]), .ZN(n41) );
  OAI22D1BWP30P140 U111 ( .A1(n2), .A2(n79), .B1(n48), .B2(n41), .ZN(N315) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[29]), .ZN(n80) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[61]), .ZN(n42) );
  OAI22D1BWP30P140 U114 ( .A1(n1), .A2(n80), .B1(n48), .B2(n42), .ZN(N316) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[8]), .ZN(n92) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[40]), .ZN(n43) );
  OAI22D1BWP30P140 U117 ( .A1(n44), .A2(n92), .B1(n48), .B2(n43), .ZN(N295) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[30]), .ZN(n81) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[62]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n44), .A2(n81), .B1(n48), .B2(n45), .ZN(N317) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[31]), .ZN(n83) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[63]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n17), .A2(n83), .B1(n48), .B2(n47), .ZN(N318) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n70) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n82), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  INVD2BWP30P140 U135 ( .I(n70), .ZN(n91) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U141 ( .I(n70), .ZN(n82) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n82), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n82), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n82), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n82), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n82), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n82), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n82), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n82), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n82), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n82), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n82), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n82), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_41 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n58), .ZN(n66) );
  CKAN2D1BWP30P140 U4 ( .A1(n4), .A2(n13), .Z(n2) );
  INR2D1BWP30P140 U5 ( .A1(i_valid[0]), .B1(n14), .ZN(n4) );
  NR2D1BWP30P140 U6 ( .A1(n14), .A2(n13), .ZN(n18) );
  CKND2D3BWP30P140 U7 ( .A1(n10), .A2(n9), .ZN(n58) );
  INVD4BWP30P140 U8 ( .I(n2), .ZN(n1) );
  INVD6BWP30P140 U9 ( .I(n66), .ZN(n80) );
  BUFFD4BWP30P140 U10 ( .I(n58), .Z(n93) );
  NR2D1BWP30P140 U11 ( .A1(n14), .A2(i_cmd[1]), .ZN(n9) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n14) );
  INVD2BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n13) );
  INVD1BWP30P140 U14 ( .I(n42), .ZN(n28) );
  INVD1BWP30P140 U15 ( .I(n85), .ZN(n7) );
  ND2D1BWP30P140 U16 ( .A1(n12), .A2(n11), .ZN(N325) );
  ND2D1BWP30P140 U17 ( .A1(n66), .A2(i_data_bus[6]), .ZN(n12) );
  ND2D1BWP30P140 U18 ( .A1(n85), .A2(i_data_bus[38]), .ZN(n11) );
  INVD1BWP30P140 U19 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U20 ( .I(i_valid[1]), .ZN(n15) );
  OAI31D1BWP30P140 U21 ( .A1(n14), .A2(n15), .A3(n13), .B(n1), .ZN(N353) );
  INVD1BWP30P140 U22 ( .I(n4), .ZN(n8) );
  INVD1BWP30P140 U23 ( .I(n14), .ZN(n5) );
  CKND2D2BWP30P140 U24 ( .A1(i_cmd[1]), .A2(n5), .ZN(n6) );
  INR2D2BWP30P140 U25 ( .A1(i_valid[1]), .B1(n6), .ZN(n92) );
  BUFFD8BWP30P140 U26 ( .I(n92), .Z(n85) );
  OAI21D1BWP30P140 U27 ( .A1(n8), .A2(i_cmd[1]), .B(n7), .ZN(N354) );
  INVD1BWP30P140 U28 ( .I(i_valid[0]), .ZN(n16) );
  MUX2NUD1BWP30P140 U29 ( .I0(n16), .I1(n15), .S(i_cmd[0]), .ZN(n10) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[0]), .ZN(n87) );
  MUX2NUD1BWP30P140 U31 ( .I0(n16), .I1(n15), .S(i_cmd[1]), .ZN(n17) );
  ND2OPTIBD1BWP30P140 U32 ( .A1(n18), .A2(n17), .ZN(n19) );
  INVD2BWP30P140 U33 ( .I(n19), .ZN(n42) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[32]), .ZN(n20) );
  OAI22D1BWP30P140 U35 ( .A1(n1), .A2(n87), .B1(n28), .B2(n20), .ZN(N287) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[4]), .ZN(n91) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[36]), .ZN(n21) );
  OAI22D1BWP30P140 U38 ( .A1(n1), .A2(n91), .B1(n28), .B2(n21), .ZN(N291) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[6]), .ZN(n23) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[38]), .ZN(n22) );
  OAI22D1BWP30P140 U41 ( .A1(n1), .A2(n23), .B1(n28), .B2(n22), .ZN(N293) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[5]), .ZN(n94) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[37]), .ZN(n24) );
  OAI22D1BWP30P140 U44 ( .A1(n1), .A2(n94), .B1(n28), .B2(n24), .ZN(N292) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[1]), .ZN(n88) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[33]), .ZN(n25) );
  OAI22D1BWP30P140 U47 ( .A1(n1), .A2(n88), .B1(n28), .B2(n25), .ZN(N288) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[3]), .ZN(n90) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[35]), .ZN(n26) );
  OAI22D1BWP30P140 U50 ( .A1(n1), .A2(n90), .B1(n28), .B2(n26), .ZN(N290) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[2]), .ZN(n89) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[34]), .ZN(n27) );
  OAI22D1BWP30P140 U53 ( .A1(n1), .A2(n89), .B1(n55), .B2(n27), .ZN(N289) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[7]), .ZN(n61) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[39]), .ZN(n59) );
  OAI22D1BWP30P140 U56 ( .A1(n1), .A2(n61), .B1(n41), .B2(n59), .ZN(N294) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[8]), .ZN(n71) );
  INVD2BWP30P140 U58 ( .I(n42), .ZN(n41) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[40]), .ZN(n29) );
  OAI22D1BWP30P140 U60 ( .A1(n1), .A2(n71), .B1(n55), .B2(n29), .ZN(N295) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[9]), .ZN(n76) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[41]), .ZN(n30) );
  OAI22D1BWP30P140 U63 ( .A1(n1), .A2(n76), .B1(n41), .B2(n30), .ZN(N296) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[10]), .ZN(n75) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[42]), .ZN(n31) );
  OAI22D1BWP30P140 U66 ( .A1(n1), .A2(n75), .B1(n55), .B2(n31), .ZN(N297) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[43]), .ZN(n32) );
  OAI22D1BWP30P140 U69 ( .A1(n1), .A2(n68), .B1(n41), .B2(n32), .ZN(N298) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[12]), .ZN(n67) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[44]), .ZN(n33) );
  OAI22D1BWP30P140 U72 ( .A1(n1), .A2(n67), .B1(n55), .B2(n33), .ZN(N299) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[13]), .ZN(n72) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[45]), .ZN(n34) );
  OAI22D1BWP30P140 U75 ( .A1(n1), .A2(n72), .B1(n41), .B2(n34), .ZN(N300) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[14]), .ZN(n86) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[46]), .ZN(n35) );
  OAI22D1BWP30P140 U78 ( .A1(n1), .A2(n86), .B1(n55), .B2(n35), .ZN(N301) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[15]), .ZN(n79) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[47]), .ZN(n36) );
  OAI22D1BWP30P140 U81 ( .A1(n1), .A2(n79), .B1(n41), .B2(n36), .ZN(N302) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[16]), .ZN(n84) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[48]), .ZN(n37) );
  OAI22D1BWP30P140 U84 ( .A1(n1), .A2(n84), .B1(n55), .B2(n37), .ZN(N303) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[17]), .ZN(n77) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[49]), .ZN(n38) );
  OAI22D1BWP30P140 U87 ( .A1(n1), .A2(n77), .B1(n41), .B2(n38), .ZN(N304) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[18]), .ZN(n83) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[50]), .ZN(n39) );
  OAI22D1BWP30P140 U90 ( .A1(n1), .A2(n83), .B1(n55), .B2(n39), .ZN(N305) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[19]), .ZN(n82) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[51]), .ZN(n40) );
  OAI22D1BWP30P140 U93 ( .A1(n1), .A2(n82), .B1(n41), .B2(n40), .ZN(N306) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[20]), .ZN(n74) );
  INVD2BWP30P140 U95 ( .I(n42), .ZN(n55) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[52]), .ZN(n43) );
  OAI22D1BWP30P140 U97 ( .A1(n1), .A2(n74), .B1(n55), .B2(n43), .ZN(N307) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[21]), .ZN(n73) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[53]), .ZN(n44) );
  OAI22D1BWP30P140 U100 ( .A1(n1), .A2(n73), .B1(n41), .B2(n44), .ZN(N308) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[22]), .ZN(n78) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[54]), .ZN(n45) );
  OAI22D1BWP30P140 U103 ( .A1(n1), .A2(n78), .B1(n55), .B2(n45), .ZN(N309) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[23]), .ZN(n63) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[55]), .ZN(n46) );
  OAI22D1BWP30P140 U106 ( .A1(n1), .A2(n63), .B1(n41), .B2(n46), .ZN(N310) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[24]), .ZN(n62) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[56]), .ZN(n47) );
  OAI22D1BWP30P140 U109 ( .A1(n1), .A2(n62), .B1(n55), .B2(n47), .ZN(N311) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[25]), .ZN(n56) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[57]), .ZN(n48) );
  OAI22D1BWP30P140 U112 ( .A1(n1), .A2(n56), .B1(n41), .B2(n48), .ZN(N312) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[26]), .ZN(n65) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[58]), .ZN(n49) );
  OAI22D1BWP30P140 U115 ( .A1(n1), .A2(n65), .B1(n55), .B2(n49), .ZN(N313) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[27]), .ZN(n64) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[59]), .ZN(n50) );
  OAI22D1BWP30P140 U118 ( .A1(n1), .A2(n64), .B1(n41), .B2(n50), .ZN(N314) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[28]), .ZN(n70) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[60]), .ZN(n51) );
  OAI22D1BWP30P140 U121 ( .A1(n1), .A2(n70), .B1(n55), .B2(n51), .ZN(N315) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[29]), .ZN(n57) );
  INVD1BWP30P140 U123 ( .I(i_data_bus[61]), .ZN(n52) );
  OAI22D1BWP30P140 U124 ( .A1(n1), .A2(n57), .B1(n41), .B2(n52), .ZN(N316) );
  INVD1BWP30P140 U125 ( .I(i_data_bus[30]), .ZN(n69) );
  INVD1BWP30P140 U126 ( .I(i_data_bus[62]), .ZN(n53) );
  OAI22D1BWP30P140 U127 ( .A1(n1), .A2(n69), .B1(n55), .B2(n53), .ZN(N317) );
  INVD1BWP30P140 U128 ( .I(i_data_bus[31]), .ZN(n81) );
  INVD1BWP30P140 U129 ( .I(i_data_bus[63]), .ZN(n54) );
  OAI22D1BWP30P140 U130 ( .A1(n1), .A2(n81), .B1(n41), .B2(n54), .ZN(N318) );
  MOAI22D1BWP30P140 U131 ( .A1(n56), .A2(n80), .B1(i_data_bus[57]), .B2(n92), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U132 ( .A1(n57), .A2(n80), .B1(i_data_bus[61]), .B2(n85), 
        .ZN(N348) );
  INVD2BWP30P140 U133 ( .I(n85), .ZN(n60) );
  OAI22D1BWP30P140 U134 ( .A1(n93), .A2(n61), .B1(n60), .B2(n59), .ZN(N326) );
  MOAI22D1BWP30P140 U135 ( .A1(n62), .A2(n80), .B1(i_data_bus[56]), .B2(n85), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U136 ( .A1(n63), .A2(n80), .B1(i_data_bus[55]), .B2(n85), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U137 ( .A1(n64), .A2(n80), .B1(i_data_bus[59]), .B2(n85), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U138 ( .A1(n65), .A2(n80), .B1(i_data_bus[58]), .B2(n85), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U139 ( .A1(n67), .A2(n80), .B1(i_data_bus[44]), .B2(n92), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U140 ( .A1(n68), .A2(n80), .B1(i_data_bus[43]), .B2(n85), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U141 ( .A1(n69), .A2(n80), .B1(i_data_bus[62]), .B2(n85), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U142 ( .A1(n70), .A2(n80), .B1(i_data_bus[60]), .B2(n85), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U143 ( .A1(n71), .A2(n80), .B1(i_data_bus[40]), .B2(n85), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U144 ( .A1(n72), .A2(n80), .B1(i_data_bus[45]), .B2(n85), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U145 ( .A1(n73), .A2(n80), .B1(i_data_bus[53]), .B2(n85), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U146 ( .A1(n74), .A2(n80), .B1(i_data_bus[52]), .B2(n85), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U147 ( .A1(n75), .A2(n93), .B1(i_data_bus[42]), .B2(n85), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U148 ( .A1(n76), .A2(n80), .B1(i_data_bus[41]), .B2(n85), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U149 ( .A1(n77), .A2(n80), .B1(i_data_bus[49]), .B2(n85), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U150 ( .A1(n78), .A2(n80), .B1(i_data_bus[54]), .B2(n85), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U151 ( .A1(n79), .A2(n58), .B1(i_data_bus[47]), .B2(n85), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n80), .B1(i_data_bus[63]), .B2(n85), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n58), .B1(i_data_bus[51]), .B2(n85), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n58), .B1(i_data_bus[50]), .B2(n85), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n58), .B1(i_data_bus[48]), .B2(n85), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n58), .B1(i_data_bus[46]), .B2(n85), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n93), .B1(i_data_bus[32]), .B2(n92), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n93), .B1(i_data_bus[33]), .B2(n92), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n93), .B1(i_data_bus[34]), .B2(n92), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n93), .B1(i_data_bus[35]), .B2(n92), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U161 ( .A1(n91), .A2(n93), .B1(i_data_bus[36]), .B2(n92), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U162 ( .A1(n94), .A2(n93), .B1(i_data_bus[37]), .B2(n92), 
        .ZN(N324) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_42 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n58), .ZN(n73) );
  CKAN2D1BWP30P140 U4 ( .A1(n4), .A2(n13), .Z(n2) );
  INR2D1BWP30P140 U5 ( .A1(i_valid[0]), .B1(n14), .ZN(n4) );
  NR2D1BWP30P140 U6 ( .A1(n14), .A2(n13), .ZN(n18) );
  CKND2D3BWP30P140 U7 ( .A1(n10), .A2(n9), .ZN(n58) );
  INVD4BWP30P140 U8 ( .I(n2), .ZN(n1) );
  INVD6BWP30P140 U9 ( .I(n73), .ZN(n71) );
  BUFFD4BWP30P140 U10 ( .I(n58), .Z(n93) );
  NR2D1BWP30P140 U11 ( .A1(n14), .A2(i_cmd[1]), .ZN(n9) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n14) );
  INVD2BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n13) );
  INVD1BWP30P140 U14 ( .I(n40), .ZN(n27) );
  INVD1BWP30P140 U15 ( .I(n85), .ZN(n7) );
  ND2D1BWP30P140 U16 ( .A1(n12), .A2(n11), .ZN(N325) );
  ND2D1BWP30P140 U17 ( .A1(n73), .A2(i_data_bus[6]), .ZN(n12) );
  ND2D1BWP30P140 U18 ( .A1(n85), .A2(i_data_bus[38]), .ZN(n11) );
  INVD1BWP30P140 U19 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U20 ( .I(i_valid[1]), .ZN(n15) );
  OAI31D1BWP30P140 U21 ( .A1(n14), .A2(n15), .A3(n13), .B(n1), .ZN(N353) );
  INVD1BWP30P140 U22 ( .I(n4), .ZN(n8) );
  INVD1BWP30P140 U23 ( .I(n14), .ZN(n5) );
  CKND2D2BWP30P140 U24 ( .A1(i_cmd[1]), .A2(n5), .ZN(n6) );
  INR2D2BWP30P140 U25 ( .A1(i_valid[1]), .B1(n6), .ZN(n92) );
  BUFFD8BWP30P140 U26 ( .I(n92), .Z(n85) );
  OAI21D1BWP30P140 U27 ( .A1(n8), .A2(i_cmd[1]), .B(n7), .ZN(N354) );
  INVD1BWP30P140 U28 ( .I(i_valid[0]), .ZN(n16) );
  MUX2NUD1BWP30P140 U29 ( .I0(n16), .I1(n15), .S(i_cmd[0]), .ZN(n10) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[5]), .ZN(n94) );
  MUX2NUD1BWP30P140 U31 ( .I0(n16), .I1(n15), .S(i_cmd[1]), .ZN(n17) );
  ND2OPTIBD1BWP30P140 U32 ( .A1(n18), .A2(n17), .ZN(n19) );
  INVD2BWP30P140 U33 ( .I(n19), .ZN(n40) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[37]), .ZN(n20) );
  OAI22D1BWP30P140 U35 ( .A1(n1), .A2(n94), .B1(n27), .B2(n20), .ZN(N292) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[4]), .ZN(n91) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[36]), .ZN(n21) );
  OAI22D1BWP30P140 U38 ( .A1(n1), .A2(n91), .B1(n27), .B2(n21), .ZN(N291) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[3]), .ZN(n90) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[35]), .ZN(n22) );
  OAI22D1BWP30P140 U41 ( .A1(n1), .A2(n90), .B1(n27), .B2(n22), .ZN(N290) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[2]), .ZN(n89) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[34]), .ZN(n23) );
  OAI22D1BWP30P140 U44 ( .A1(n1), .A2(n89), .B1(n27), .B2(n23), .ZN(N289) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[1]), .ZN(n88) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[33]), .ZN(n24) );
  OAI22D1BWP30P140 U47 ( .A1(n1), .A2(n88), .B1(n27), .B2(n24), .ZN(N288) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[0]), .ZN(n87) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[32]), .ZN(n25) );
  OAI22D1BWP30P140 U50 ( .A1(n1), .A2(n87), .B1(n27), .B2(n25), .ZN(N287) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[7]), .ZN(n61) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[39]), .ZN(n59) );
  OAI22D1BWP30P140 U53 ( .A1(n1), .A2(n61), .B1(n55), .B2(n59), .ZN(N294) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[6]), .ZN(n28) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[38]), .ZN(n26) );
  OAI22D1BWP30P140 U56 ( .A1(n1), .A2(n28), .B1(n53), .B2(n26), .ZN(N293) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[10]), .ZN(n83) );
  INVD2BWP30P140 U58 ( .I(n40), .ZN(n53) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[42]), .ZN(n29) );
  OAI22D1BWP30P140 U60 ( .A1(n1), .A2(n83), .B1(n55), .B2(n29), .ZN(N297) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[11]), .ZN(n82) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[43]), .ZN(n30) );
  OAI22D1BWP30P140 U63 ( .A1(n1), .A2(n82), .B1(n53), .B2(n30), .ZN(N298) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[12]), .ZN(n81) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[44]), .ZN(n31) );
  OAI22D1BWP30P140 U66 ( .A1(n1), .A2(n81), .B1(n55), .B2(n31), .ZN(N299) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[13]), .ZN(n80) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[45]), .ZN(n32) );
  OAI22D1BWP30P140 U69 ( .A1(n1), .A2(n80), .B1(n53), .B2(n32), .ZN(N300) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[8]), .ZN(n86) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[40]), .ZN(n33) );
  OAI22D1BWP30P140 U72 ( .A1(n1), .A2(n86), .B1(n55), .B2(n33), .ZN(N295) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[9]), .ZN(n84) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[41]), .ZN(n34) );
  OAI22D1BWP30P140 U75 ( .A1(n1), .A2(n84), .B1(n53), .B2(n34), .ZN(N296) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[15]), .ZN(n78) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[47]), .ZN(n35) );
  OAI22D1BWP30P140 U78 ( .A1(n1), .A2(n78), .B1(n55), .B2(n35), .ZN(N302) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[14]), .ZN(n79) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[46]), .ZN(n36) );
  OAI22D1BWP30P140 U81 ( .A1(n1), .A2(n79), .B1(n53), .B2(n36), .ZN(N301) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[17]), .ZN(n76) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[49]), .ZN(n37) );
  OAI22D1BWP30P140 U84 ( .A1(n1), .A2(n76), .B1(n55), .B2(n37), .ZN(N304) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[50]), .ZN(n38) );
  OAI22D1BWP30P140 U87 ( .A1(n1), .A2(n75), .B1(n53), .B2(n38), .ZN(N305) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[19]), .ZN(n74) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[51]), .ZN(n39) );
  OAI22D1BWP30P140 U90 ( .A1(n1), .A2(n74), .B1(n55), .B2(n39), .ZN(N306) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[20]), .ZN(n72) );
  INVD2BWP30P140 U92 ( .I(n40), .ZN(n55) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[52]), .ZN(n41) );
  OAI22D1BWP30P140 U94 ( .A1(n1), .A2(n72), .B1(n55), .B2(n41), .ZN(N307) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[21]), .ZN(n70) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[53]), .ZN(n42) );
  OAI22D1BWP30P140 U97 ( .A1(n1), .A2(n70), .B1(n53), .B2(n42), .ZN(N308) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[22]), .ZN(n69) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[54]), .ZN(n43) );
  OAI22D1BWP30P140 U100 ( .A1(n1), .A2(n69), .B1(n55), .B2(n43), .ZN(N309) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[23]), .ZN(n68) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[55]), .ZN(n44) );
  OAI22D1BWP30P140 U103 ( .A1(n1), .A2(n68), .B1(n53), .B2(n44), .ZN(N310) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[24]), .ZN(n66) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[56]), .ZN(n45) );
  OAI22D1BWP30P140 U106 ( .A1(n1), .A2(n66), .B1(n55), .B2(n45), .ZN(N311) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[25]), .ZN(n56) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[57]), .ZN(n46) );
  OAI22D1BWP30P140 U109 ( .A1(n1), .A2(n56), .B1(n53), .B2(n46), .ZN(N312) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[26]), .ZN(n67) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[58]), .ZN(n47) );
  OAI22D1BWP30P140 U112 ( .A1(n1), .A2(n67), .B1(n55), .B2(n47), .ZN(N313) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[28]), .ZN(n64) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[60]), .ZN(n48) );
  OAI22D1BWP30P140 U115 ( .A1(n1), .A2(n64), .B1(n53), .B2(n48), .ZN(N315) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[29]), .ZN(n57) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[61]), .ZN(n49) );
  OAI22D1BWP30P140 U118 ( .A1(n1), .A2(n57), .B1(n55), .B2(n49), .ZN(N316) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[30]), .ZN(n63) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[62]), .ZN(n50) );
  OAI22D1BWP30P140 U121 ( .A1(n1), .A2(n63), .B1(n53), .B2(n50), .ZN(N317) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[31]), .ZN(n62) );
  INVD1BWP30P140 U123 ( .I(i_data_bus[63]), .ZN(n51) );
  OAI22D1BWP30P140 U124 ( .A1(n1), .A2(n62), .B1(n55), .B2(n51), .ZN(N318) );
  INVD1BWP30P140 U125 ( .I(i_data_bus[16]), .ZN(n77) );
  INVD1BWP30P140 U126 ( .I(i_data_bus[48]), .ZN(n52) );
  OAI22D1BWP30P140 U127 ( .A1(n1), .A2(n77), .B1(n53), .B2(n52), .ZN(N303) );
  INVD1BWP30P140 U128 ( .I(i_data_bus[27]), .ZN(n65) );
  INVD1BWP30P140 U129 ( .I(i_data_bus[59]), .ZN(n54) );
  OAI22D1BWP30P140 U130 ( .A1(n1), .A2(n65), .B1(n53), .B2(n54), .ZN(N314) );
  MOAI22D1BWP30P140 U131 ( .A1(n56), .A2(n71), .B1(i_data_bus[57]), .B2(n92), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U132 ( .A1(n57), .A2(n71), .B1(i_data_bus[61]), .B2(n85), 
        .ZN(N348) );
  INVD2BWP30P140 U133 ( .I(n85), .ZN(n60) );
  OAI22D1BWP30P140 U134 ( .A1(n93), .A2(n61), .B1(n60), .B2(n59), .ZN(N326) );
  MOAI22D1BWP30P140 U135 ( .A1(n62), .A2(n71), .B1(i_data_bus[63]), .B2(n85), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U136 ( .A1(n63), .A2(n71), .B1(i_data_bus[62]), .B2(n85), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U137 ( .A1(n64), .A2(n71), .B1(i_data_bus[60]), .B2(n85), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U138 ( .A1(n65), .A2(n71), .B1(i_data_bus[59]), .B2(n85), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U139 ( .A1(n66), .A2(n71), .B1(i_data_bus[56]), .B2(n92), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U140 ( .A1(n67), .A2(n71), .B1(i_data_bus[58]), .B2(n85), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U141 ( .A1(n68), .A2(n71), .B1(i_data_bus[55]), .B2(n85), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U142 ( .A1(n69), .A2(n71), .B1(i_data_bus[54]), .B2(n85), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U143 ( .A1(n70), .A2(n71), .B1(i_data_bus[53]), .B2(n85), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U144 ( .A1(n72), .A2(n71), .B1(i_data_bus[52]), .B2(n85), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n71), .B1(i_data_bus[51]), .B2(n85), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n71), .B1(i_data_bus[50]), .B2(n85), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n71), .B1(i_data_bus[49]), .B2(n85), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n71), .B1(i_data_bus[48]), .B2(n85), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n93), .B1(i_data_bus[47]), .B2(n85), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n71), .B1(i_data_bus[46]), .B2(n85), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n71), .B1(i_data_bus[45]), .B2(n85), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n58), .B1(i_data_bus[44]), .B2(n85), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n58), .B1(i_data_bus[43]), .B2(n85), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n58), .B1(i_data_bus[42]), .B2(n85), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n58), .B1(i_data_bus[41]), .B2(n85), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n58), .B1(i_data_bus[40]), .B2(n85), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n93), .B1(i_data_bus[32]), .B2(n92), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n93), .B1(i_data_bus[33]), .B2(n92), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n93), .B1(i_data_bus[34]), .B2(n92), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n93), .B1(i_data_bus[35]), .B2(n92), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U161 ( .A1(n91), .A2(n93), .B1(i_data_bus[36]), .B2(n92), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U162 ( .A1(n94), .A2(n93), .B1(i_data_bus[37]), .B2(n92), 
        .ZN(N324) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_43 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n58), .ZN(n62) );
  CKAN2D1BWP30P140 U4 ( .A1(n4), .A2(n13), .Z(n2) );
  INR2D1BWP30P140 U5 ( .A1(i_valid[0]), .B1(n14), .ZN(n4) );
  NR2D1BWP30P140 U6 ( .A1(n14), .A2(n13), .ZN(n18) );
  CKND2D3BWP30P140 U7 ( .A1(n10), .A2(n9), .ZN(n58) );
  INVD4BWP30P140 U8 ( .I(n2), .ZN(n1) );
  INVD6BWP30P140 U9 ( .I(n62), .ZN(n85) );
  BUFFD4BWP30P140 U10 ( .I(n58), .Z(n93) );
  NR2D1BWP30P140 U11 ( .A1(n14), .A2(i_cmd[1]), .ZN(n9) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n14) );
  INVD2BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n13) );
  INVD1BWP30P140 U14 ( .I(n42), .ZN(n28) );
  INVD1BWP30P140 U15 ( .I(n84), .ZN(n7) );
  ND2D1BWP30P140 U16 ( .A1(n12), .A2(n11), .ZN(N325) );
  ND2D1BWP30P140 U17 ( .A1(n62), .A2(i_data_bus[6]), .ZN(n12) );
  ND2D1BWP30P140 U18 ( .A1(n84), .A2(i_data_bus[38]), .ZN(n11) );
  INVD1BWP30P140 U19 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U20 ( .I(i_valid[1]), .ZN(n15) );
  OAI31D1BWP30P140 U21 ( .A1(n14), .A2(n15), .A3(n13), .B(n1), .ZN(N353) );
  INVD1BWP30P140 U22 ( .I(n4), .ZN(n8) );
  INVD1BWP30P140 U23 ( .I(n14), .ZN(n5) );
  CKND2D2BWP30P140 U24 ( .A1(i_cmd[1]), .A2(n5), .ZN(n6) );
  INR2D2BWP30P140 U25 ( .A1(i_valid[1]), .B1(n6), .ZN(n92) );
  BUFFD8BWP30P140 U26 ( .I(n92), .Z(n84) );
  OAI21D1BWP30P140 U27 ( .A1(n8), .A2(i_cmd[1]), .B(n7), .ZN(N354) );
  INVD1BWP30P140 U28 ( .I(i_valid[0]), .ZN(n16) );
  MUX2NUD1BWP30P140 U29 ( .I0(n16), .I1(n15), .S(i_cmd[0]), .ZN(n10) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[3]), .ZN(n90) );
  MUX2NUD1BWP30P140 U31 ( .I0(n16), .I1(n15), .S(i_cmd[1]), .ZN(n17) );
  ND2OPTIBD1BWP30P140 U32 ( .A1(n18), .A2(n17), .ZN(n19) );
  INVD2BWP30P140 U33 ( .I(n19), .ZN(n42) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[35]), .ZN(n20) );
  OAI22D1BWP30P140 U35 ( .A1(n1), .A2(n90), .B1(n28), .B2(n20), .ZN(N290) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[2]), .ZN(n89) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[34]), .ZN(n21) );
  OAI22D1BWP30P140 U38 ( .A1(n1), .A2(n89), .B1(n28), .B2(n21), .ZN(N289) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[5]), .ZN(n94) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[37]), .ZN(n22) );
  OAI22D1BWP30P140 U41 ( .A1(n1), .A2(n94), .B1(n28), .B2(n22), .ZN(N292) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[4]), .ZN(n91) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[36]), .ZN(n23) );
  OAI22D1BWP30P140 U44 ( .A1(n1), .A2(n91), .B1(n28), .B2(n23), .ZN(N291) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[1]), .ZN(n88) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[33]), .ZN(n24) );
  OAI22D1BWP30P140 U47 ( .A1(n1), .A2(n88), .B1(n28), .B2(n24), .ZN(N288) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[0]), .ZN(n87) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[32]), .ZN(n25) );
  OAI22D1BWP30P140 U50 ( .A1(n1), .A2(n87), .B1(n28), .B2(n25), .ZN(N287) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[6]), .ZN(n27) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[38]), .ZN(n26) );
  OAI22D1BWP30P140 U53 ( .A1(n1), .A2(n27), .B1(n41), .B2(n26), .ZN(N293) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[7]), .ZN(n61) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[39]), .ZN(n59) );
  OAI22D1BWP30P140 U56 ( .A1(n1), .A2(n61), .B1(n55), .B2(n59), .ZN(N294) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[31]), .ZN(n74) );
  INVD2BWP30P140 U58 ( .I(n42), .ZN(n41) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[63]), .ZN(n29) );
  OAI22D1BWP30P140 U60 ( .A1(n1), .A2(n74), .B1(n41), .B2(n29), .ZN(N318) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[30]), .ZN(n69) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[62]), .ZN(n30) );
  OAI22D1BWP30P140 U63 ( .A1(n1), .A2(n69), .B1(n55), .B2(n30), .ZN(N317) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[29]), .ZN(n57) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[61]), .ZN(n31) );
  OAI22D1BWP30P140 U66 ( .A1(n1), .A2(n57), .B1(n41), .B2(n31), .ZN(N316) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[28]), .ZN(n82) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[60]), .ZN(n32) );
  OAI22D1BWP30P140 U69 ( .A1(n1), .A2(n82), .B1(n55), .B2(n32), .ZN(N315) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[27]), .ZN(n83) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[59]), .ZN(n33) );
  OAI22D1BWP30P140 U72 ( .A1(n1), .A2(n83), .B1(n41), .B2(n33), .ZN(N314) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[26]), .ZN(n86) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[58]), .ZN(n34) );
  OAI22D1BWP30P140 U75 ( .A1(n1), .A2(n86), .B1(n55), .B2(n34), .ZN(N313) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[25]), .ZN(n56) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[57]), .ZN(n35) );
  OAI22D1BWP30P140 U78 ( .A1(n1), .A2(n56), .B1(n41), .B2(n35), .ZN(N312) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[24]), .ZN(n81) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[56]), .ZN(n36) );
  OAI22D1BWP30P140 U81 ( .A1(n1), .A2(n81), .B1(n55), .B2(n36), .ZN(N311) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[23]), .ZN(n76) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[55]), .ZN(n37) );
  OAI22D1BWP30P140 U84 ( .A1(n1), .A2(n76), .B1(n41), .B2(n37), .ZN(N310) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[22]), .ZN(n75) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[54]), .ZN(n38) );
  OAI22D1BWP30P140 U87 ( .A1(n1), .A2(n75), .B1(n55), .B2(n38), .ZN(N309) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[21]), .ZN(n68) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[53]), .ZN(n39) );
  OAI22D1BWP30P140 U90 ( .A1(n1), .A2(n68), .B1(n41), .B2(n39), .ZN(N308) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[20]), .ZN(n71) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[52]), .ZN(n40) );
  OAI22D1BWP30P140 U93 ( .A1(n1), .A2(n71), .B1(n55), .B2(n40), .ZN(N307) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[19]), .ZN(n72) );
  INVD2BWP30P140 U95 ( .I(n42), .ZN(n55) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[51]), .ZN(n43) );
  OAI22D1BWP30P140 U97 ( .A1(n1), .A2(n72), .B1(n41), .B2(n43), .ZN(N306) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[18]), .ZN(n73) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[50]), .ZN(n44) );
  OAI22D1BWP30P140 U100 ( .A1(n1), .A2(n73), .B1(n55), .B2(n44), .ZN(N305) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[17]), .ZN(n70) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[49]), .ZN(n45) );
  OAI22D1BWP30P140 U103 ( .A1(n1), .A2(n70), .B1(n41), .B2(n45), .ZN(N304) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[16]), .ZN(n63) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[48]), .ZN(n46) );
  OAI22D1BWP30P140 U106 ( .A1(n1), .A2(n63), .B1(n55), .B2(n46), .ZN(N303) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[15]), .ZN(n64) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[47]), .ZN(n47) );
  OAI22D1BWP30P140 U109 ( .A1(n1), .A2(n64), .B1(n41), .B2(n47), .ZN(N302) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[14]), .ZN(n66) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[46]), .ZN(n48) );
  OAI22D1BWP30P140 U112 ( .A1(n1), .A2(n66), .B1(n55), .B2(n48), .ZN(N301) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[13]), .ZN(n65) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[45]), .ZN(n49) );
  OAI22D1BWP30P140 U115 ( .A1(n1), .A2(n65), .B1(n41), .B2(n49), .ZN(N300) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[12]), .ZN(n67) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[44]), .ZN(n50) );
  OAI22D1BWP30P140 U118 ( .A1(n1), .A2(n67), .B1(n55), .B2(n50), .ZN(N299) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[11]), .ZN(n80) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[43]), .ZN(n51) );
  OAI22D1BWP30P140 U121 ( .A1(n1), .A2(n80), .B1(n41), .B2(n51), .ZN(N298) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[10]), .ZN(n79) );
  INVD1BWP30P140 U123 ( .I(i_data_bus[42]), .ZN(n52) );
  OAI22D1BWP30P140 U124 ( .A1(n1), .A2(n79), .B1(n55), .B2(n52), .ZN(N297) );
  INVD1BWP30P140 U125 ( .I(i_data_bus[9]), .ZN(n78) );
  INVD1BWP30P140 U126 ( .I(i_data_bus[41]), .ZN(n53) );
  OAI22D1BWP30P140 U127 ( .A1(n1), .A2(n78), .B1(n41), .B2(n53), .ZN(N296) );
  INVD1BWP30P140 U128 ( .I(i_data_bus[8]), .ZN(n77) );
  INVD1BWP30P140 U129 ( .I(i_data_bus[40]), .ZN(n54) );
  OAI22D1BWP30P140 U130 ( .A1(n1), .A2(n77), .B1(n55), .B2(n54), .ZN(N295) );
  MOAI22D1BWP30P140 U131 ( .A1(n56), .A2(n85), .B1(i_data_bus[57]), .B2(n92), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U132 ( .A1(n57), .A2(n85), .B1(i_data_bus[61]), .B2(n84), 
        .ZN(N348) );
  INVD2BWP30P140 U133 ( .I(n84), .ZN(n60) );
  OAI22D1BWP30P140 U134 ( .A1(n93), .A2(n61), .B1(n60), .B2(n59), .ZN(N326) );
  MOAI22D1BWP30P140 U135 ( .A1(n63), .A2(n85), .B1(i_data_bus[48]), .B2(n84), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U136 ( .A1(n64), .A2(n85), .B1(i_data_bus[47]), .B2(n84), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U137 ( .A1(n65), .A2(n85), .B1(i_data_bus[45]), .B2(n84), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U138 ( .A1(n66), .A2(n85), .B1(i_data_bus[46]), .B2(n84), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U139 ( .A1(n67), .A2(n93), .B1(i_data_bus[44]), .B2(n92), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U140 ( .A1(n68), .A2(n85), .B1(i_data_bus[53]), .B2(n84), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U141 ( .A1(n69), .A2(n85), .B1(i_data_bus[62]), .B2(n84), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U142 ( .A1(n70), .A2(n85), .B1(i_data_bus[49]), .B2(n84), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U143 ( .A1(n71), .A2(n85), .B1(i_data_bus[52]), .B2(n84), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U144 ( .A1(n72), .A2(n85), .B1(i_data_bus[51]), .B2(n84), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U145 ( .A1(n73), .A2(n58), .B1(i_data_bus[50]), .B2(n84), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U146 ( .A1(n74), .A2(n85), .B1(i_data_bus[63]), .B2(n84), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U147 ( .A1(n75), .A2(n85), .B1(i_data_bus[54]), .B2(n84), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U148 ( .A1(n76), .A2(n85), .B1(i_data_bus[55]), .B2(n84), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U149 ( .A1(n77), .A2(n58), .B1(i_data_bus[40]), .B2(n84), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U150 ( .A1(n78), .A2(n58), .B1(i_data_bus[41]), .B2(n84), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U151 ( .A1(n79), .A2(n58), .B1(i_data_bus[42]), .B2(n84), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U152 ( .A1(n80), .A2(n58), .B1(i_data_bus[43]), .B2(n84), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U153 ( .A1(n81), .A2(n85), .B1(i_data_bus[56]), .B2(n84), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n82), .A2(n85), .B1(i_data_bus[60]), .B2(n84), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U155 ( .A1(n83), .A2(n85), .B1(i_data_bus[59]), .B2(n84), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n85), .B1(i_data_bus[58]), .B2(n84), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n93), .B1(i_data_bus[32]), .B2(n92), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n93), .B1(i_data_bus[33]), .B2(n92), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n93), .B1(i_data_bus[34]), .B2(n92), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n93), .B1(i_data_bus[35]), .B2(n92), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U161 ( .A1(n91), .A2(n93), .B1(i_data_bus[36]), .B2(n92), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U162 ( .A1(n94), .A2(n93), .B1(i_data_bus[37]), .B2(n92), 
        .ZN(N324) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_44 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD4BWP30P140 U3 ( .I(n57), .ZN(n84) );
  BUFFD8BWP30P140 U4 ( .I(n91), .Z(n83) );
  CKAN2D1BWP30P140 U5 ( .A1(n9), .A2(n13), .Z(n3) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n14), .ZN(n9) );
  NR2D1BWP30P140 U7 ( .A1(n14), .A2(n13), .ZN(n18) );
  INVD2BWP30P140 U8 ( .I(n83), .ZN(n1) );
  CKND2D3BWP30P140 U9 ( .A1(n6), .A2(n5), .ZN(n60) );
  INVD4BWP30P140 U10 ( .I(n3), .ZN(n2) );
  INVD4BWP30P140 U11 ( .I(n60), .ZN(n57) );
  BUFFD4BWP30P140 U12 ( .I(n60), .Z(n92) );
  NR2D1BWP30P140 U13 ( .A1(n14), .A2(i_cmd[1]), .ZN(n5) );
  ND2D1BWP30P140 U14 ( .A1(n4), .A2(i_en), .ZN(n14) );
  INVD2BWP30P140 U15 ( .I(i_cmd[0]), .ZN(n13) );
  INVD1BWP30P140 U16 ( .I(n33), .ZN(n28) );
  ND2D1BWP30P140 U17 ( .A1(n12), .A2(n11), .ZN(N325) );
  ND2D1BWP30P140 U18 ( .A1(n57), .A2(i_data_bus[6]), .ZN(n12) );
  ND2D1BWP30P140 U19 ( .A1(n83), .A2(i_data_bus[38]), .ZN(n11) );
  MOAI22D1BWP30P140 U20 ( .A1(n49), .A2(n84), .B1(i_data_bus[50]), .B2(n83), 
        .ZN(N337) );
  INVD1BWP30P140 U21 ( .I(i_data_bus[18]), .ZN(n49) );
  INVD1BWP30P140 U22 ( .I(i_valid[0]), .ZN(n16) );
  INVD2BWP30P140 U23 ( .I(i_valid[1]), .ZN(n15) );
  MUX2NUD1BWP30P140 U24 ( .I0(n16), .I1(n15), .S(i_cmd[0]), .ZN(n6) );
  INVD1BWP30P140 U25 ( .I(rst), .ZN(n4) );
  INVD1BWP30P140 U26 ( .I(n14), .ZN(n7) );
  CKND2D2BWP30P140 U27 ( .A1(i_cmd[1]), .A2(n7), .ZN(n8) );
  INR2D2BWP30P140 U28 ( .A1(i_valid[1]), .B1(n8), .ZN(n91) );
  OAI31D1BWP30P140 U29 ( .A1(n14), .A2(n15), .A3(n13), .B(n2), .ZN(N353) );
  INVD1BWP30P140 U30 ( .I(n9), .ZN(n10) );
  OAI21D1BWP30P140 U31 ( .A1(n10), .A2(i_cmd[1]), .B(n1), .ZN(N354) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[0]), .ZN(n86) );
  MUX2NUD1BWP30P140 U33 ( .I0(n16), .I1(n15), .S(i_cmd[1]), .ZN(n17) );
  ND2OPTIBD1BWP30P140 U34 ( .A1(n18), .A2(n17), .ZN(n19) );
  INVD2BWP30P140 U35 ( .I(n19), .ZN(n33) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[32]), .ZN(n20) );
  OAI22D1BWP30P140 U37 ( .A1(n2), .A2(n86), .B1(n28), .B2(n20), .ZN(N287) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[6]), .ZN(n22) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[38]), .ZN(n21) );
  OAI22D1BWP30P140 U40 ( .A1(n2), .A2(n22), .B1(n28), .B2(n21), .ZN(N293) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[5]), .ZN(n93) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[37]), .ZN(n23) );
  OAI22D1BWP30P140 U43 ( .A1(n2), .A2(n93), .B1(n28), .B2(n23), .ZN(N292) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[4]), .ZN(n90) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[36]), .ZN(n24) );
  OAI22D1BWP30P140 U46 ( .A1(n2), .A2(n90), .B1(n28), .B2(n24), .ZN(N291) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[1]), .ZN(n87) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[33]), .ZN(n25) );
  OAI22D1BWP30P140 U49 ( .A1(n2), .A2(n87), .B1(n28), .B2(n25), .ZN(N288) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[7]), .ZN(n62) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[39]), .ZN(n61) );
  OAI22D1BWP30P140 U52 ( .A1(n2), .A2(n62), .B1(n28), .B2(n61), .ZN(N294) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[3]), .ZN(n89) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[35]), .ZN(n26) );
  OAI22D1BWP30P140 U55 ( .A1(n2), .A2(n89), .B1(n56), .B2(n26), .ZN(N290) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[2]), .ZN(n88) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[34]), .ZN(n27) );
  OAI22D1BWP30P140 U58 ( .A1(n2), .A2(n88), .B1(n54), .B2(n27), .ZN(N289) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[31]), .ZN(n85) );
  INVD2BWP30P140 U60 ( .I(n33), .ZN(n56) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[63]), .ZN(n29) );
  OAI22D1BWP30P140 U62 ( .A1(n2), .A2(n85), .B1(n56), .B2(n29), .ZN(N318) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[30]), .ZN(n81) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[62]), .ZN(n30) );
  OAI22D1BWP30P140 U65 ( .A1(n2), .A2(n81), .B1(n54), .B2(n30), .ZN(N317) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[23]), .ZN(n74) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[55]), .ZN(n31) );
  OAI22D1BWP30P140 U68 ( .A1(n2), .A2(n74), .B1(n56), .B2(n31), .ZN(N310) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[22]), .ZN(n73) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[54]), .ZN(n32) );
  OAI22D1BWP30P140 U71 ( .A1(n2), .A2(n73), .B1(n54), .B2(n32), .ZN(N309) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[9]), .ZN(n64) );
  INVD2BWP30P140 U73 ( .I(n33), .ZN(n54) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[41]), .ZN(n34) );
  OAI22D1BWP30P140 U75 ( .A1(n2), .A2(n64), .B1(n56), .B2(n34), .ZN(N296) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[8]), .ZN(n63) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[40]), .ZN(n35) );
  OAI22D1BWP30P140 U78 ( .A1(n2), .A2(n63), .B1(n54), .B2(n35), .ZN(N295) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[19]), .ZN(n70) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[51]), .ZN(n36) );
  OAI22D1BWP30P140 U81 ( .A1(n2), .A2(n70), .B1(n56), .B2(n36), .ZN(N306) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[27]), .ZN(n77) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[59]), .ZN(n37) );
  OAI22D1BWP30P140 U84 ( .A1(n2), .A2(n77), .B1(n56), .B2(n37), .ZN(N314) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[29]), .ZN(n58) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[61]), .ZN(n38) );
  OAI22D1BWP30P140 U87 ( .A1(n2), .A2(n58), .B1(n54), .B2(n38), .ZN(N316) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[25]), .ZN(n59) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[57]), .ZN(n39) );
  OAI22D1BWP30P140 U90 ( .A1(n2), .A2(n59), .B1(n56), .B2(n39), .ZN(N312) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[11]), .ZN(n66) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[43]), .ZN(n40) );
  OAI22D1BWP30P140 U93 ( .A1(n2), .A2(n66), .B1(n54), .B2(n40), .ZN(N298) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[12]), .ZN(n67) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[44]), .ZN(n41) );
  OAI22D1BWP30P140 U96 ( .A1(n2), .A2(n67), .B1(n56), .B2(n41), .ZN(N299) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[13]), .ZN(n79) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[45]), .ZN(n42) );
  OAI22D1BWP30P140 U99 ( .A1(n2), .A2(n79), .B1(n54), .B2(n42), .ZN(N300) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[16]), .ZN(n82) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[48]), .ZN(n43) );
  OAI22D1BWP30P140 U102 ( .A1(n2), .A2(n82), .B1(n56), .B2(n43), .ZN(N303) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[14]), .ZN(n80) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[46]), .ZN(n44) );
  OAI22D1BWP30P140 U105 ( .A1(n2), .A2(n80), .B1(n54), .B2(n44), .ZN(N301) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[28]), .ZN(n78) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[60]), .ZN(n45) );
  OAI22D1BWP30P140 U108 ( .A1(n2), .A2(n78), .B1(n54), .B2(n45), .ZN(N315) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[24]), .ZN(n75) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[56]), .ZN(n46) );
  OAI22D1BWP30P140 U111 ( .A1(n2), .A2(n75), .B1(n56), .B2(n46), .ZN(N311) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[17]), .ZN(n69) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[49]), .ZN(n47) );
  OAI22D1BWP30P140 U114 ( .A1(n2), .A2(n69), .B1(n56), .B2(n47), .ZN(N304) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[50]), .ZN(n48) );
  OAI22D1BWP30P140 U116 ( .A1(n2), .A2(n49), .B1(n54), .B2(n48), .ZN(N305) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[21]), .ZN(n72) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[53]), .ZN(n50) );
  OAI22D1BWP30P140 U119 ( .A1(n2), .A2(n72), .B1(n54), .B2(n50), .ZN(N308) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[10]), .ZN(n65) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[42]), .ZN(n51) );
  OAI22D1BWP30P140 U122 ( .A1(n2), .A2(n65), .B1(n56), .B2(n51), .ZN(N297) );
  INVD1BWP30P140 U123 ( .I(i_data_bus[20]), .ZN(n71) );
  INVD1BWP30P140 U124 ( .I(i_data_bus[52]), .ZN(n52) );
  OAI22D1BWP30P140 U125 ( .A1(n2), .A2(n71), .B1(n56), .B2(n52), .ZN(N307) );
  INVD1BWP30P140 U126 ( .I(i_data_bus[15]), .ZN(n68) );
  INVD1BWP30P140 U127 ( .I(i_data_bus[47]), .ZN(n53) );
  OAI22D1BWP30P140 U128 ( .A1(n2), .A2(n68), .B1(n54), .B2(n53), .ZN(N302) );
  INVD1BWP30P140 U129 ( .I(i_data_bus[26]), .ZN(n76) );
  INVD1BWP30P140 U130 ( .I(i_data_bus[58]), .ZN(n55) );
  OAI22D1BWP30P140 U131 ( .A1(n2), .A2(n76), .B1(n54), .B2(n55), .ZN(N313) );
  MOAI22D1BWP30P140 U132 ( .A1(n58), .A2(n84), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U133 ( .A1(n59), .A2(n84), .B1(i_data_bus[57]), .B2(n83), 
        .ZN(N344) );
  OAI22D1BWP30P140 U134 ( .A1(n92), .A2(n62), .B1(n1), .B2(n61), .ZN(N326) );
  MOAI22D1BWP30P140 U135 ( .A1(n63), .A2(n84), .B1(i_data_bus[40]), .B2(n83), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U136 ( .A1(n64), .A2(n84), .B1(i_data_bus[41]), .B2(n83), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U137 ( .A1(n65), .A2(n84), .B1(i_data_bus[42]), .B2(n83), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U138 ( .A1(n66), .A2(n92), .B1(i_data_bus[43]), .B2(n83), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U139 ( .A1(n67), .A2(n84), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U140 ( .A1(n68), .A2(n84), .B1(i_data_bus[47]), .B2(n83), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U141 ( .A1(n69), .A2(n60), .B1(i_data_bus[49]), .B2(n83), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U142 ( .A1(n70), .A2(n60), .B1(i_data_bus[51]), .B2(n83), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U143 ( .A1(n71), .A2(n84), .B1(i_data_bus[52]), .B2(n83), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U144 ( .A1(n72), .A2(n84), .B1(i_data_bus[53]), .B2(n83), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U145 ( .A1(n73), .A2(n84), .B1(i_data_bus[54]), .B2(n83), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n74), .A2(n84), .B1(i_data_bus[55]), .B2(n83), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U147 ( .A1(n75), .A2(n84), .B1(i_data_bus[56]), .B2(n83), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U148 ( .A1(n76), .A2(n84), .B1(i_data_bus[58]), .B2(n83), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U149 ( .A1(n77), .A2(n84), .B1(i_data_bus[59]), .B2(n83), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U150 ( .A1(n78), .A2(n84), .B1(i_data_bus[60]), .B2(n83), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U151 ( .A1(n79), .A2(n60), .B1(i_data_bus[45]), .B2(n83), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U152 ( .A1(n80), .A2(n60), .B1(i_data_bus[46]), .B2(n83), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U153 ( .A1(n81), .A2(n84), .B1(i_data_bus[62]), .B2(n83), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U154 ( .A1(n82), .A2(n60), .B1(i_data_bus[48]), .B2(n83), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n84), .B1(i_data_bus[63]), .B2(n83), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_45 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  INVD1BWP30P140 U4 ( .I(n4), .ZN(n9) );
  NR2D1BWP30P140 U5 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  INVD1BWP30P140 U7 ( .I(n9), .ZN(n1) );
  INVD1BWP30P140 U8 ( .I(n9), .ZN(n2) );
  BUFFD12BWP30P140 U9 ( .I(n46), .Z(n48) );
  CKND2D3BWP30P140 U10 ( .A1(n7), .A2(n6), .ZN(n46) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U14 ( .I(n9), .ZN(n49) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n9), .ZN(n44) );
  INVD1BWP30P140 U18 ( .I(n78), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n44), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U24 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[36]), .ZN(n8) );
  OAI22D1BWP30P140 U26 ( .A1(n44), .A2(n59), .B1(n48), .B2(n8), .ZN(N291) );
  INVD1BWP30P140 U27 ( .I(n9), .ZN(n14) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[32]), .ZN(n10) );
  OAI22D1BWP30P140 U30 ( .A1(n2), .A2(n64), .B1(n48), .B2(n10), .ZN(N287) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[1]), .ZN(n62) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[33]), .ZN(n11) );
  OAI22D1BWP30P140 U33 ( .A1(n1), .A2(n62), .B1(n48), .B2(n11), .ZN(N288) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[2]), .ZN(n61) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[34]), .ZN(n12) );
  OAI22D1BWP30P140 U36 ( .A1(n49), .A2(n61), .B1(n48), .B2(n12), .ZN(N289) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[35]), .ZN(n13) );
  OAI22D1BWP30P140 U39 ( .A1(n14), .A2(n60), .B1(n48), .B2(n13), .ZN(N290) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[5]), .ZN(n58) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[37]), .ZN(n15) );
  OAI22D1BWP30P140 U42 ( .A1(n44), .A2(n58), .B1(n48), .B2(n15), .ZN(N292) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[6]), .ZN(n57) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[38]), .ZN(n16) );
  OAI22D1BWP30P140 U45 ( .A1(n44), .A2(n57), .B1(n48), .B2(n16), .ZN(N293) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[39]), .ZN(n17) );
  OAI22D1BWP30P140 U48 ( .A1(n44), .A2(n56), .B1(n46), .B2(n17), .ZN(N294) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[11]), .ZN(n87) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n44), .A2(n87), .B1(n48), .B2(n22), .ZN(N298) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[13]), .ZN(n85) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n1), .A2(n85), .B1(n48), .B2(n23), .ZN(N300) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[16]), .ZN(n82) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[48]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n49), .A2(n82), .B1(n48), .B2(n24), .ZN(N303) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[42]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n14), .A2(n88), .B1(n48), .B2(n25), .ZN(N297) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[44]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n2), .A2(n86), .B1(n48), .B2(n26), .ZN(N299) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[17]), .ZN(n81) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[49]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n1), .A2(n81), .B1(n48), .B2(n27), .ZN(N304) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[14]), .ZN(n84) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[46]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n49), .A2(n84), .B1(n48), .B2(n28), .ZN(N301) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[15]), .ZN(n83) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[47]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n14), .A2(n83), .B1(n48), .B2(n29), .ZN(N302) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[18]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[50]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n2), .A2(n80), .B1(n48), .B2(n30), .ZN(N305) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[19]), .ZN(n79) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[51]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n14), .A2(n79), .B1(n48), .B2(n31), .ZN(N306) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[52]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n2), .A2(n77), .B1(n48), .B2(n32), .ZN(N307) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[21]), .ZN(n75) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[53]), .ZN(n33) );
  OAI22D1BWP30P140 U87 ( .A1(n1), .A2(n75), .B1(n48), .B2(n33), .ZN(N308) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[23]), .ZN(n73) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[55]), .ZN(n34) );
  OAI22D1BWP30P140 U90 ( .A1(n49), .A2(n73), .B1(n48), .B2(n34), .ZN(N310) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[24]), .ZN(n72) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[56]), .ZN(n35) );
  OAI22D1BWP30P140 U93 ( .A1(n14), .A2(n72), .B1(n48), .B2(n35), .ZN(N311) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[25]), .ZN(n71) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[57]), .ZN(n36) );
  OAI22D1BWP30P140 U96 ( .A1(n2), .A2(n71), .B1(n48), .B2(n36), .ZN(N312) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[26]), .ZN(n70) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[58]), .ZN(n37) );
  OAI22D1BWP30P140 U99 ( .A1(n1), .A2(n70), .B1(n48), .B2(n37), .ZN(N313) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[59]), .ZN(n38) );
  OAI22D1BWP30P140 U102 ( .A1(n49), .A2(n69), .B1(n48), .B2(n38), .ZN(N314) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[28]), .ZN(n68) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[60]), .ZN(n39) );
  OAI22D1BWP30P140 U105 ( .A1(n14), .A2(n68), .B1(n48), .B2(n39), .ZN(N315) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[29]), .ZN(n67) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[61]), .ZN(n40) );
  OAI22D1BWP30P140 U108 ( .A1(n2), .A2(n67), .B1(n46), .B2(n40), .ZN(N316) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[30]), .ZN(n66) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[62]), .ZN(n41) );
  OAI22D1BWP30P140 U111 ( .A1(n1), .A2(n66), .B1(n48), .B2(n41), .ZN(N317) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[31]), .ZN(n65) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[63]), .ZN(n42) );
  OAI22D1BWP30P140 U114 ( .A1(n49), .A2(n65), .B1(n48), .B2(n42), .ZN(N318) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[54]), .ZN(n43) );
  OAI22D1BWP30P140 U117 ( .A1(n14), .A2(n74), .B1(n48), .B2(n43), .ZN(N309) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[8]), .ZN(n92) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[40]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n1), .A2(n92), .B1(n48), .B2(n45), .ZN(N295) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[9]), .ZN(n89) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[41]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n49), .A2(n89), .B1(n48), .B2(n47), .ZN(N296) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n78) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  INVD2BWP30P140 U135 ( .I(n78), .ZN(n76) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_46 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  INVD1BWP30P140 U4 ( .I(n4), .ZN(n13) );
  NR2D1BWP30P140 U5 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  INVD1BWP30P140 U7 ( .I(n13), .ZN(n1) );
  INVD1BWP30P140 U8 ( .I(n13), .ZN(n2) );
  BUFFD12BWP30P140 U9 ( .I(n46), .Z(n48) );
  CKND2D3BWP30P140 U10 ( .A1(n7), .A2(n6), .ZN(n46) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U14 ( .I(n13), .ZN(n33) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n13), .ZN(n49) );
  INVD1BWP30P140 U18 ( .I(n78), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n49), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n13), .ZN(n12) );
  INVD1BWP30P140 U24 ( .I(i_data_bus[0]), .ZN(n56) );
  INVD1BWP30P140 U25 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[32]), .ZN(n8) );
  OAI22D1BWP30P140 U27 ( .A1(n2), .A2(n56), .B1(n48), .B2(n8), .ZN(N287) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[1]), .ZN(n64) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[33]), .ZN(n9) );
  OAI22D1BWP30P140 U30 ( .A1(n1), .A2(n64), .B1(n48), .B2(n9), .ZN(N288) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[34]), .ZN(n10) );
  OAI22D1BWP30P140 U33 ( .A1(n33), .A2(n62), .B1(n48), .B2(n10), .ZN(N289) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[35]), .ZN(n11) );
  OAI22D1BWP30P140 U36 ( .A1(n12), .A2(n61), .B1(n48), .B2(n11), .ZN(N290) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[36]), .ZN(n14) );
  OAI22D1BWP30P140 U39 ( .A1(n49), .A2(n60), .B1(n48), .B2(n14), .ZN(N291) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[37]), .ZN(n15) );
  OAI22D1BWP30P140 U42 ( .A1(n49), .A2(n59), .B1(n48), .B2(n15), .ZN(N292) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[38]), .ZN(n16) );
  OAI22D1BWP30P140 U45 ( .A1(n49), .A2(n58), .B1(n48), .B2(n16), .ZN(N293) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[39]), .ZN(n17) );
  OAI22D1BWP30P140 U48 ( .A1(n49), .A2(n57), .B1(n46), .B2(n17), .ZN(N294) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[8]), .ZN(n92) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[40]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n49), .A2(n92), .B1(n48), .B2(n22), .ZN(N295) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[9]), .ZN(n89) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[41]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n1), .A2(n89), .B1(n48), .B2(n23), .ZN(N296) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[42]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n33), .A2(n88), .B1(n48), .B2(n24), .ZN(N297) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[11]), .ZN(n87) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[43]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n12), .A2(n87), .B1(n48), .B2(n25), .ZN(N298) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[44]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n2), .A2(n86), .B1(n48), .B2(n26), .ZN(N299) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[13]), .ZN(n85) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[45]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n1), .A2(n85), .B1(n48), .B2(n27), .ZN(N300) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[14]), .ZN(n84) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[46]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n33), .A2(n84), .B1(n48), .B2(n28), .ZN(N301) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[15]), .ZN(n83) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[47]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n12), .A2(n83), .B1(n48), .B2(n29), .ZN(N302) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[16]), .ZN(n82) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[48]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n2), .A2(n82), .B1(n46), .B2(n30), .ZN(N303) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[17]), .ZN(n81) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[49]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n1), .A2(n81), .B1(n48), .B2(n31), .ZN(N304) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[18]), .ZN(n80) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[50]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n33), .A2(n80), .B1(n48), .B2(n32), .ZN(N305) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[19]), .ZN(n79) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[51]), .ZN(n34) );
  OAI22D1BWP30P140 U87 ( .A1(n12), .A2(n79), .B1(n48), .B2(n34), .ZN(N306) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[52]), .ZN(n35) );
  OAI22D1BWP30P140 U90 ( .A1(n2), .A2(n77), .B1(n48), .B2(n35), .ZN(N307) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[21]), .ZN(n75) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[53]), .ZN(n36) );
  OAI22D1BWP30P140 U93 ( .A1(n1), .A2(n75), .B1(n48), .B2(n36), .ZN(N308) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[54]), .ZN(n37) );
  OAI22D1BWP30P140 U96 ( .A1(n33), .A2(n74), .B1(n48), .B2(n37), .ZN(N309) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[23]), .ZN(n73) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[55]), .ZN(n38) );
  OAI22D1BWP30P140 U99 ( .A1(n12), .A2(n73), .B1(n48), .B2(n38), .ZN(N310) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[24]), .ZN(n72) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[56]), .ZN(n39) );
  OAI22D1BWP30P140 U102 ( .A1(n2), .A2(n72), .B1(n48), .B2(n39), .ZN(N311) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[25]), .ZN(n71) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[57]), .ZN(n40) );
  OAI22D1BWP30P140 U105 ( .A1(n1), .A2(n71), .B1(n48), .B2(n40), .ZN(N312) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[26]), .ZN(n70) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[58]), .ZN(n41) );
  OAI22D1BWP30P140 U108 ( .A1(n33), .A2(n70), .B1(n48), .B2(n41), .ZN(N313) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[59]), .ZN(n42) );
  OAI22D1BWP30P140 U111 ( .A1(n12), .A2(n69), .B1(n48), .B2(n42), .ZN(N314) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[28]), .ZN(n68) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[60]), .ZN(n43) );
  OAI22D1BWP30P140 U114 ( .A1(n2), .A2(n68), .B1(n48), .B2(n43), .ZN(N315) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[29]), .ZN(n67) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[61]), .ZN(n44) );
  OAI22D1BWP30P140 U117 ( .A1(n1), .A2(n67), .B1(n48), .B2(n44), .ZN(N316) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[30]), .ZN(n66) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[62]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n33), .A2(n66), .B1(n48), .B2(n45), .ZN(N317) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[31]), .ZN(n65) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[63]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n12), .A2(n65), .B1(n48), .B2(n47), .ZN(N318) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n78) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n91), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  INVD2BWP30P140 U135 ( .I(n78), .ZN(n76) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_47 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  INVD1BWP30P140 U4 ( .I(n4), .ZN(n10) );
  NR2D1BWP30P140 U5 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  INVD1BWP30P140 U7 ( .I(n10), .ZN(n1) );
  INVD1BWP30P140 U8 ( .I(n10), .ZN(n2) );
  BUFFD12BWP30P140 U9 ( .I(n46), .Z(n48) );
  CKND2D3BWP30P140 U10 ( .A1(n7), .A2(n6), .ZN(n46) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U14 ( .I(n10), .ZN(n49) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n10), .ZN(n44) );
  INVD1BWP30P140 U18 ( .I(n78), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n44), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n10), .ZN(n17) );
  INVD1BWP30P140 U24 ( .I(i_data_bus[2]), .ZN(n61) );
  INVD1BWP30P140 U25 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[34]), .ZN(n8) );
  OAI22D1BWP30P140 U27 ( .A1(n1), .A2(n61), .B1(n48), .B2(n8), .ZN(N289) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[1]), .ZN(n62) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[33]), .ZN(n9) );
  OAI22D1BWP30P140 U30 ( .A1(n49), .A2(n62), .B1(n48), .B2(n9), .ZN(N288) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[36]), .ZN(n11) );
  OAI22D1BWP30P140 U33 ( .A1(n44), .A2(n59), .B1(n48), .B2(n11), .ZN(N291) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[5]), .ZN(n58) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[37]), .ZN(n12) );
  OAI22D1BWP30P140 U36 ( .A1(n44), .A2(n58), .B1(n48), .B2(n12), .ZN(N292) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[6]), .ZN(n57) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[38]), .ZN(n13) );
  OAI22D1BWP30P140 U39 ( .A1(n44), .A2(n57), .B1(n48), .B2(n13), .ZN(N293) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[39]), .ZN(n14) );
  OAI22D1BWP30P140 U42 ( .A1(n44), .A2(n56), .B1(n48), .B2(n14), .ZN(N294) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[35]), .ZN(n15) );
  OAI22D1BWP30P140 U45 ( .A1(n17), .A2(n60), .B1(n48), .B2(n15), .ZN(N290) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[32]), .ZN(n16) );
  OAI22D1BWP30P140 U48 ( .A1(n2), .A2(n64), .B1(n46), .B2(n16), .ZN(N287) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[42]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n44), .A2(n88), .B1(n48), .B2(n22), .ZN(N297) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[11]), .ZN(n87) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[43]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n1), .A2(n87), .B1(n48), .B2(n23), .ZN(N298) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[44]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n49), .A2(n86), .B1(n48), .B2(n24), .ZN(N299) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[13]), .ZN(n85) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[45]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n17), .A2(n85), .B1(n48), .B2(n25), .ZN(N300) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[14]), .ZN(n84) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[46]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n2), .A2(n84), .B1(n48), .B2(n26), .ZN(N301) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[15]), .ZN(n83) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[47]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n1), .A2(n83), .B1(n48), .B2(n27), .ZN(N302) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[16]), .ZN(n82) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[48]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n49), .A2(n82), .B1(n48), .B2(n28), .ZN(N303) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[17]), .ZN(n81) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[49]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n17), .A2(n81), .B1(n48), .B2(n29), .ZN(N304) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[18]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[50]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n2), .A2(n80), .B1(n48), .B2(n30), .ZN(N305) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[19]), .ZN(n79) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[51]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n17), .A2(n79), .B1(n48), .B2(n31), .ZN(N306) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[52]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n2), .A2(n77), .B1(n48), .B2(n32), .ZN(N307) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[21]), .ZN(n75) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[53]), .ZN(n33) );
  OAI22D1BWP30P140 U87 ( .A1(n1), .A2(n75), .B1(n48), .B2(n33), .ZN(N308) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[54]), .ZN(n34) );
  OAI22D1BWP30P140 U90 ( .A1(n49), .A2(n74), .B1(n48), .B2(n34), .ZN(N309) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[23]), .ZN(n73) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[55]), .ZN(n35) );
  OAI22D1BWP30P140 U93 ( .A1(n17), .A2(n73), .B1(n48), .B2(n35), .ZN(N310) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[24]), .ZN(n72) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[56]), .ZN(n36) );
  OAI22D1BWP30P140 U96 ( .A1(n2), .A2(n72), .B1(n48), .B2(n36), .ZN(N311) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[25]), .ZN(n71) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[57]), .ZN(n37) );
  OAI22D1BWP30P140 U99 ( .A1(n1), .A2(n71), .B1(n48), .B2(n37), .ZN(N312) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[26]), .ZN(n70) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[58]), .ZN(n38) );
  OAI22D1BWP30P140 U102 ( .A1(n49), .A2(n70), .B1(n48), .B2(n38), .ZN(N313) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[59]), .ZN(n39) );
  OAI22D1BWP30P140 U105 ( .A1(n17), .A2(n69), .B1(n48), .B2(n39), .ZN(N314) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[28]), .ZN(n68) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[60]), .ZN(n40) );
  OAI22D1BWP30P140 U108 ( .A1(n2), .A2(n68), .B1(n46), .B2(n40), .ZN(N315) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[29]), .ZN(n67) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[61]), .ZN(n41) );
  OAI22D1BWP30P140 U111 ( .A1(n1), .A2(n67), .B1(n48), .B2(n41), .ZN(N316) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[30]), .ZN(n66) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[62]), .ZN(n42) );
  OAI22D1BWP30P140 U114 ( .A1(n49), .A2(n66), .B1(n48), .B2(n42), .ZN(N317) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[31]), .ZN(n65) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[63]), .ZN(n43) );
  OAI22D1BWP30P140 U117 ( .A1(n17), .A2(n65), .B1(n48), .B2(n43), .ZN(N318) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[9]), .ZN(n89) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[41]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n1), .A2(n89), .B1(n48), .B2(n45), .ZN(N296) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[8]), .ZN(n92) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[40]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n49), .A2(n92), .B1(n48), .B2(n47), .ZN(N295) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n78) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  INVD2BWP30P140 U135 ( .I(n78), .ZN(n76) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_48 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  AN3D4BWP30P140 U3 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n19), .Z(n90) );
  INVD1BWP30P140 U4 ( .I(n4), .ZN(n10) );
  NR2D1BWP30P140 U5 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  INR2D1BWP30P140 U6 ( .A1(i_valid[0]), .B1(n50), .ZN(n18) );
  INVD1BWP30P140 U7 ( .I(n10), .ZN(n1) );
  INVD1BWP30P140 U8 ( .I(n10), .ZN(n2) );
  BUFFD12BWP30P140 U9 ( .I(n46), .Z(n48) );
  CKND2D3BWP30P140 U10 ( .A1(n7), .A2(n6), .ZN(n46) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n18), .A2(n5), .ZN(n4) );
  ND2D1BWP30P140 U12 ( .A1(n3), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U14 ( .I(n10), .ZN(n49) );
  MUX2NUD1BWP30P140 U15 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n7) );
  NR2D1BWP30P140 U16 ( .A1(n50), .A2(n5), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n10), .ZN(n35) );
  INVD1BWP30P140 U18 ( .I(n78), .ZN(n63) );
  INVD1BWP30P140 U19 ( .I(n90), .ZN(n20) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(i_valid[1]), .ZN(n51) );
  OAI31D1BWP30P140 U22 ( .A1(n50), .A2(n51), .A3(n5), .B(n35), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n10), .ZN(n15) );
  INVD1BWP30P140 U24 ( .I(i_data_bus[2]), .ZN(n58) );
  INVD1BWP30P140 U25 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[34]), .ZN(n8) );
  OAI22D1BWP30P140 U27 ( .A1(n2), .A2(n58), .B1(n48), .B2(n8), .ZN(N289) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[0]), .ZN(n56) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[32]), .ZN(n9) );
  OAI22D1BWP30P140 U30 ( .A1(n1), .A2(n56), .B1(n48), .B2(n9), .ZN(N287) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[5]), .ZN(n61) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[37]), .ZN(n11) );
  OAI22D1BWP30P140 U33 ( .A1(n35), .A2(n61), .B1(n48), .B2(n11), .ZN(N292) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[36]), .ZN(n12) );
  OAI22D1BWP30P140 U36 ( .A1(n35), .A2(n60), .B1(n48), .B2(n12), .ZN(N291) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[3]), .ZN(n59) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[35]), .ZN(n13) );
  OAI22D1BWP30P140 U39 ( .A1(n49), .A2(n59), .B1(n48), .B2(n13), .ZN(N290) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[1]), .ZN(n57) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[33]), .ZN(n14) );
  OAI22D1BWP30P140 U42 ( .A1(n15), .A2(n57), .B1(n48), .B2(n14), .ZN(N288) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[6]), .ZN(n62) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[38]), .ZN(n16) );
  OAI22D1BWP30P140 U45 ( .A1(n35), .A2(n62), .B1(n48), .B2(n16), .ZN(N293) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[39]), .ZN(n17) );
  OAI22D1BWP30P140 U48 ( .A1(n35), .A2(n64), .B1(n46), .B2(n17), .ZN(N294) );
  INVD1BWP30P140 U49 ( .I(n18), .ZN(n21) );
  INVD1BWP30P140 U50 ( .I(n50), .ZN(n19) );
  OAI21D1BWP30P140 U51 ( .A1(n21), .A2(i_cmd[1]), .B(n20), .ZN(N354) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[63]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n15), .A2(n92), .B1(n48), .B2(n22), .ZN(N318) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[62]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n2), .A2(n89), .B1(n48), .B2(n23), .ZN(N317) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[61]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n1), .A2(n88), .B1(n48), .B2(n24), .ZN(N316) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[60]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n49), .A2(n87), .B1(n48), .B2(n25), .ZN(N315) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[59]), .ZN(n26) );
  OAI22D1BWP30P140 U66 ( .A1(n15), .A2(n86), .B1(n48), .B2(n26), .ZN(N314) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[58]), .ZN(n27) );
  OAI22D1BWP30P140 U69 ( .A1(n2), .A2(n85), .B1(n48), .B2(n27), .ZN(N313) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[57]), .ZN(n28) );
  OAI22D1BWP30P140 U72 ( .A1(n1), .A2(n84), .B1(n48), .B2(n28), .ZN(N312) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[56]), .ZN(n29) );
  OAI22D1BWP30P140 U75 ( .A1(n49), .A2(n83), .B1(n48), .B2(n29), .ZN(N311) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[55]), .ZN(n30) );
  OAI22D1BWP30P140 U78 ( .A1(n15), .A2(n82), .B1(n46), .B2(n30), .ZN(N310) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[54]), .ZN(n31) );
  OAI22D1BWP30P140 U81 ( .A1(n2), .A2(n81), .B1(n48), .B2(n31), .ZN(N309) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[53]), .ZN(n32) );
  OAI22D1BWP30P140 U84 ( .A1(n1), .A2(n80), .B1(n48), .B2(n32), .ZN(N308) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[52]), .ZN(n33) );
  OAI22D1BWP30P140 U87 ( .A1(n49), .A2(n79), .B1(n48), .B2(n33), .ZN(N307) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[19]), .ZN(n77) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[51]), .ZN(n34) );
  OAI22D1BWP30P140 U90 ( .A1(n15), .A2(n77), .B1(n48), .B2(n34), .ZN(N306) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[50]), .ZN(n36) );
  OAI22D1BWP30P140 U93 ( .A1(n35), .A2(n75), .B1(n48), .B2(n36), .ZN(N305) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[49]), .ZN(n37) );
  OAI22D1BWP30P140 U96 ( .A1(n1), .A2(n74), .B1(n48), .B2(n37), .ZN(N304) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[48]), .ZN(n38) );
  OAI22D1BWP30P140 U99 ( .A1(n49), .A2(n73), .B1(n48), .B2(n38), .ZN(N303) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[47]), .ZN(n39) );
  OAI22D1BWP30P140 U102 ( .A1(n15), .A2(n72), .B1(n48), .B2(n39), .ZN(N302) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[46]), .ZN(n40) );
  OAI22D1BWP30P140 U105 ( .A1(n2), .A2(n71), .B1(n48), .B2(n40), .ZN(N301) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[45]), .ZN(n41) );
  OAI22D1BWP30P140 U108 ( .A1(n1), .A2(n70), .B1(n48), .B2(n41), .ZN(N300) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[44]), .ZN(n42) );
  OAI22D1BWP30P140 U111 ( .A1(n49), .A2(n69), .B1(n48), .B2(n42), .ZN(N299) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[43]), .ZN(n43) );
  OAI22D1BWP30P140 U114 ( .A1(n15), .A2(n68), .B1(n48), .B2(n43), .ZN(N298) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[42]), .ZN(n44) );
  OAI22D1BWP30P140 U117 ( .A1(n2), .A2(n67), .B1(n48), .B2(n44), .ZN(N297) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[41]), .ZN(n45) );
  OAI22D1BWP30P140 U120 ( .A1(n1), .A2(n66), .B1(n48), .B2(n45), .ZN(N296) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[40]), .ZN(n47) );
  OAI22D1BWP30P140 U123 ( .A1(n49), .A2(n65), .B1(n48), .B2(n47), .ZN(N295) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n78) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n91), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  INVD2BWP30P140 U135 ( .I(n78), .ZN(n76) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_49 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  ND2OPTPAD6BWP30P140 U3 ( .A1(n35), .A2(n34), .ZN(n69) );
  INVD6BWP30P140 U4 ( .I(n36), .ZN(n68) );
  INVD3BWP30P140 U5 ( .I(n32), .ZN(n35) );
  NR2D2BWP30P140 U6 ( .A1(i_cmd[1]), .A2(n33), .ZN(n34) );
  CKND2D4BWP30P140 U7 ( .A1(n25), .A2(n1), .ZN(n71) );
  ND2OPTPAD4BWP30P140 U8 ( .A1(n30), .A2(n7), .ZN(n14) );
  INVD3BWP30P140 U9 ( .I(n3), .ZN(n30) );
  CKND2D3BWP30P140 U10 ( .A1(i_valid[0]), .A2(n11), .ZN(n3) );
  INVD4BWP30P140 U11 ( .I(i_valid[1]), .ZN(n9) );
  ND2D1BWP30P140 U12 ( .A1(n29), .A2(n28), .ZN(N295) );
  BUFFD1BWP30P140 U13 ( .I(i_valid[1]), .Z(n4) );
  ND2D1BWP30P140 U14 ( .A1(n2), .A2(i_en), .ZN(n33) );
  INVD6BWP30P140 U15 ( .I(n14), .ZN(n93) );
  ND2OPTIBD1BWP30P140 U16 ( .A1(n14), .A2(n8), .ZN(N353) );
  IND2D1BWP30P140 U17 ( .A1(n7), .B1(n6), .ZN(n8) );
  NR2D1BWP30P140 U18 ( .A1(n5), .A2(n33), .ZN(n6) );
  INVD1BWP30P140 U19 ( .I(n4), .ZN(n5) );
  OAI22D1BWP30P140 U20 ( .A1(n22), .A2(n12), .B1(n14), .B2(n52), .ZN(N304) );
  OAI22D1BWP30P140 U21 ( .A1(n22), .A2(n13), .B1(n14), .B2(n40), .ZN(N316) );
  AN2D4BWP30P140 U22 ( .A1(i_cmd[0]), .A2(n11), .Z(n1) );
  INVD1BWP30P140 U23 ( .I(n33), .ZN(n11) );
  INVD1BWP30P140 U24 ( .I(rst), .ZN(n2) );
  INVD2BWP30P140 U25 ( .I(i_cmd[0]), .ZN(n7) );
  INVD2BWP30P140 U26 ( .I(i_valid[0]), .ZN(n10) );
  MUX2NOPTD4BWP30P140 U27 ( .I0(n10), .I1(n9), .S(i_cmd[1]), .ZN(n25) );
  BUFFD4BWP30P140 U28 ( .I(n71), .Z(n22) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[49]), .ZN(n12) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[17]), .ZN(n52) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[61]), .ZN(n13) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[29]), .ZN(n40) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[62]), .ZN(n15) );
  MOAI22D1BWP30P140 U34 ( .A1(n22), .A2(n15), .B1(n93), .B2(i_data_bus[30]), 
        .ZN(N317) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[63]), .ZN(n16) );
  MOAI22D1BWP30P140 U36 ( .A1(n22), .A2(n16), .B1(n93), .B2(i_data_bus[31]), 
        .ZN(N318) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[35]), .ZN(n17) );
  MOAI22D1BWP30P140 U38 ( .A1(n22), .A2(n17), .B1(n93), .B2(i_data_bus[3]), 
        .ZN(N290) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[36]), .ZN(n18) );
  MOAI22D1BWP30P140 U40 ( .A1(n22), .A2(n18), .B1(n93), .B2(i_data_bus[4]), 
        .ZN(N291) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[37]), .ZN(n19) );
  MOAI22D1BWP30P140 U42 ( .A1(n22), .A2(n19), .B1(n93), .B2(i_data_bus[5]), 
        .ZN(N292) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[38]), .ZN(n20) );
  MOAI22D1BWP30P140 U44 ( .A1(n22), .A2(n20), .B1(n93), .B2(i_data_bus[6]), 
        .ZN(N293) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[39]), .ZN(n21) );
  MOAI22D1BWP30P140 U46 ( .A1(n22), .A2(n21), .B1(n93), .B2(i_data_bus[7]), 
        .ZN(N294) );
  BUFFD4BWP30P140 U47 ( .I(n71), .Z(n92) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[50]), .ZN(n23) );
  MOAI22D1BWP30P140 U49 ( .A1(n92), .A2(n23), .B1(n93), .B2(i_data_bus[18]), 
        .ZN(N305) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[51]), .ZN(n24) );
  MOAI22D1BWP30P140 U51 ( .A1(n92), .A2(n24), .B1(n93), .B2(i_data_bus[19]), 
        .ZN(N306) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[40]), .ZN(n27) );
  CKBD1BWP30P140 U53 ( .I(n25), .Z(n26) );
  IND3D1BWP30P140 U54 ( .A1(n27), .B1(n1), .B2(n26), .ZN(n29) );
  ND2D1BWP30P140 U55 ( .A1(n93), .A2(i_data_bus[8]), .ZN(n28) );
  INVD1BWP30P140 U56 ( .I(n30), .ZN(n31) );
  ND3OPTPAD4BWP30P140 U57 ( .A1(i_cmd[1]), .A2(i_valid[1]), .A3(n11), .ZN(n36)
         );
  OAI21D1BWP30P140 U58 ( .A1(n31), .A2(i_cmd[1]), .B(n36), .ZN(N354) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[0]), .ZN(n37) );
  MUX2NOPTD2BWP30P140 U60 ( .I0(i_valid[0]), .I1(i_valid[1]), .S(i_cmd[0]), 
        .ZN(n32) );
  MOAI22D1BWP30P140 U61 ( .A1(n37), .A2(n69), .B1(i_data_bus[32]), .B2(n68), 
        .ZN(N319) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[31]), .ZN(n38) );
  MOAI22D1BWP30P140 U63 ( .A1(n38), .A2(n69), .B1(i_data_bus[63]), .B2(n68), 
        .ZN(N350) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[30]), .ZN(n39) );
  MOAI22D1BWP30P140 U65 ( .A1(n39), .A2(n69), .B1(i_data_bus[62]), .B2(n68), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U66 ( .A1(n40), .A2(n69), .B1(i_data_bus[61]), .B2(n68), 
        .ZN(N348) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[28]), .ZN(n41) );
  MOAI22D1BWP30P140 U68 ( .A1(n41), .A2(n69), .B1(i_data_bus[60]), .B2(n68), 
        .ZN(N347) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[27]), .ZN(n42) );
  MOAI22D1BWP30P140 U70 ( .A1(n42), .A2(n69), .B1(i_data_bus[59]), .B2(n68), 
        .ZN(N346) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[26]), .ZN(n43) );
  MOAI22D1BWP30P140 U72 ( .A1(n43), .A2(n69), .B1(i_data_bus[58]), .B2(n68), 
        .ZN(N345) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[25]), .ZN(n44) );
  MOAI22D1BWP30P140 U74 ( .A1(n44), .A2(n69), .B1(i_data_bus[57]), .B2(n68), 
        .ZN(N344) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[24]), .ZN(n45) );
  MOAI22D1BWP30P140 U76 ( .A1(n45), .A2(n69), .B1(i_data_bus[56]), .B2(n68), 
        .ZN(N343) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[23]), .ZN(n46) );
  MOAI22D1BWP30P140 U78 ( .A1(n46), .A2(n69), .B1(i_data_bus[55]), .B2(n68), 
        .ZN(N342) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[22]), .ZN(n47) );
  MOAI22D1BWP30P140 U80 ( .A1(n47), .A2(n69), .B1(i_data_bus[54]), .B2(n68), 
        .ZN(N341) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[21]), .ZN(n48) );
  MOAI22D1BWP30P140 U82 ( .A1(n48), .A2(n69), .B1(i_data_bus[53]), .B2(n68), 
        .ZN(N340) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[20]), .ZN(n49) );
  MOAI22D1BWP30P140 U84 ( .A1(n49), .A2(n69), .B1(i_data_bus[52]), .B2(n68), 
        .ZN(N339) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[19]), .ZN(n50) );
  MOAI22D1BWP30P140 U86 ( .A1(n50), .A2(n69), .B1(i_data_bus[51]), .B2(n68), 
        .ZN(N338) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[18]), .ZN(n51) );
  MOAI22D1BWP30P140 U88 ( .A1(n51), .A2(n69), .B1(i_data_bus[50]), .B2(n68), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U89 ( .A1(n52), .A2(n69), .B1(i_data_bus[49]), .B2(n68), 
        .ZN(N336) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[16]), .ZN(n53) );
  MOAI22D1BWP30P140 U91 ( .A1(n53), .A2(n69), .B1(i_data_bus[48]), .B2(n68), 
        .ZN(N335) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[15]), .ZN(n54) );
  MOAI22D1BWP30P140 U93 ( .A1(n54), .A2(n69), .B1(i_data_bus[47]), .B2(n68), 
        .ZN(N334) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[14]), .ZN(n55) );
  MOAI22D1BWP30P140 U95 ( .A1(n55), .A2(n69), .B1(i_data_bus[46]), .B2(n68), 
        .ZN(N333) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[13]), .ZN(n56) );
  MOAI22D1BWP30P140 U97 ( .A1(n56), .A2(n69), .B1(i_data_bus[45]), .B2(n68), 
        .ZN(N332) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[12]), .ZN(n57) );
  MOAI22D1BWP30P140 U99 ( .A1(n57), .A2(n69), .B1(i_data_bus[44]), .B2(n68), 
        .ZN(N331) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[11]), .ZN(n58) );
  MOAI22D1BWP30P140 U101 ( .A1(n58), .A2(n69), .B1(i_data_bus[43]), .B2(n68), 
        .ZN(N330) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[10]), .ZN(n59) );
  MOAI22D1BWP30P140 U103 ( .A1(n59), .A2(n69), .B1(i_data_bus[42]), .B2(n68), 
        .ZN(N329) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[9]), .ZN(n60) );
  MOAI22D1BWP30P140 U105 ( .A1(n60), .A2(n69), .B1(i_data_bus[41]), .B2(n68), 
        .ZN(N328) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[8]), .ZN(n61) );
  MOAI22D1BWP30P140 U107 ( .A1(n61), .A2(n69), .B1(i_data_bus[40]), .B2(n68), 
        .ZN(N327) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[7]), .ZN(n62) );
  MOAI22D1BWP30P140 U109 ( .A1(n62), .A2(n69), .B1(i_data_bus[39]), .B2(n68), 
        .ZN(N326) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[6]), .ZN(n63) );
  MOAI22D1BWP30P140 U111 ( .A1(n63), .A2(n69), .B1(i_data_bus[38]), .B2(n68), 
        .ZN(N325) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[5]), .ZN(n64) );
  MOAI22D1BWP30P140 U113 ( .A1(n64), .A2(n69), .B1(i_data_bus[37]), .B2(n68), 
        .ZN(N324) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[4]), .ZN(n65) );
  MOAI22D1BWP30P140 U115 ( .A1(n65), .A2(n69), .B1(i_data_bus[36]), .B2(n68), 
        .ZN(N323) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[3]), .ZN(n66) );
  MOAI22D1BWP30P140 U117 ( .A1(n66), .A2(n69), .B1(i_data_bus[35]), .B2(n68), 
        .ZN(N322) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[2]), .ZN(n67) );
  MOAI22D1BWP30P140 U119 ( .A1(n67), .A2(n69), .B1(i_data_bus[34]), .B2(n68), 
        .ZN(N321) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[1]), .ZN(n70) );
  MOAI22D1BWP30P140 U121 ( .A1(n70), .A2(n69), .B1(i_data_bus[33]), .B2(n68), 
        .ZN(N320) );
  INVD2BWP30P140 U122 ( .I(n71), .ZN(n72) );
  INVD4BWP30P140 U123 ( .I(n72), .ZN(n95) );
  INVD1BWP30P140 U124 ( .I(i_data_bus[60]), .ZN(n73) );
  MOAI22D1BWP30P140 U125 ( .A1(n95), .A2(n73), .B1(n93), .B2(i_data_bus[28]), 
        .ZN(N315) );
  INVD1BWP30P140 U126 ( .I(i_data_bus[48]), .ZN(n74) );
  MOAI22D1BWP30P140 U127 ( .A1(n92), .A2(n74), .B1(n93), .B2(i_data_bus[16]), 
        .ZN(N303) );
  INVD1BWP30P140 U128 ( .I(i_data_bus[34]), .ZN(n75) );
  MOAI22D1BWP30P140 U129 ( .A1(n95), .A2(n75), .B1(n93), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140 U130 ( .I(i_data_bus[59]), .ZN(n76) );
  MOAI22D1BWP30P140 U131 ( .A1(n95), .A2(n76), .B1(n93), .B2(i_data_bus[27]), 
        .ZN(N314) );
  INVD1BWP30P140 U132 ( .I(i_data_bus[47]), .ZN(n77) );
  MOAI22D1BWP30P140 U133 ( .A1(n92), .A2(n77), .B1(n93), .B2(i_data_bus[15]), 
        .ZN(N302) );
  INVD1BWP30P140 U134 ( .I(i_data_bus[33]), .ZN(n78) );
  MOAI22D1BWP30P140 U135 ( .A1(n95), .A2(n78), .B1(n93), .B2(i_data_bus[1]), 
        .ZN(N288) );
  INVD1BWP30P140 U136 ( .I(i_data_bus[58]), .ZN(n79) );
  MOAI22D1BWP30P140 U137 ( .A1(n95), .A2(n79), .B1(n93), .B2(i_data_bus[26]), 
        .ZN(N313) );
  INVD1BWP30P140 U138 ( .I(i_data_bus[46]), .ZN(n80) );
  MOAI22D1BWP30P140 U139 ( .A1(n92), .A2(n80), .B1(n93), .B2(i_data_bus[14]), 
        .ZN(N301) );
  INVD1BWP30P140 U140 ( .I(i_data_bus[32]), .ZN(n81) );
  MOAI22D1BWP30P140 U141 ( .A1(n95), .A2(n81), .B1(n93), .B2(i_data_bus[0]), 
        .ZN(N287) );
  INVD1BWP30P140 U142 ( .I(i_data_bus[57]), .ZN(n82) );
  MOAI22D1BWP30P140 U143 ( .A1(n95), .A2(n82), .B1(n93), .B2(i_data_bus[25]), 
        .ZN(N312) );
  INVD1BWP30P140 U144 ( .I(i_data_bus[45]), .ZN(n83) );
  MOAI22D1BWP30P140 U145 ( .A1(n92), .A2(n83), .B1(n93), .B2(i_data_bus[13]), 
        .ZN(N300) );
  INVD1BWP30P140 U146 ( .I(i_data_bus[56]), .ZN(n84) );
  MOAI22D1BWP30P140 U147 ( .A1(n95), .A2(n84), .B1(n93), .B2(i_data_bus[24]), 
        .ZN(N311) );
  INVD1BWP30P140 U148 ( .I(i_data_bus[44]), .ZN(n85) );
  MOAI22D1BWP30P140 U149 ( .A1(n92), .A2(n85), .B1(n93), .B2(i_data_bus[12]), 
        .ZN(N299) );
  INVD1BWP30P140 U150 ( .I(i_data_bus[55]), .ZN(n86) );
  MOAI22D1BWP30P140 U151 ( .A1(n95), .A2(n86), .B1(n93), .B2(i_data_bus[23]), 
        .ZN(N310) );
  INVD1BWP30P140 U152 ( .I(i_data_bus[43]), .ZN(n87) );
  MOAI22D1BWP30P140 U153 ( .A1(n92), .A2(n87), .B1(n93), .B2(i_data_bus[11]), 
        .ZN(N298) );
  INVD1BWP30P140 U154 ( .I(i_data_bus[54]), .ZN(n88) );
  MOAI22D1BWP30P140 U155 ( .A1(n95), .A2(n88), .B1(n93), .B2(i_data_bus[22]), 
        .ZN(N309) );
  INVD1BWP30P140 U156 ( .I(i_data_bus[42]), .ZN(n89) );
  MOAI22D1BWP30P140 U157 ( .A1(n92), .A2(n89), .B1(n93), .B2(i_data_bus[10]), 
        .ZN(N297) );
  INVD1BWP30P140 U158 ( .I(i_data_bus[53]), .ZN(n90) );
  MOAI22D1BWP30P140 U159 ( .A1(n95), .A2(n90), .B1(n93), .B2(i_data_bus[21]), 
        .ZN(N308) );
  INVD1BWP30P140 U160 ( .I(i_data_bus[41]), .ZN(n91) );
  MOAI22D1BWP30P140 U161 ( .A1(n92), .A2(n91), .B1(n93), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140 U162 ( .I(i_data_bus[52]), .ZN(n94) );
  MOAI22D1BWP30P140 U163 ( .A1(n95), .A2(n94), .B1(n93), .B2(i_data_bus[20]), 
        .ZN(N307) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_50 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  INVD3BWP30P140 U3 ( .I(n82), .ZN(n126) );
  INVD6BWP30P140 U4 ( .I(n106), .ZN(n127) );
  INVD3BWP30P140 U5 ( .I(n35), .ZN(n82) );
  INVD1BWP30P140 U6 ( .I(n13), .ZN(n14) );
  INR2D6BWP30P140 U7 ( .A1(i_valid[1]), .B1(n16), .ZN(n93) );
  CKND2D4BWP30P140 U8 ( .A1(n92), .A2(n90), .ZN(n106) );
  CKND2D3BWP30P140 U9 ( .A1(n10), .A2(n9), .ZN(n35) );
  CKND2D3BWP30P140 U10 ( .A1(i_cmd[1]), .A2(n6), .ZN(n16) );
  NR2D1BWP30P140 U11 ( .A1(i_cmd[1]), .A2(n87), .ZN(n13) );
  NR2OPTPAD2BWP30P140 U12 ( .A1(n8), .A2(n7), .ZN(n10) );
  INVD2BWP30P140 U13 ( .I(n11), .ZN(n92) );
  ND2OPTIBD2BWP30P140 U14 ( .A1(n88), .A2(i_cmd[1]), .ZN(n9) );
  NR2D1P5BWP30P140 U15 ( .A1(i_cmd[1]), .A2(i_valid[0]), .ZN(n8) );
  OAI22D2BWP30P140 U16 ( .A1(n1), .A2(n97), .B1(n118), .B2(n96), .ZN(N294) );
  INVD4BWP30P140 U17 ( .I(n82), .ZN(n118) );
  ND2D1BWP30P140 U18 ( .A1(n2), .A2(n91), .ZN(N353) );
  INVD1BWP30P140 U19 ( .I(n127), .ZN(n1) );
  CKND2D3BWP30P140 U20 ( .A1(i_valid[0]), .A2(n6), .ZN(n11) );
  ND2OPTIBD1BWP30P140 U21 ( .A1(n92), .A2(n90), .ZN(n2) );
  INVD1BWP30P140 U22 ( .I(i_cmd[0]), .ZN(n90) );
  BUFFD4BWP30P140 U23 ( .I(n35), .Z(n129) );
  CKND2D3BWP30P140 U24 ( .A1(i_cmd[0]), .A2(n6), .ZN(n7) );
  ND2D1BWP30P140 U25 ( .A1(n5), .A2(i_en), .ZN(n87) );
  INVD1BWP30P140 U26 ( .I(n93), .ZN(n94) );
  IND2D1BWP30P140 U27 ( .A1(n90), .B1(n89), .ZN(n91) );
  NR2D1BWP30P140 U28 ( .A1(n88), .A2(n87), .ZN(n89) );
  INVD1BWP30P140 U29 ( .I(i_valid[1]), .ZN(n88) );
  OAI21D1BWP30P140 U30 ( .A1(n118), .A2(n84), .B(n83), .ZN(N288) );
  ND2OPTIBD1BWP30P140 U31 ( .A1(n127), .A2(i_data_bus[1]), .ZN(n83) );
  OAI22D1BWP30P140 U32 ( .A1(n35), .A2(n34), .B1(n2), .B2(n53), .ZN(N304) );
  OAI22D1BWP30P140 U33 ( .A1(n129), .A2(n31), .B1(n2), .B2(n55), .ZN(N305) );
  OAI22D1BWP30P140 U34 ( .A1(n129), .A2(n30), .B1(n2), .B2(n57), .ZN(N306) );
  ND2D1BWP30P140 U35 ( .A1(n93), .A2(i_data_bus[53]), .ZN(n60) );
  ND2D1BWP30P140 U36 ( .A1(n93), .A2(i_data_bus[54]), .ZN(n62) );
  ND2D1BWP30P140 U37 ( .A1(n93), .A2(i_data_bus[55]), .ZN(n64) );
  ND2D1BWP30P140 U38 ( .A1(n93), .A2(i_data_bus[56]), .ZN(n66) );
  ND2D1BWP30P140 U39 ( .A1(n93), .A2(i_data_bus[57]), .ZN(n68) );
  ND2D1BWP30P140 U40 ( .A1(n93), .A2(i_data_bus[58]), .ZN(n70) );
  ND2D1BWP30P140 U41 ( .A1(n93), .A2(i_data_bus[59]), .ZN(n72) );
  ND2D1BWP30P140 U42 ( .A1(n93), .A2(i_data_bus[60]), .ZN(n74) );
  ND2D1BWP30P140 U43 ( .A1(n93), .A2(i_data_bus[61]), .ZN(n76) );
  ND2D1BWP30P140 U44 ( .A1(n93), .A2(i_data_bus[62]), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U45 ( .A1(n93), .A2(i_data_bus[63]), .ZN(n80) );
  MOAI22D1BWP30P140 U46 ( .A1(n118), .A2(n104), .B1(n127), .B2(i_data_bus[6]), 
        .ZN(N293) );
  MOAI22D1BWP30P140 U47 ( .A1(n118), .A2(n98), .B1(n127), .B2(i_data_bus[5]), 
        .ZN(N292) );
  MOAI22D1BWP30P140 U48 ( .A1(n126), .A2(n32), .B1(n127), .B2(i_data_bus[31]), 
        .ZN(N318) );
  MOAI22D1BWP30P140 U49 ( .A1(n118), .A2(n100), .B1(n127), .B2(i_data_bus[4]), 
        .ZN(N291) );
  MOAI22D1BWP30P140 U50 ( .A1(n118), .A2(n102), .B1(n127), .B2(i_data_bus[3]), 
        .ZN(N290) );
  MOAI22D1BWP30P140 U51 ( .A1(n126), .A2(n33), .B1(n127), .B2(i_data_bus[29]), 
        .ZN(N316) );
  OR2D4BWP30P140 U52 ( .A1(n15), .A2(n14), .Z(n3) );
  MOAI22D1BWP30P140 U53 ( .A1(n126), .A2(n12), .B1(n127), .B2(i_data_bus[30]), 
        .ZN(N317) );
  OR2D4BWP30P140 U54 ( .A1(n15), .A2(n14), .Z(n4) );
  INVD1BWP30P140 U55 ( .I(n87), .ZN(n6) );
  INVD1BWP30P140 U56 ( .I(rst), .ZN(n5) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[62]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[30]), .ZN(n79) );
  MUX2NOPTD2BWP30P140 U59 ( .I0(i_valid[0]), .I1(i_valid[1]), .S(i_cmd[0]), 
        .ZN(n15) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[0]), .ZN(n18) );
  ND2OPTIBD1BWP30P140 U61 ( .A1(n93), .A2(i_data_bus[32]), .ZN(n17) );
  OAI21D1BWP30P140 U62 ( .A1(n4), .A2(n18), .B(n17), .ZN(N319) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[1]), .ZN(n20) );
  ND2OPTIBD1BWP30P140 U64 ( .A1(n93), .A2(i_data_bus[33]), .ZN(n19) );
  OAI21D1BWP30P140 U65 ( .A1(n4), .A2(n20), .B(n19), .ZN(N320) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[2]), .ZN(n22) );
  ND2OPTIBD1BWP30P140 U67 ( .A1(n93), .A2(i_data_bus[34]), .ZN(n21) );
  OAI21D1BWP30P140 U68 ( .A1(n4), .A2(n22), .B(n21), .ZN(N321) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[3]), .ZN(n103) );
  ND2OPTIBD1BWP30P140 U70 ( .A1(n93), .A2(i_data_bus[35]), .ZN(n23) );
  OAI21D1BWP30P140 U71 ( .A1(n4), .A2(n103), .B(n23), .ZN(N322) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[4]), .ZN(n101) );
  ND2OPTIBD1BWP30P140 U73 ( .A1(n93), .A2(i_data_bus[36]), .ZN(n24) );
  OAI21D1BWP30P140 U74 ( .A1(n4), .A2(n101), .B(n24), .ZN(N323) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[5]), .ZN(n99) );
  ND2OPTIBD1BWP30P140 U76 ( .A1(n93), .A2(i_data_bus[37]), .ZN(n25) );
  OAI21D1BWP30P140 U77 ( .A1(n4), .A2(n99), .B(n25), .ZN(N324) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[6]), .ZN(n105) );
  ND2OPTIBD1BWP30P140 U79 ( .A1(n93), .A2(i_data_bus[38]), .ZN(n26) );
  OAI21D1BWP30P140 U80 ( .A1(n4), .A2(n105), .B(n26), .ZN(N325) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[7]), .ZN(n97) );
  ND2OPTIBD1BWP30P140 U82 ( .A1(n93), .A2(i_data_bus[39]), .ZN(n27) );
  OAI21D1BWP30P140 U83 ( .A1(n4), .A2(n97), .B(n27), .ZN(N326) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[8]), .ZN(n29) );
  ND2OPTIBD1BWP30P140 U85 ( .A1(n93), .A2(i_data_bus[40]), .ZN(n28) );
  OAI21D1BWP30P140 U86 ( .A1(n4), .A2(n29), .B(n28), .ZN(N327) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[51]), .ZN(n30) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[19]), .ZN(n57) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[50]), .ZN(n31) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[18]), .ZN(n55) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[63]), .ZN(n32) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[31]), .ZN(n81) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[61]), .ZN(n33) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[29]), .ZN(n77) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[49]), .ZN(n34) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[17]), .ZN(n53) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[9]), .ZN(n37) );
  ND2OPTIBD1BWP30P140 U98 ( .A1(n93), .A2(i_data_bus[41]), .ZN(n36) );
  OAI21D1BWP30P140 U99 ( .A1(n4), .A2(n37), .B(n36), .ZN(N328) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[10]), .ZN(n39) );
  ND2OPTIBD1BWP30P140 U101 ( .A1(n93), .A2(i_data_bus[42]), .ZN(n38) );
  OAI21D1BWP30P140 U102 ( .A1(n4), .A2(n39), .B(n38), .ZN(N329) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[11]), .ZN(n41) );
  ND2OPTIBD1BWP30P140 U104 ( .A1(n93), .A2(i_data_bus[43]), .ZN(n40) );
  OAI21D1BWP30P140 U105 ( .A1(n4), .A2(n41), .B(n40), .ZN(N330) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[12]), .ZN(n43) );
  ND2OPTIBD1BWP30P140 U107 ( .A1(n93), .A2(i_data_bus[44]), .ZN(n42) );
  OAI21D1BWP30P140 U108 ( .A1(n4), .A2(n43), .B(n42), .ZN(N331) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[13]), .ZN(n45) );
  ND2OPTIBD1BWP30P140 U110 ( .A1(n93), .A2(i_data_bus[45]), .ZN(n44) );
  OAI21D1BWP30P140 U111 ( .A1(n4), .A2(n45), .B(n44), .ZN(N332) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[14]), .ZN(n47) );
  ND2OPTIBD1BWP30P140 U113 ( .A1(n93), .A2(i_data_bus[46]), .ZN(n46) );
  OAI21D1BWP30P140 U114 ( .A1(n4), .A2(n47), .B(n46), .ZN(N333) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[15]), .ZN(n49) );
  ND2OPTIBD1BWP30P140 U116 ( .A1(n93), .A2(i_data_bus[47]), .ZN(n48) );
  OAI21D1BWP30P140 U117 ( .A1(n4), .A2(n49), .B(n48), .ZN(N334) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[16]), .ZN(n51) );
  ND2OPTIBD1BWP30P140 U119 ( .A1(n93), .A2(i_data_bus[48]), .ZN(n50) );
  OAI21D1BWP30P140 U120 ( .A1(n3), .A2(n51), .B(n50), .ZN(N335) );
  ND2OPTIBD1BWP30P140 U121 ( .A1(n93), .A2(i_data_bus[49]), .ZN(n52) );
  OAI21D1BWP30P140 U122 ( .A1(n3), .A2(n53), .B(n52), .ZN(N336) );
  ND2OPTIBD1BWP30P140 U123 ( .A1(n93), .A2(i_data_bus[50]), .ZN(n54) );
  OAI21D1BWP30P140 U124 ( .A1(n3), .A2(n55), .B(n54), .ZN(N337) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n93), .A2(i_data_bus[51]), .ZN(n56) );
  OAI21D1BWP30P140 U126 ( .A1(n3), .A2(n57), .B(n56), .ZN(N338) );
  INVD1BWP30P140 U127 ( .I(i_data_bus[20]), .ZN(n59) );
  ND2OPTIBD1BWP30P140 U128 ( .A1(n93), .A2(i_data_bus[52]), .ZN(n58) );
  OAI21D1BWP30P140 U129 ( .A1(n3), .A2(n59), .B(n58), .ZN(N339) );
  INVD1BWP30P140 U130 ( .I(i_data_bus[21]), .ZN(n61) );
  OAI21D1BWP30P140 U131 ( .A1(n3), .A2(n61), .B(n60), .ZN(N340) );
  INVD1BWP30P140 U132 ( .I(i_data_bus[22]), .ZN(n63) );
  OAI21D1BWP30P140 U133 ( .A1(n3), .A2(n63), .B(n62), .ZN(N341) );
  INVD1BWP30P140 U134 ( .I(i_data_bus[23]), .ZN(n65) );
  OAI21D1BWP30P140 U135 ( .A1(n3), .A2(n65), .B(n64), .ZN(N342) );
  INVD1BWP30P140 U136 ( .I(i_data_bus[24]), .ZN(n67) );
  OAI21D1BWP30P140 U137 ( .A1(n3), .A2(n67), .B(n66), .ZN(N343) );
  INVD1BWP30P140 U138 ( .I(i_data_bus[25]), .ZN(n69) );
  OAI21D1BWP30P140 U139 ( .A1(n3), .A2(n69), .B(n68), .ZN(N344) );
  INVD1BWP30P140 U140 ( .I(i_data_bus[26]), .ZN(n71) );
  OAI21D1BWP30P140 U141 ( .A1(n3), .A2(n71), .B(n70), .ZN(N345) );
  INVD1BWP30P140 U142 ( .I(i_data_bus[27]), .ZN(n73) );
  OAI21D1BWP30P140 U143 ( .A1(n3), .A2(n73), .B(n72), .ZN(N346) );
  INVD1BWP30P140 U144 ( .I(i_data_bus[28]), .ZN(n75) );
  OAI21D1BWP30P140 U145 ( .A1(n3), .A2(n75), .B(n74), .ZN(N347) );
  OAI21D1BWP30P140 U146 ( .A1(n3), .A2(n77), .B(n76), .ZN(N348) );
  OAI21D1BWP30P140 U147 ( .A1(n3), .A2(n79), .B(n78), .ZN(N349) );
  OAI21D1BWP30P140 U148 ( .A1(n3), .A2(n81), .B(n80), .ZN(N350) );
  INVD1BWP30P140 U149 ( .I(i_data_bus[33]), .ZN(n84) );
  INVD1BWP30P140 U150 ( .I(i_data_bus[32]), .ZN(n86) );
  IND2D1BWP30P140 U151 ( .A1(n106), .B1(i_data_bus[0]), .ZN(n85) );
  OAI21D1BWP30P140 U152 ( .A1(n118), .A2(n86), .B(n85), .ZN(N287) );
  INVD1BWP30P140 U153 ( .I(n92), .ZN(n95) );
  OAI21D1BWP30P140 U154 ( .A1(n95), .A2(i_cmd[1]), .B(n94), .ZN(N354) );
  INVD1BWP30P140 U155 ( .I(i_data_bus[39]), .ZN(n96) );
  INVD1BWP30P140 U156 ( .I(i_data_bus[37]), .ZN(n98) );
  INVD1BWP30P140 U157 ( .I(i_data_bus[36]), .ZN(n100) );
  INVD1BWP30P140 U158 ( .I(i_data_bus[35]), .ZN(n102) );
  INVD1BWP30P140 U159 ( .I(i_data_bus[38]), .ZN(n104) );
  INVD1BWP30P140 U160 ( .I(i_data_bus[60]), .ZN(n107) );
  MOAI22D1BWP30P140 U161 ( .A1(n126), .A2(n107), .B1(n127), .B2(i_data_bus[28]), .ZN(N315) );
  INVD1BWP30P140 U162 ( .I(i_data_bus[48]), .ZN(n108) );
  MOAI22D1BWP30P140 U163 ( .A1(n129), .A2(n108), .B1(n127), .B2(i_data_bus[16]), .ZN(N303) );
  INVD1BWP30P140 U164 ( .I(i_data_bus[34]), .ZN(n109) );
  MOAI22D1BWP30P140 U165 ( .A1(n118), .A2(n109), .B1(n127), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140 U166 ( .I(i_data_bus[59]), .ZN(n110) );
  MOAI22D1BWP30P140 U167 ( .A1(n126), .A2(n110), .B1(n127), .B2(i_data_bus[27]), .ZN(N314) );
  INVD1BWP30P140 U168 ( .I(i_data_bus[47]), .ZN(n111) );
  MOAI22D1BWP30P140 U169 ( .A1(n129), .A2(n111), .B1(n127), .B2(i_data_bus[15]), .ZN(N302) );
  INVD1BWP30P140 U170 ( .I(i_data_bus[58]), .ZN(n112) );
  MOAI22D1BWP30P140 U171 ( .A1(n126), .A2(n112), .B1(n127), .B2(i_data_bus[26]), .ZN(N313) );
  INVD1BWP30P140 U172 ( .I(i_data_bus[46]), .ZN(n113) );
  MOAI22D1BWP30P140 U173 ( .A1(n129), .A2(n113), .B1(n127), .B2(i_data_bus[14]), .ZN(N301) );
  INVD1BWP30P140 U174 ( .I(i_data_bus[57]), .ZN(n114) );
  MOAI22D1BWP30P140 U175 ( .A1(n126), .A2(n114), .B1(n127), .B2(i_data_bus[25]), .ZN(N312) );
  INVD1BWP30P140 U176 ( .I(i_data_bus[45]), .ZN(n115) );
  MOAI22D1BWP30P140 U177 ( .A1(n129), .A2(n115), .B1(n127), .B2(i_data_bus[13]), .ZN(N300) );
  INVD1BWP30P140 U178 ( .I(i_data_bus[56]), .ZN(n116) );
  MOAI22D1BWP30P140 U179 ( .A1(n126), .A2(n116), .B1(n127), .B2(i_data_bus[24]), .ZN(N311) );
  INVD1BWP30P140 U180 ( .I(i_data_bus[44]), .ZN(n117) );
  MOAI22D1BWP30P140 U181 ( .A1(n118), .A2(n117), .B1(n127), .B2(i_data_bus[12]), .ZN(N299) );
  INVD1BWP30P140 U182 ( .I(i_data_bus[55]), .ZN(n119) );
  MOAI22D1BWP30P140 U183 ( .A1(n126), .A2(n119), .B1(n127), .B2(i_data_bus[23]), .ZN(N310) );
  INVD1BWP30P140 U184 ( .I(i_data_bus[43]), .ZN(n120) );
  MOAI22D1BWP30P140 U185 ( .A1(n129), .A2(n120), .B1(n127), .B2(i_data_bus[11]), .ZN(N298) );
  INVD1BWP30P140 U186 ( .I(i_data_bus[54]), .ZN(n121) );
  MOAI22D1BWP30P140 U187 ( .A1(n126), .A2(n121), .B1(n127), .B2(i_data_bus[22]), .ZN(N309) );
  INVD1BWP30P140 U188 ( .I(i_data_bus[42]), .ZN(n122) );
  MOAI22D1BWP30P140 U189 ( .A1(n129), .A2(n122), .B1(n127), .B2(i_data_bus[10]), .ZN(N297) );
  INVD1BWP30P140 U190 ( .I(i_data_bus[53]), .ZN(n123) );
  MOAI22D1BWP30P140 U191 ( .A1(n126), .A2(n123), .B1(n127), .B2(i_data_bus[21]), .ZN(N308) );
  INVD1BWP30P140 U192 ( .I(i_data_bus[41]), .ZN(n124) );
  MOAI22D1BWP30P140 U193 ( .A1(n129), .A2(n124), .B1(n127), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140 U194 ( .I(i_data_bus[52]), .ZN(n125) );
  MOAI22D1BWP30P140 U195 ( .A1(n126), .A2(n125), .B1(n127), .B2(i_data_bus[20]), .ZN(N307) );
  INVD1BWP30P140 U196 ( .I(i_data_bus[40]), .ZN(n128) );
  MOAI22D1BWP30P140 U197 ( .A1(n129), .A2(n128), .B1(n127), .B2(i_data_bus[8]), 
        .ZN(N295) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_51 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  INVD3BWP30P140 U3 ( .I(n17), .ZN(n105) );
  NR2D4BWP30P140 U4 ( .A1(n13), .A2(n12), .ZN(n17) );
  NR2D1BWP30P140 U5 ( .A1(i_cmd[1]), .A2(n91), .ZN(n24) );
  INVD6BWP30P140 U6 ( .I(n39), .ZN(n1) );
  ND2OPTPAD1BWP30P140 U7 ( .A1(i_cmd[0]), .A2(n11), .ZN(n12) );
  AN2D1BWP30P140 U8 ( .A1(i_valid[0]), .A2(n11), .Z(n8) );
  MUX2NOPTD2BWP30P140 U9 ( .I0(i_valid[0]), .I1(i_valid[1]), .S(i_cmd[1]), 
        .ZN(n13) );
  MUX2NOPTD2BWP30P140 U10 ( .I0(i_valid[0]), .I1(i_valid[1]), .S(i_cmd[0]), 
        .ZN(n23) );
  OR2D8BWP30P140 U11 ( .A1(n14), .A2(i_cmd[0]), .Z(n107) );
  CKND2D4BWP30P140 U12 ( .A1(i_valid[0]), .A2(n11), .ZN(n14) );
  INVD2BWP30P140 U13 ( .I(n107), .ZN(n9) );
  INVD8BWP30P140 U14 ( .I(n107), .ZN(n126) );
  INVD1BWP30P140 U15 ( .I(i_cmd[0]), .ZN(n94) );
  ND3OPTPAD2BWP30P140 U16 ( .A1(i_cmd[1]), .A2(i_valid[1]), .A3(n11), .ZN(n96)
         );
  ND2D1BWP30P140 U17 ( .A1(n10), .A2(i_en), .ZN(n91) );
  ND2D1BWP30P140 U18 ( .A1(n107), .A2(n95), .ZN(N353) );
  IND2D1BWP30P140 U19 ( .A1(n94), .B1(n93), .ZN(n95) );
  NR2D1BWP30P140 U20 ( .A1(n92), .A2(n91), .ZN(n93) );
  INVD1BWP30P140 U21 ( .I(i_valid[1]), .ZN(n92) );
  OAI21D1BWP30P140 U22 ( .A1(n105), .A2(n90), .B(n89), .ZN(N287) );
  OAI21D1BWP30P140 U23 ( .A1(n105), .A2(n88), .B(n87), .ZN(N288) );
  ND2D1BWP30P140 U24 ( .A1(n9), .A2(i_data_bus[1]), .ZN(n87) );
  ND2D1BWP30P140 U25 ( .A1(n84), .A2(i_data_bus[47]), .ZN(n52) );
  ND2D1BWP30P140 U26 ( .A1(n84), .A2(i_data_bus[51]), .ZN(n60) );
  ND2D1BWP30P140 U27 ( .A1(n84), .A2(i_data_bus[52]), .ZN(n62) );
  ND2D1BWP30P140 U28 ( .A1(n84), .A2(i_data_bus[53]), .ZN(n64) );
  ND2D1BWP30P140 U29 ( .A1(n84), .A2(i_data_bus[54]), .ZN(n66) );
  ND2D1BWP30P140 U30 ( .A1(n84), .A2(i_data_bus[55]), .ZN(n68) );
  ND2D1BWP30P140 U31 ( .A1(n84), .A2(i_data_bus[56]), .ZN(n70) );
  ND2D1BWP30P140 U32 ( .A1(n84), .A2(i_data_bus[57]), .ZN(n72) );
  ND2D1BWP30P140 U33 ( .A1(n84), .A2(i_data_bus[58]), .ZN(n74) );
  ND2D1BWP30P140 U34 ( .A1(n84), .A2(i_data_bus[59]), .ZN(n76) );
  ND2D1BWP30P140 U35 ( .A1(n84), .A2(i_data_bus[60]), .ZN(n78) );
  ND2D1BWP30P140 U36 ( .A1(n84), .A2(i_data_bus[61]), .ZN(n80) );
  ND2D1BWP30P140 U37 ( .A1(n84), .A2(i_data_bus[62]), .ZN(n82) );
  ND2D1BWP30P140 U38 ( .A1(n84), .A2(i_data_bus[63]), .ZN(n85) );
  OAI22D1BWP30P140 U39 ( .A1(n128), .A2(n22), .B1(n107), .B2(n61), .ZN(N306)
         );
  OAI22D1BWP30P140 U40 ( .A1(n128), .A2(n21), .B1(n107), .B2(n57), .ZN(N304)
         );
  OAI22D1BWP30P140 U41 ( .A1(n128), .A2(n20), .B1(n107), .B2(n81), .ZN(N316)
         );
  OAI22D1BWP30P140 U42 ( .A1(n128), .A2(n19), .B1(n107), .B2(n83), .ZN(N317)
         );
  OAI22D1BWP30P140 U43 ( .A1(n107), .A2(n32), .B1(n105), .B2(n18), .ZN(N290)
         );
  INR2D4BWP30P140 U44 ( .A1(n24), .B1(n23), .ZN(n39) );
  INVD1BWP30P140 U45 ( .I(n91), .ZN(n11) );
  INVD1BWP30P140 U46 ( .I(rst), .ZN(n10) );
  INVD6BWP30P140 U47 ( .I(n17), .ZN(n128) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[63]), .ZN(n15) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[31]), .ZN(n86) );
  OAI22D1BWP30P140 U50 ( .A1(n128), .A2(n15), .B1(n107), .B2(n86), .ZN(N318)
         );
  INVD1BWP30P140 U51 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[18]), .ZN(n59) );
  OAI22D1BWP30P140 U53 ( .A1(n128), .A2(n16), .B1(n107), .B2(n59), .ZN(N305)
         );
  INVD1BWP30P140 U54 ( .I(i_data_bus[3]), .ZN(n32) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[35]), .ZN(n18) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[62]), .ZN(n19) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[30]), .ZN(n83) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[61]), .ZN(n20) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[29]), .ZN(n81) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[49]), .ZN(n21) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[17]), .ZN(n57) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[51]), .ZN(n22) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[19]), .ZN(n61) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[0]), .ZN(n26) );
  INVD6BWP30P140 U65 ( .I(n96), .ZN(n84) );
  ND2OPTIBD1BWP30P140 U66 ( .A1(n84), .A2(i_data_bus[32]), .ZN(n25) );
  OAI21D1BWP30P140 U67 ( .A1(n1), .A2(n26), .B(n25), .ZN(N319) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[1]), .ZN(n28) );
  ND2OPTIBD1BWP30P140 U69 ( .A1(n84), .A2(i_data_bus[33]), .ZN(n27) );
  OAI21D1BWP30P140 U70 ( .A1(n1), .A2(n28), .B(n27), .ZN(N320) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[2]), .ZN(n30) );
  ND2OPTIBD1BWP30P140 U72 ( .A1(n84), .A2(i_data_bus[34]), .ZN(n29) );
  OAI21D1BWP30P140 U73 ( .A1(n1), .A2(n30), .B(n29), .ZN(N321) );
  ND2OPTIBD1BWP30P140 U74 ( .A1(n84), .A2(i_data_bus[35]), .ZN(n31) );
  OAI21D1BWP30P140 U75 ( .A1(n1), .A2(n32), .B(n31), .ZN(N322) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[4]), .ZN(n99) );
  ND2OPTIBD1BWP30P140 U77 ( .A1(n84), .A2(i_data_bus[36]), .ZN(n33) );
  OAI21D1BWP30P140 U78 ( .A1(n1), .A2(n99), .B(n33), .ZN(N323) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[5]), .ZN(n103) );
  ND2OPTIBD1BWP30P140 U80 ( .A1(n84), .A2(i_data_bus[37]), .ZN(n34) );
  OAI21D1BWP30P140 U81 ( .A1(n1), .A2(n103), .B(n34), .ZN(N324) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[6]), .ZN(n101) );
  ND2OPTIBD1BWP30P140 U83 ( .A1(n84), .A2(i_data_bus[38]), .ZN(n35) );
  OAI21D1BWP30P140 U84 ( .A1(n1), .A2(n101), .B(n35), .ZN(N325) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[7]), .ZN(n106) );
  ND2OPTIBD1BWP30P140 U86 ( .A1(n84), .A2(i_data_bus[39]), .ZN(n36) );
  OAI21D1BWP30P140 U87 ( .A1(n1), .A2(n106), .B(n36), .ZN(N326) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[8]), .ZN(n38) );
  ND2OPTIBD1BWP30P140 U89 ( .A1(n84), .A2(i_data_bus[40]), .ZN(n37) );
  OAI21D1BWP30P140 U90 ( .A1(n1), .A2(n38), .B(n37), .ZN(N327) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[9]), .ZN(n41) );
  ND2OPTIBD1BWP30P140 U92 ( .A1(n84), .A2(i_data_bus[41]), .ZN(n40) );
  OAI21D1BWP30P140 U93 ( .A1(n1), .A2(n41), .B(n40), .ZN(N328) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[10]), .ZN(n43) );
  ND2OPTIBD1BWP30P140 U95 ( .A1(n84), .A2(i_data_bus[42]), .ZN(n42) );
  OAI21D1BWP30P140 U96 ( .A1(n1), .A2(n43), .B(n42), .ZN(N329) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[11]), .ZN(n45) );
  ND2OPTIBD1BWP30P140 U98 ( .A1(n84), .A2(i_data_bus[43]), .ZN(n44) );
  OAI21D1BWP30P140 U99 ( .A1(n1), .A2(n45), .B(n44), .ZN(N330) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[12]), .ZN(n47) );
  ND2OPTIBD1BWP30P140 U101 ( .A1(n84), .A2(i_data_bus[44]), .ZN(n46) );
  OAI21D1BWP30P140 U102 ( .A1(n1), .A2(n47), .B(n46), .ZN(N331) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[13]), .ZN(n49) );
  ND2OPTIBD1BWP30P140 U104 ( .A1(n84), .A2(i_data_bus[45]), .ZN(n48) );
  OAI21D1BWP30P140 U105 ( .A1(n1), .A2(n49), .B(n48), .ZN(N332) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[14]), .ZN(n51) );
  ND2OPTIBD1BWP30P140 U107 ( .A1(n84), .A2(i_data_bus[46]), .ZN(n50) );
  OAI21D1BWP30P140 U108 ( .A1(n1), .A2(n51), .B(n50), .ZN(N333) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[15]), .ZN(n53) );
  OAI21D1BWP30P140 U110 ( .A1(n1), .A2(n53), .B(n52), .ZN(N334) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[16]), .ZN(n55) );
  ND2OPTIBD1BWP30P140 U112 ( .A1(n84), .A2(i_data_bus[48]), .ZN(n54) );
  OAI21D1BWP30P140 U113 ( .A1(n1), .A2(n55), .B(n54), .ZN(N335) );
  ND2OPTIBD1BWP30P140 U114 ( .A1(n84), .A2(i_data_bus[49]), .ZN(n56) );
  OAI21D1BWP30P140 U115 ( .A1(n1), .A2(n57), .B(n56), .ZN(N336) );
  ND2OPTIBD1BWP30P140 U116 ( .A1(n84), .A2(i_data_bus[50]), .ZN(n58) );
  OAI21D1BWP30P140 U117 ( .A1(n1), .A2(n59), .B(n58), .ZN(N337) );
  OAI21D1BWP30P140 U118 ( .A1(n1), .A2(n61), .B(n60), .ZN(N338) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[20]), .ZN(n63) );
  OAI21D1BWP30P140 U120 ( .A1(n1), .A2(n63), .B(n62), .ZN(N339) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[21]), .ZN(n65) );
  OAI21D1BWP30P140 U122 ( .A1(n1), .A2(n65), .B(n64), .ZN(N340) );
  INVD1BWP30P140 U123 ( .I(i_data_bus[22]), .ZN(n67) );
  OAI21D1BWP30P140 U124 ( .A1(n1), .A2(n67), .B(n66), .ZN(N341) );
  INVD1BWP30P140 U125 ( .I(i_data_bus[23]), .ZN(n69) );
  OAI21D1BWP30P140 U126 ( .A1(n1), .A2(n69), .B(n68), .ZN(N342) );
  INVD1BWP30P140 U127 ( .I(i_data_bus[24]), .ZN(n71) );
  OAI21D1BWP30P140 U128 ( .A1(n1), .A2(n71), .B(n70), .ZN(N343) );
  INVD1BWP30P140 U129 ( .I(i_data_bus[25]), .ZN(n73) );
  OAI21D1BWP30P140 U130 ( .A1(n1), .A2(n73), .B(n72), .ZN(N344) );
  INVD1BWP30P140 U131 ( .I(i_data_bus[26]), .ZN(n75) );
  OAI21D1BWP30P140 U132 ( .A1(n1), .A2(n75), .B(n74), .ZN(N345) );
  INVD1BWP30P140 U133 ( .I(i_data_bus[27]), .ZN(n77) );
  OAI21D1BWP30P140 U134 ( .A1(n1), .A2(n77), .B(n76), .ZN(N346) );
  INVD1BWP30P140 U135 ( .I(i_data_bus[28]), .ZN(n79) );
  OAI21D1BWP30P140 U136 ( .A1(n1), .A2(n79), .B(n78), .ZN(N347) );
  OAI21D1BWP30P140 U137 ( .A1(n1), .A2(n81), .B(n80), .ZN(N348) );
  OAI21D1BWP30P140 U138 ( .A1(n1), .A2(n83), .B(n82), .ZN(N349) );
  OAI21D1BWP30P140 U139 ( .A1(n1), .A2(n86), .B(n85), .ZN(N350) );
  INVD1BWP30P140 U140 ( .I(i_data_bus[33]), .ZN(n88) );
  INVD1BWP30P140 U141 ( .I(i_data_bus[32]), .ZN(n90) );
  IND2D2BWP30P140 U142 ( .A1(n107), .B1(i_data_bus[0]), .ZN(n89) );
  INVD1BWP30P140 U143 ( .I(n8), .ZN(n97) );
  OAI21D1BWP30P140 U144 ( .A1(n97), .A2(i_cmd[1]), .B(n96), .ZN(N354) );
  INVD1BWP30P140 U145 ( .I(i_data_bus[36]), .ZN(n98) );
  OAI22D1BWP30P140 U146 ( .A1(n107), .A2(n99), .B1(n105), .B2(n98), .ZN(N291)
         );
  INVD1BWP30P140 U147 ( .I(i_data_bus[38]), .ZN(n100) );
  OAI22D1BWP30P140 U148 ( .A1(n107), .A2(n101), .B1(n105), .B2(n100), .ZN(N293) );
  INVD1BWP30P140 U149 ( .I(i_data_bus[37]), .ZN(n102) );
  OAI22D1BWP30P140 U150 ( .A1(n107), .A2(n103), .B1(n105), .B2(n102), .ZN(N292) );
  INVD1BWP30P140 U151 ( .I(i_data_bus[39]), .ZN(n104) );
  OAI22D1BWP30P140 U152 ( .A1(n107), .A2(n106), .B1(n105), .B2(n104), .ZN(N294) );
  INVD1BWP30P140 U153 ( .I(i_data_bus[60]), .ZN(n108) );
  MOAI22D1BWP30P140 U154 ( .A1(n128), .A2(n108), .B1(n126), .B2(i_data_bus[28]), .ZN(N315) );
  INVD1BWP30P140 U155 ( .I(i_data_bus[48]), .ZN(n109) );
  MOAI22D1BWP30P140 U156 ( .A1(n128), .A2(n109), .B1(n126), .B2(i_data_bus[16]), .ZN(N303) );
  INVD1BWP30P140 U157 ( .I(i_data_bus[34]), .ZN(n110) );
  MOAI22D1BWP30P140 U158 ( .A1(n128), .A2(n110), .B1(n126), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140 U159 ( .I(i_data_bus[59]), .ZN(n111) );
  MOAI22D1BWP30P140 U160 ( .A1(n128), .A2(n111), .B1(n126), .B2(i_data_bus[27]), .ZN(N314) );
  INVD1BWP30P140 U161 ( .I(i_data_bus[47]), .ZN(n112) );
  MOAI22D1BWP30P140 U162 ( .A1(n128), .A2(n112), .B1(n126), .B2(i_data_bus[15]), .ZN(N302) );
  INVD1BWP30P140 U163 ( .I(i_data_bus[58]), .ZN(n113) );
  MOAI22D1BWP30P140 U164 ( .A1(n128), .A2(n113), .B1(n126), .B2(i_data_bus[26]), .ZN(N313) );
  INVD1BWP30P140 U165 ( .I(i_data_bus[46]), .ZN(n114) );
  MOAI22D1BWP30P140 U166 ( .A1(n128), .A2(n114), .B1(n126), .B2(i_data_bus[14]), .ZN(N301) );
  INVD1BWP30P140 U167 ( .I(i_data_bus[57]), .ZN(n115) );
  MOAI22D1BWP30P140 U168 ( .A1(n128), .A2(n115), .B1(n126), .B2(i_data_bus[25]), .ZN(N312) );
  INVD1BWP30P140 U169 ( .I(i_data_bus[45]), .ZN(n116) );
  MOAI22D1BWP30P140 U170 ( .A1(n128), .A2(n116), .B1(n126), .B2(i_data_bus[13]), .ZN(N300) );
  INVD1BWP30P140 U171 ( .I(i_data_bus[56]), .ZN(n117) );
  MOAI22D1BWP30P140 U172 ( .A1(n128), .A2(n117), .B1(n126), .B2(i_data_bus[24]), .ZN(N311) );
  INVD1BWP30P140 U173 ( .I(i_data_bus[44]), .ZN(n118) );
  MOAI22D1BWP30P140 U174 ( .A1(n128), .A2(n118), .B1(n126), .B2(i_data_bus[12]), .ZN(N299) );
  INVD1BWP30P140 U175 ( .I(i_data_bus[55]), .ZN(n119) );
  MOAI22D1BWP30P140 U176 ( .A1(n128), .A2(n119), .B1(n126), .B2(i_data_bus[23]), .ZN(N310) );
  INVD1BWP30P140 U177 ( .I(i_data_bus[43]), .ZN(n120) );
  MOAI22D1BWP30P140 U178 ( .A1(n128), .A2(n120), .B1(n126), .B2(i_data_bus[11]), .ZN(N298) );
  INVD1BWP30P140 U179 ( .I(i_data_bus[54]), .ZN(n121) );
  MOAI22D1BWP30P140 U180 ( .A1(n128), .A2(n121), .B1(n126), .B2(i_data_bus[22]), .ZN(N309) );
  INVD1BWP30P140 U181 ( .I(i_data_bus[42]), .ZN(n122) );
  MOAI22D1BWP30P140 U182 ( .A1(n128), .A2(n122), .B1(n126), .B2(i_data_bus[10]), .ZN(N297) );
  INVD1BWP30P140 U183 ( .I(i_data_bus[53]), .ZN(n123) );
  MOAI22D1BWP30P140 U184 ( .A1(n128), .A2(n123), .B1(n126), .B2(i_data_bus[21]), .ZN(N308) );
  INVD1BWP30P140 U185 ( .I(i_data_bus[41]), .ZN(n124) );
  MOAI22D1BWP30P140 U186 ( .A1(n128), .A2(n124), .B1(n126), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140 U187 ( .I(i_data_bus[52]), .ZN(n125) );
  MOAI22D1BWP30P140 U188 ( .A1(n128), .A2(n125), .B1(n126), .B2(i_data_bus[20]), .ZN(N307) );
  INVD1BWP30P140 U189 ( .I(i_data_bus[40]), .ZN(n127) );
  MOAI22D1BWP30P140 U190 ( .A1(n128), .A2(n127), .B1(n9), .B2(i_data_bus[8]), 
        .ZN(N295) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_52 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  INVD3BWP30P140 U3 ( .I(n17), .ZN(n105) );
  NR2D4BWP30P140 U4 ( .A1(n13), .A2(n12), .ZN(n17) );
  NR2D1BWP30P140 U5 ( .A1(i_cmd[1]), .A2(n91), .ZN(n24) );
  INVD6BWP30P140 U6 ( .I(n35), .ZN(n1) );
  ND2OPTPAD1BWP30P140 U7 ( .A1(i_cmd[0]), .A2(n11), .ZN(n12) );
  AN2D1BWP30P140 U8 ( .A1(i_valid[0]), .A2(n11), .Z(n8) );
  MUX2NOPTD2BWP30P140 U9 ( .I0(i_valid[0]), .I1(i_valid[1]), .S(i_cmd[1]), 
        .ZN(n13) );
  MUX2NOPTD2BWP30P140 U10 ( .I0(i_valid[0]), .I1(i_valid[1]), .S(i_cmd[0]), 
        .ZN(n23) );
  OR2D8BWP30P140 U11 ( .A1(n14), .A2(i_cmd[0]), .Z(n107) );
  CKND2D4BWP30P140 U12 ( .A1(i_valid[0]), .A2(n11), .ZN(n14) );
  INVD2BWP30P140 U13 ( .I(n107), .ZN(n9) );
  INVD8BWP30P140 U14 ( .I(n107), .ZN(n126) );
  INVD1BWP30P140 U15 ( .I(i_cmd[0]), .ZN(n94) );
  ND3OPTPAD2BWP30P140 U16 ( .A1(i_cmd[1]), .A2(i_valid[1]), .A3(n11), .ZN(n96)
         );
  ND2D1BWP30P140 U17 ( .A1(n10), .A2(i_en), .ZN(n91) );
  ND2D1BWP30P140 U18 ( .A1(n107), .A2(n95), .ZN(N353) );
  IND2D1BWP30P140 U19 ( .A1(n94), .B1(n93), .ZN(n95) );
  NR2D1BWP30P140 U20 ( .A1(n92), .A2(n91), .ZN(n93) );
  INVD1BWP30P140 U21 ( .I(i_valid[1]), .ZN(n92) );
  OAI21D1BWP30P140 U22 ( .A1(n105), .A2(n90), .B(n89), .ZN(N287) );
  OAI21D1BWP30P140 U23 ( .A1(n105), .A2(n88), .B(n87), .ZN(N288) );
  ND2D1BWP30P140 U24 ( .A1(n9), .A2(i_data_bus[1]), .ZN(n87) );
  ND2D1BWP30P140 U25 ( .A1(n84), .A2(i_data_bus[47]), .ZN(n48) );
  ND2D1BWP30P140 U26 ( .A1(n84), .A2(i_data_bus[51]), .ZN(n56) );
  ND2D1BWP30P140 U27 ( .A1(n84), .A2(i_data_bus[52]), .ZN(n58) );
  ND2D1BWP30P140 U28 ( .A1(n84), .A2(i_data_bus[53]), .ZN(n60) );
  ND2D1BWP30P140 U29 ( .A1(n84), .A2(i_data_bus[54]), .ZN(n62) );
  ND2D1BWP30P140 U30 ( .A1(n84), .A2(i_data_bus[55]), .ZN(n64) );
  ND2D1BWP30P140 U31 ( .A1(n84), .A2(i_data_bus[56]), .ZN(n66) );
  ND2D1BWP30P140 U32 ( .A1(n84), .A2(i_data_bus[57]), .ZN(n68) );
  ND2D1BWP30P140 U33 ( .A1(n84), .A2(i_data_bus[58]), .ZN(n70) );
  ND2D1BWP30P140 U34 ( .A1(n84), .A2(i_data_bus[59]), .ZN(n72) );
  ND2D1BWP30P140 U35 ( .A1(n84), .A2(i_data_bus[60]), .ZN(n74) );
  ND2D1BWP30P140 U36 ( .A1(n84), .A2(i_data_bus[61]), .ZN(n76) );
  ND2D1BWP30P140 U37 ( .A1(n84), .A2(i_data_bus[62]), .ZN(n78) );
  ND2D1BWP30P140 U38 ( .A1(n84), .A2(i_data_bus[63]), .ZN(n80) );
  OAI22D1BWP30P140 U39 ( .A1(n128), .A2(n22), .B1(n107), .B2(n79), .ZN(N317)
         );
  OAI22D1BWP30P140 U40 ( .A1(n128), .A2(n21), .B1(n107), .B2(n77), .ZN(N316)
         );
  OAI22D1BWP30P140 U41 ( .A1(n128), .A2(n20), .B1(n107), .B2(n57), .ZN(N306)
         );
  OAI22D1BWP30P140 U42 ( .A1(n128), .A2(n19), .B1(n107), .B2(n53), .ZN(N304)
         );
  OAI22D1BWP30P140 U43 ( .A1(n107), .A2(n31), .B1(n105), .B2(n18), .ZN(N293)
         );
  INR2D4BWP30P140 U44 ( .A1(n24), .B1(n23), .ZN(n35) );
  INVD1BWP30P140 U45 ( .I(n91), .ZN(n11) );
  INVD1BWP30P140 U46 ( .I(rst), .ZN(n10) );
  INVD6BWP30P140 U47 ( .I(n17), .ZN(n128) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[50]), .ZN(n15) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[18]), .ZN(n55) );
  OAI22D1BWP30P140 U50 ( .A1(n128), .A2(n15), .B1(n107), .B2(n55), .ZN(N305)
         );
  INVD1BWP30P140 U51 ( .I(i_data_bus[63]), .ZN(n16) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[31]), .ZN(n81) );
  OAI22D1BWP30P140 U53 ( .A1(n128), .A2(n16), .B1(n107), .B2(n81), .ZN(N318)
         );
  INVD1BWP30P140 U54 ( .I(i_data_bus[6]), .ZN(n31) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[38]), .ZN(n18) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[49]), .ZN(n19) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[17]), .ZN(n53) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[51]), .ZN(n20) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[19]), .ZN(n57) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[61]), .ZN(n21) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[29]), .ZN(n77) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[62]), .ZN(n22) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[30]), .ZN(n79) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[2]), .ZN(n26) );
  INVD6BWP30P140 U65 ( .I(n96), .ZN(n84) );
  ND2OPTIBD1BWP30P140 U66 ( .A1(n84), .A2(i_data_bus[34]), .ZN(n25) );
  OAI21D1BWP30P140 U67 ( .A1(n1), .A2(n26), .B(n25), .ZN(N321) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[3]), .ZN(n99) );
  ND2OPTIBD1BWP30P140 U69 ( .A1(n84), .A2(i_data_bus[35]), .ZN(n27) );
  OAI21D1BWP30P140 U70 ( .A1(n1), .A2(n99), .B(n27), .ZN(N322) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[4]), .ZN(n103) );
  ND2OPTIBD1BWP30P140 U72 ( .A1(n84), .A2(i_data_bus[36]), .ZN(n28) );
  OAI21D1BWP30P140 U73 ( .A1(n1), .A2(n103), .B(n28), .ZN(N323) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[5]), .ZN(n106) );
  ND2OPTIBD1BWP30P140 U75 ( .A1(n84), .A2(i_data_bus[37]), .ZN(n29) );
  OAI21D1BWP30P140 U76 ( .A1(n1), .A2(n106), .B(n29), .ZN(N324) );
  ND2OPTIBD1BWP30P140 U77 ( .A1(n84), .A2(i_data_bus[38]), .ZN(n30) );
  OAI21D1BWP30P140 U78 ( .A1(n1), .A2(n31), .B(n30), .ZN(N325) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[7]), .ZN(n101) );
  ND2OPTIBD1BWP30P140 U80 ( .A1(n84), .A2(i_data_bus[39]), .ZN(n32) );
  OAI21D1BWP30P140 U81 ( .A1(n1), .A2(n101), .B(n32), .ZN(N326) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[8]), .ZN(n34) );
  ND2OPTIBD1BWP30P140 U83 ( .A1(n84), .A2(i_data_bus[40]), .ZN(n33) );
  OAI21D1BWP30P140 U84 ( .A1(n1), .A2(n34), .B(n33), .ZN(N327) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[9]), .ZN(n37) );
  ND2OPTIBD1BWP30P140 U86 ( .A1(n84), .A2(i_data_bus[41]), .ZN(n36) );
  OAI21D1BWP30P140 U87 ( .A1(n1), .A2(n37), .B(n36), .ZN(N328) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[10]), .ZN(n39) );
  ND2OPTIBD1BWP30P140 U89 ( .A1(n84), .A2(i_data_bus[42]), .ZN(n38) );
  OAI21D1BWP30P140 U90 ( .A1(n1), .A2(n39), .B(n38), .ZN(N329) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[11]), .ZN(n41) );
  ND2OPTIBD1BWP30P140 U92 ( .A1(n84), .A2(i_data_bus[43]), .ZN(n40) );
  OAI21D1BWP30P140 U93 ( .A1(n1), .A2(n41), .B(n40), .ZN(N330) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[12]), .ZN(n43) );
  ND2OPTIBD1BWP30P140 U95 ( .A1(n84), .A2(i_data_bus[44]), .ZN(n42) );
  OAI21D1BWP30P140 U96 ( .A1(n1), .A2(n43), .B(n42), .ZN(N331) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[13]), .ZN(n45) );
  ND2OPTIBD1BWP30P140 U98 ( .A1(n84), .A2(i_data_bus[45]), .ZN(n44) );
  OAI21D1BWP30P140 U99 ( .A1(n1), .A2(n45), .B(n44), .ZN(N332) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[14]), .ZN(n47) );
  ND2OPTIBD1BWP30P140 U101 ( .A1(n84), .A2(i_data_bus[46]), .ZN(n46) );
  OAI21D1BWP30P140 U102 ( .A1(n1), .A2(n47), .B(n46), .ZN(N333) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[15]), .ZN(n49) );
  OAI21D1BWP30P140 U104 ( .A1(n1), .A2(n49), .B(n48), .ZN(N334) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[16]), .ZN(n51) );
  ND2OPTIBD1BWP30P140 U106 ( .A1(n84), .A2(i_data_bus[48]), .ZN(n50) );
  OAI21D1BWP30P140 U107 ( .A1(n1), .A2(n51), .B(n50), .ZN(N335) );
  ND2OPTIBD1BWP30P140 U108 ( .A1(n84), .A2(i_data_bus[49]), .ZN(n52) );
  OAI21D1BWP30P140 U109 ( .A1(n1), .A2(n53), .B(n52), .ZN(N336) );
  ND2OPTIBD1BWP30P140 U110 ( .A1(n84), .A2(i_data_bus[50]), .ZN(n54) );
  OAI21D1BWP30P140 U111 ( .A1(n1), .A2(n55), .B(n54), .ZN(N337) );
  OAI21D1BWP30P140 U112 ( .A1(n1), .A2(n57), .B(n56), .ZN(N338) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[20]), .ZN(n59) );
  OAI21D1BWP30P140 U114 ( .A1(n1), .A2(n59), .B(n58), .ZN(N339) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[21]), .ZN(n61) );
  OAI21D1BWP30P140 U116 ( .A1(n1), .A2(n61), .B(n60), .ZN(N340) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[22]), .ZN(n63) );
  OAI21D1BWP30P140 U118 ( .A1(n1), .A2(n63), .B(n62), .ZN(N341) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[23]), .ZN(n65) );
  OAI21D1BWP30P140 U120 ( .A1(n1), .A2(n65), .B(n64), .ZN(N342) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[24]), .ZN(n67) );
  OAI21D1BWP30P140 U122 ( .A1(n1), .A2(n67), .B(n66), .ZN(N343) );
  INVD1BWP30P140 U123 ( .I(i_data_bus[25]), .ZN(n69) );
  OAI21D1BWP30P140 U124 ( .A1(n1), .A2(n69), .B(n68), .ZN(N344) );
  INVD1BWP30P140 U125 ( .I(i_data_bus[26]), .ZN(n71) );
  OAI21D1BWP30P140 U126 ( .A1(n1), .A2(n71), .B(n70), .ZN(N345) );
  INVD1BWP30P140 U127 ( .I(i_data_bus[27]), .ZN(n73) );
  OAI21D1BWP30P140 U128 ( .A1(n1), .A2(n73), .B(n72), .ZN(N346) );
  INVD1BWP30P140 U129 ( .I(i_data_bus[28]), .ZN(n75) );
  OAI21D1BWP30P140 U130 ( .A1(n1), .A2(n75), .B(n74), .ZN(N347) );
  OAI21D1BWP30P140 U131 ( .A1(n1), .A2(n77), .B(n76), .ZN(N348) );
  OAI21D1BWP30P140 U132 ( .A1(n1), .A2(n79), .B(n78), .ZN(N349) );
  OAI21D1BWP30P140 U133 ( .A1(n1), .A2(n81), .B(n80), .ZN(N350) );
  INVD1BWP30P140 U134 ( .I(i_data_bus[1]), .ZN(n83) );
  ND2OPTIBD1BWP30P140 U135 ( .A1(n84), .A2(i_data_bus[33]), .ZN(n82) );
  OAI21D1BWP30P140 U136 ( .A1(n1), .A2(n83), .B(n82), .ZN(N320) );
  INVD1BWP30P140 U137 ( .I(i_data_bus[0]), .ZN(n86) );
  ND2OPTIBD1BWP30P140 U138 ( .A1(n84), .A2(i_data_bus[32]), .ZN(n85) );
  OAI21D1BWP30P140 U139 ( .A1(n1), .A2(n86), .B(n85), .ZN(N319) );
  INVD1BWP30P140 U140 ( .I(i_data_bus[33]), .ZN(n88) );
  INVD1BWP30P140 U141 ( .I(i_data_bus[32]), .ZN(n90) );
  IND2D2BWP30P140 U142 ( .A1(n107), .B1(i_data_bus[0]), .ZN(n89) );
  INVD1BWP30P140 U143 ( .I(n8), .ZN(n97) );
  OAI21D1BWP30P140 U144 ( .A1(n97), .A2(i_cmd[1]), .B(n96), .ZN(N354) );
  INVD1BWP30P140 U145 ( .I(i_data_bus[35]), .ZN(n98) );
  OAI22D1BWP30P140 U146 ( .A1(n107), .A2(n99), .B1(n105), .B2(n98), .ZN(N290)
         );
  INVD1BWP30P140 U147 ( .I(i_data_bus[39]), .ZN(n100) );
  OAI22D1BWP30P140 U148 ( .A1(n107), .A2(n101), .B1(n105), .B2(n100), .ZN(N294) );
  INVD1BWP30P140 U149 ( .I(i_data_bus[36]), .ZN(n102) );
  OAI22D1BWP30P140 U150 ( .A1(n107), .A2(n103), .B1(n105), .B2(n102), .ZN(N291) );
  INVD1BWP30P140 U151 ( .I(i_data_bus[37]), .ZN(n104) );
  OAI22D1BWP30P140 U152 ( .A1(n107), .A2(n106), .B1(n105), .B2(n104), .ZN(N292) );
  INVD1BWP30P140 U153 ( .I(i_data_bus[60]), .ZN(n108) );
  MOAI22D1BWP30P140 U154 ( .A1(n128), .A2(n108), .B1(n126), .B2(i_data_bus[28]), .ZN(N315) );
  INVD1BWP30P140 U155 ( .I(i_data_bus[48]), .ZN(n109) );
  MOAI22D1BWP30P140 U156 ( .A1(n128), .A2(n109), .B1(n126), .B2(i_data_bus[16]), .ZN(N303) );
  INVD1BWP30P140 U157 ( .I(i_data_bus[34]), .ZN(n110) );
  MOAI22D1BWP30P140 U158 ( .A1(n128), .A2(n110), .B1(n126), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140 U159 ( .I(i_data_bus[59]), .ZN(n111) );
  MOAI22D1BWP30P140 U160 ( .A1(n128), .A2(n111), .B1(n126), .B2(i_data_bus[27]), .ZN(N314) );
  INVD1BWP30P140 U161 ( .I(i_data_bus[47]), .ZN(n112) );
  MOAI22D1BWP30P140 U162 ( .A1(n128), .A2(n112), .B1(n126), .B2(i_data_bus[15]), .ZN(N302) );
  INVD1BWP30P140 U163 ( .I(i_data_bus[58]), .ZN(n113) );
  MOAI22D1BWP30P140 U164 ( .A1(n128), .A2(n113), .B1(n126), .B2(i_data_bus[26]), .ZN(N313) );
  INVD1BWP30P140 U165 ( .I(i_data_bus[46]), .ZN(n114) );
  MOAI22D1BWP30P140 U166 ( .A1(n128), .A2(n114), .B1(n126), .B2(i_data_bus[14]), .ZN(N301) );
  INVD1BWP30P140 U167 ( .I(i_data_bus[57]), .ZN(n115) );
  MOAI22D1BWP30P140 U168 ( .A1(n128), .A2(n115), .B1(n126), .B2(i_data_bus[25]), .ZN(N312) );
  INVD1BWP30P140 U169 ( .I(i_data_bus[45]), .ZN(n116) );
  MOAI22D1BWP30P140 U170 ( .A1(n128), .A2(n116), .B1(n126), .B2(i_data_bus[13]), .ZN(N300) );
  INVD1BWP30P140 U171 ( .I(i_data_bus[56]), .ZN(n117) );
  MOAI22D1BWP30P140 U172 ( .A1(n128), .A2(n117), .B1(n126), .B2(i_data_bus[24]), .ZN(N311) );
  INVD1BWP30P140 U173 ( .I(i_data_bus[44]), .ZN(n118) );
  MOAI22D1BWP30P140 U174 ( .A1(n128), .A2(n118), .B1(n126), .B2(i_data_bus[12]), .ZN(N299) );
  INVD1BWP30P140 U175 ( .I(i_data_bus[55]), .ZN(n119) );
  MOAI22D1BWP30P140 U176 ( .A1(n128), .A2(n119), .B1(n126), .B2(i_data_bus[23]), .ZN(N310) );
  INVD1BWP30P140 U177 ( .I(i_data_bus[43]), .ZN(n120) );
  MOAI22D1BWP30P140 U178 ( .A1(n128), .A2(n120), .B1(n126), .B2(i_data_bus[11]), .ZN(N298) );
  INVD1BWP30P140 U179 ( .I(i_data_bus[54]), .ZN(n121) );
  MOAI22D1BWP30P140 U180 ( .A1(n128), .A2(n121), .B1(n126), .B2(i_data_bus[22]), .ZN(N309) );
  INVD1BWP30P140 U181 ( .I(i_data_bus[42]), .ZN(n122) );
  MOAI22D1BWP30P140 U182 ( .A1(n128), .A2(n122), .B1(n126), .B2(i_data_bus[10]), .ZN(N297) );
  INVD1BWP30P140 U183 ( .I(i_data_bus[53]), .ZN(n123) );
  MOAI22D1BWP30P140 U184 ( .A1(n128), .A2(n123), .B1(n126), .B2(i_data_bus[21]), .ZN(N308) );
  INVD1BWP30P140 U185 ( .I(i_data_bus[41]), .ZN(n124) );
  MOAI22D1BWP30P140 U186 ( .A1(n128), .A2(n124), .B1(n126), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140 U187 ( .I(i_data_bus[52]), .ZN(n125) );
  MOAI22D1BWP30P140 U188 ( .A1(n128), .A2(n125), .B1(n126), .B2(i_data_bus[20]), .ZN(N307) );
  INVD1BWP30P140 U189 ( .I(i_data_bus[40]), .ZN(n127) );
  MOAI22D1BWP30P140 U190 ( .A1(n128), .A2(n127), .B1(n9), .B2(i_data_bus[8]), 
        .ZN(N295) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_53 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  INVD3BWP30P140 U3 ( .I(n17), .ZN(n104) );
  NR2D4BWP30P140 U4 ( .A1(n13), .A2(n12), .ZN(n17) );
  NR2D1BWP30P140 U5 ( .A1(i_cmd[1]), .A2(n91), .ZN(n24) );
  ND2OPTIBD1BWP30P140 U6 ( .A1(i_valid[0]), .A2(n11), .ZN(n1) );
  INVD6BWP30P140 U7 ( .I(n36), .ZN(n2) );
  ND2OPTPAD1BWP30P140 U8 ( .A1(i_cmd[0]), .A2(n11), .ZN(n12) );
  MUX2NOPTD2BWP30P140 U9 ( .I0(i_valid[0]), .I1(i_valid[1]), .S(i_cmd[1]), 
        .ZN(n13) );
  MUX2NOPTD2BWP30P140 U10 ( .I0(i_valid[0]), .I1(i_valid[1]), .S(i_cmd[0]), 
        .ZN(n23) );
  OR2D8BWP30P140 U11 ( .A1(n14), .A2(i_cmd[0]), .Z(n106) );
  CKND2D4BWP30P140 U12 ( .A1(i_valid[0]), .A2(n11), .ZN(n14) );
  INVD2BWP30P140 U13 ( .I(n106), .ZN(n9) );
  INVD8BWP30P140 U14 ( .I(n106), .ZN(n125) );
  INVD1BWP30P140 U15 ( .I(i_cmd[0]), .ZN(n94) );
  ND3OPTPAD2BWP30P140 U16 ( .A1(i_cmd[1]), .A2(i_valid[1]), .A3(n11), .ZN(n96)
         );
  ND2D1BWP30P140 U17 ( .A1(n10), .A2(i_en), .ZN(n91) );
  ND2D1BWP30P140 U18 ( .A1(n106), .A2(n95), .ZN(N353) );
  IND2D1BWP30P140 U19 ( .A1(n94), .B1(n93), .ZN(n95) );
  NR2D1BWP30P140 U20 ( .A1(n92), .A2(n91), .ZN(n93) );
  INVD1BWP30P140 U21 ( .I(i_valid[1]), .ZN(n92) );
  OAI21D1BWP30P140 U22 ( .A1(n104), .A2(n90), .B(n89), .ZN(N287) );
  OAI21D1BWP30P140 U23 ( .A1(n104), .A2(n88), .B(n87), .ZN(N288) );
  ND2D1BWP30P140 U24 ( .A1(n9), .A2(i_data_bus[1]), .ZN(n87) );
  ND2D1BWP30P140 U25 ( .A1(n84), .A2(i_data_bus[47]), .ZN(n50) );
  ND2D1BWP30P140 U26 ( .A1(n84), .A2(i_data_bus[51]), .ZN(n58) );
  ND2D1BWP30P140 U27 ( .A1(n84), .A2(i_data_bus[52]), .ZN(n60) );
  ND2D1BWP30P140 U28 ( .A1(n84), .A2(i_data_bus[53]), .ZN(n62) );
  ND2D1BWP30P140 U29 ( .A1(n84), .A2(i_data_bus[54]), .ZN(n64) );
  ND2D1BWP30P140 U30 ( .A1(n84), .A2(i_data_bus[55]), .ZN(n66) );
  ND2D1BWP30P140 U31 ( .A1(n84), .A2(i_data_bus[56]), .ZN(n85) );
  ND2D1BWP30P140 U32 ( .A1(n84), .A2(i_data_bus[57]), .ZN(n82) );
  ND2D1BWP30P140 U33 ( .A1(n84), .A2(i_data_bus[58]), .ZN(n80) );
  ND2D1BWP30P140 U34 ( .A1(n84), .A2(i_data_bus[59]), .ZN(n78) );
  ND2D1BWP30P140 U35 ( .A1(n84), .A2(i_data_bus[60]), .ZN(n76) );
  ND2D1BWP30P140 U36 ( .A1(n84), .A2(i_data_bus[61]), .ZN(n74) );
  ND2D1BWP30P140 U37 ( .A1(n84), .A2(i_data_bus[62]), .ZN(n72) );
  ND2D1BWP30P140 U38 ( .A1(n84), .A2(i_data_bus[63]), .ZN(n68) );
  OAI22D1BWP30P140 U39 ( .A1(n127), .A2(n22), .B1(n106), .B2(n69), .ZN(N318)
         );
  OAI22D1BWP30P140 U40 ( .A1(n127), .A2(n21), .B1(n106), .B2(n59), .ZN(N306)
         );
  OAI22D1BWP30P140 U41 ( .A1(n127), .A2(n20), .B1(n106), .B2(n57), .ZN(N305)
         );
  OAI22D1BWP30P140 U42 ( .A1(n127), .A2(n19), .B1(n106), .B2(n73), .ZN(N317)
         );
  OAI22D1BWP30P140 U43 ( .A1(n106), .A2(n30), .B1(n104), .B2(n18), .ZN(N291)
         );
  INR2D4BWP30P140 U44 ( .A1(n24), .B1(n23), .ZN(n36) );
  INVD1BWP30P140 U45 ( .I(n91), .ZN(n11) );
  INVD1BWP30P140 U46 ( .I(rst), .ZN(n10) );
  INVD6BWP30P140 U47 ( .I(n17), .ZN(n127) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[61]), .ZN(n15) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[29]), .ZN(n75) );
  OAI22D1BWP30P140 U50 ( .A1(n127), .A2(n15), .B1(n106), .B2(n75), .ZN(N316)
         );
  INVD1BWP30P140 U51 ( .I(i_data_bus[49]), .ZN(n16) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[17]), .ZN(n55) );
  OAI22D1BWP30P140 U53 ( .A1(n127), .A2(n16), .B1(n106), .B2(n55), .ZN(N304)
         );
  INVD1BWP30P140 U54 ( .I(i_data_bus[4]), .ZN(n30) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[36]), .ZN(n18) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[62]), .ZN(n19) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[30]), .ZN(n73) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[50]), .ZN(n20) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[18]), .ZN(n57) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[51]), .ZN(n21) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[19]), .ZN(n59) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[63]), .ZN(n22) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[31]), .ZN(n69) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[1]), .ZN(n26) );
  INVD6BWP30P140 U65 ( .I(n96), .ZN(n84) );
  ND2OPTIBD1BWP30P140 U66 ( .A1(n84), .A2(i_data_bus[33]), .ZN(n25) );
  OAI21D1BWP30P140 U67 ( .A1(n2), .A2(n26), .B(n25), .ZN(N320) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[2]), .ZN(n28) );
  ND2OPTIBD1BWP30P140 U69 ( .A1(n84), .A2(i_data_bus[34]), .ZN(n27) );
  OAI21D1BWP30P140 U70 ( .A1(n2), .A2(n28), .B(n27), .ZN(N321) );
  ND2OPTIBD1BWP30P140 U71 ( .A1(n84), .A2(i_data_bus[36]), .ZN(n29) );
  OAI21D1BWP30P140 U72 ( .A1(n2), .A2(n30), .B(n29), .ZN(N323) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[5]), .ZN(n98) );
  ND2OPTIBD1BWP30P140 U74 ( .A1(n84), .A2(i_data_bus[37]), .ZN(n31) );
  OAI21D1BWP30P140 U75 ( .A1(n2), .A2(n98), .B(n31), .ZN(N324) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[6]), .ZN(n100) );
  ND2OPTIBD1BWP30P140 U77 ( .A1(n84), .A2(i_data_bus[38]), .ZN(n32) );
  OAI21D1BWP30P140 U78 ( .A1(n2), .A2(n100), .B(n32), .ZN(N325) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[7]), .ZN(n102) );
  ND2OPTIBD1BWP30P140 U80 ( .A1(n84), .A2(i_data_bus[39]), .ZN(n33) );
  OAI21D1BWP30P140 U81 ( .A1(n2), .A2(n102), .B(n33), .ZN(N326) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[8]), .ZN(n35) );
  ND2OPTIBD1BWP30P140 U83 ( .A1(n84), .A2(i_data_bus[40]), .ZN(n34) );
  OAI21D1BWP30P140 U84 ( .A1(n2), .A2(n35), .B(n34), .ZN(N327) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[9]), .ZN(n38) );
  ND2OPTIBD1BWP30P140 U86 ( .A1(n84), .A2(i_data_bus[41]), .ZN(n37) );
  OAI21D1BWP30P140 U87 ( .A1(n2), .A2(n38), .B(n37), .ZN(N328) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[10]), .ZN(n40) );
  ND2OPTIBD1BWP30P140 U89 ( .A1(n84), .A2(i_data_bus[42]), .ZN(n39) );
  OAI21D1BWP30P140 U90 ( .A1(n2), .A2(n40), .B(n39), .ZN(N329) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[11]), .ZN(n42) );
  ND2OPTIBD1BWP30P140 U92 ( .A1(n84), .A2(i_data_bus[43]), .ZN(n41) );
  OAI21D1BWP30P140 U93 ( .A1(n2), .A2(n42), .B(n41), .ZN(N330) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[12]), .ZN(n44) );
  ND2OPTIBD1BWP30P140 U95 ( .A1(n84), .A2(i_data_bus[44]), .ZN(n43) );
  OAI21D1BWP30P140 U96 ( .A1(n2), .A2(n44), .B(n43), .ZN(N331) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[3]), .ZN(n105) );
  ND2OPTIBD1BWP30P140 U98 ( .A1(n84), .A2(i_data_bus[35]), .ZN(n45) );
  OAI21D1BWP30P140 U99 ( .A1(n2), .A2(n105), .B(n45), .ZN(N322) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[13]), .ZN(n47) );
  ND2OPTIBD1BWP30P140 U101 ( .A1(n84), .A2(i_data_bus[45]), .ZN(n46) );
  OAI21D1BWP30P140 U102 ( .A1(n2), .A2(n47), .B(n46), .ZN(N332) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[14]), .ZN(n49) );
  ND2OPTIBD1BWP30P140 U104 ( .A1(n84), .A2(i_data_bus[46]), .ZN(n48) );
  OAI21D1BWP30P140 U105 ( .A1(n2), .A2(n49), .B(n48), .ZN(N333) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[15]), .ZN(n51) );
  OAI21D1BWP30P140 U107 ( .A1(n2), .A2(n51), .B(n50), .ZN(N334) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[16]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U109 ( .A1(n84), .A2(i_data_bus[48]), .ZN(n52) );
  OAI21D1BWP30P140 U110 ( .A1(n2), .A2(n53), .B(n52), .ZN(N335) );
  ND2OPTIBD1BWP30P140 U111 ( .A1(n84), .A2(i_data_bus[49]), .ZN(n54) );
  OAI21D1BWP30P140 U112 ( .A1(n2), .A2(n55), .B(n54), .ZN(N336) );
  ND2OPTIBD1BWP30P140 U113 ( .A1(n84), .A2(i_data_bus[50]), .ZN(n56) );
  OAI21D1BWP30P140 U114 ( .A1(n2), .A2(n57), .B(n56), .ZN(N337) );
  OAI21D1BWP30P140 U115 ( .A1(n2), .A2(n59), .B(n58), .ZN(N338) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[20]), .ZN(n61) );
  OAI21D1BWP30P140 U117 ( .A1(n2), .A2(n61), .B(n60), .ZN(N339) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[21]), .ZN(n63) );
  OAI21D1BWP30P140 U119 ( .A1(n2), .A2(n63), .B(n62), .ZN(N340) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[22]), .ZN(n65) );
  OAI21D1BWP30P140 U121 ( .A1(n2), .A2(n65), .B(n64), .ZN(N341) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[23]), .ZN(n67) );
  OAI21D1BWP30P140 U123 ( .A1(n2), .A2(n67), .B(n66), .ZN(N342) );
  OAI21D1BWP30P140 U124 ( .A1(n2), .A2(n69), .B(n68), .ZN(N350) );
  INVD1BWP30P140 U125 ( .I(i_data_bus[0]), .ZN(n71) );
  ND2OPTIBD1BWP30P140 U126 ( .A1(n84), .A2(i_data_bus[32]), .ZN(n70) );
  OAI21D1BWP30P140 U127 ( .A1(n2), .A2(n71), .B(n70), .ZN(N319) );
  OAI21D1BWP30P140 U128 ( .A1(n2), .A2(n73), .B(n72), .ZN(N349) );
  OAI21D1BWP30P140 U129 ( .A1(n2), .A2(n75), .B(n74), .ZN(N348) );
  INVD1BWP30P140 U130 ( .I(i_data_bus[28]), .ZN(n77) );
  OAI21D1BWP30P140 U131 ( .A1(n2), .A2(n77), .B(n76), .ZN(N347) );
  INVD1BWP30P140 U132 ( .I(i_data_bus[27]), .ZN(n79) );
  OAI21D1BWP30P140 U133 ( .A1(n2), .A2(n79), .B(n78), .ZN(N346) );
  INVD1BWP30P140 U134 ( .I(i_data_bus[26]), .ZN(n81) );
  OAI21D1BWP30P140 U135 ( .A1(n2), .A2(n81), .B(n80), .ZN(N345) );
  INVD1BWP30P140 U136 ( .I(i_data_bus[25]), .ZN(n83) );
  OAI21D1BWP30P140 U137 ( .A1(n2), .A2(n83), .B(n82), .ZN(N344) );
  INVD1BWP30P140 U138 ( .I(i_data_bus[24]), .ZN(n86) );
  OAI21D1BWP30P140 U139 ( .A1(n2), .A2(n86), .B(n85), .ZN(N343) );
  INVD1BWP30P140 U140 ( .I(i_data_bus[33]), .ZN(n88) );
  INVD1BWP30P140 U141 ( .I(i_data_bus[32]), .ZN(n90) );
  IND2D2BWP30P140 U142 ( .A1(n106), .B1(i_data_bus[0]), .ZN(n89) );
  OAI21D1BWP30P140 U143 ( .A1(n1), .A2(i_cmd[1]), .B(n96), .ZN(N354) );
  INVD1BWP30P140 U144 ( .I(i_data_bus[37]), .ZN(n97) );
  OAI22D1BWP30P140 U145 ( .A1(n106), .A2(n98), .B1(n104), .B2(n97), .ZN(N292)
         );
  INVD1BWP30P140 U146 ( .I(i_data_bus[38]), .ZN(n99) );
  OAI22D1BWP30P140 U147 ( .A1(n106), .A2(n100), .B1(n104), .B2(n99), .ZN(N293)
         );
  INVD1BWP30P140 U148 ( .I(i_data_bus[39]), .ZN(n101) );
  OAI22D1BWP30P140 U149 ( .A1(n106), .A2(n102), .B1(n104), .B2(n101), .ZN(N294) );
  INVD1BWP30P140 U150 ( .I(i_data_bus[35]), .ZN(n103) );
  OAI22D1BWP30P140 U151 ( .A1(n106), .A2(n105), .B1(n104), .B2(n103), .ZN(N290) );
  INVD1BWP30P140 U152 ( .I(i_data_bus[60]), .ZN(n107) );
  MOAI22D1BWP30P140 U153 ( .A1(n127), .A2(n107), .B1(n125), .B2(i_data_bus[28]), .ZN(N315) );
  INVD1BWP30P140 U154 ( .I(i_data_bus[48]), .ZN(n108) );
  MOAI22D1BWP30P140 U155 ( .A1(n127), .A2(n108), .B1(n125), .B2(i_data_bus[16]), .ZN(N303) );
  INVD1BWP30P140 U156 ( .I(i_data_bus[34]), .ZN(n109) );
  MOAI22D1BWP30P140 U157 ( .A1(n127), .A2(n109), .B1(n125), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140 U158 ( .I(i_data_bus[59]), .ZN(n110) );
  MOAI22D1BWP30P140 U159 ( .A1(n127), .A2(n110), .B1(n125), .B2(i_data_bus[27]), .ZN(N314) );
  INVD1BWP30P140 U160 ( .I(i_data_bus[47]), .ZN(n111) );
  MOAI22D1BWP30P140 U161 ( .A1(n127), .A2(n111), .B1(n125), .B2(i_data_bus[15]), .ZN(N302) );
  INVD1BWP30P140 U162 ( .I(i_data_bus[58]), .ZN(n112) );
  MOAI22D1BWP30P140 U163 ( .A1(n127), .A2(n112), .B1(n125), .B2(i_data_bus[26]), .ZN(N313) );
  INVD1BWP30P140 U164 ( .I(i_data_bus[46]), .ZN(n113) );
  MOAI22D1BWP30P140 U165 ( .A1(n127), .A2(n113), .B1(n125), .B2(i_data_bus[14]), .ZN(N301) );
  INVD1BWP30P140 U166 ( .I(i_data_bus[57]), .ZN(n114) );
  MOAI22D1BWP30P140 U167 ( .A1(n127), .A2(n114), .B1(n125), .B2(i_data_bus[25]), .ZN(N312) );
  INVD1BWP30P140 U168 ( .I(i_data_bus[45]), .ZN(n115) );
  MOAI22D1BWP30P140 U169 ( .A1(n127), .A2(n115), .B1(n125), .B2(i_data_bus[13]), .ZN(N300) );
  INVD1BWP30P140 U170 ( .I(i_data_bus[56]), .ZN(n116) );
  MOAI22D1BWP30P140 U171 ( .A1(n127), .A2(n116), .B1(n125), .B2(i_data_bus[24]), .ZN(N311) );
  INVD1BWP30P140 U172 ( .I(i_data_bus[44]), .ZN(n117) );
  MOAI22D1BWP30P140 U173 ( .A1(n127), .A2(n117), .B1(n125), .B2(i_data_bus[12]), .ZN(N299) );
  INVD1BWP30P140 U174 ( .I(i_data_bus[55]), .ZN(n118) );
  MOAI22D1BWP30P140 U175 ( .A1(n127), .A2(n118), .B1(n125), .B2(i_data_bus[23]), .ZN(N310) );
  INVD1BWP30P140 U176 ( .I(i_data_bus[43]), .ZN(n119) );
  MOAI22D1BWP30P140 U177 ( .A1(n127), .A2(n119), .B1(n125), .B2(i_data_bus[11]), .ZN(N298) );
  INVD1BWP30P140 U178 ( .I(i_data_bus[54]), .ZN(n120) );
  MOAI22D1BWP30P140 U179 ( .A1(n127), .A2(n120), .B1(n125), .B2(i_data_bus[22]), .ZN(N309) );
  INVD1BWP30P140 U180 ( .I(i_data_bus[42]), .ZN(n121) );
  MOAI22D1BWP30P140 U181 ( .A1(n127), .A2(n121), .B1(n125), .B2(i_data_bus[10]), .ZN(N297) );
  INVD1BWP30P140 U182 ( .I(i_data_bus[53]), .ZN(n122) );
  MOAI22D1BWP30P140 U183 ( .A1(n127), .A2(n122), .B1(n125), .B2(i_data_bus[21]), .ZN(N308) );
  INVD1BWP30P140 U184 ( .I(i_data_bus[41]), .ZN(n123) );
  MOAI22D1BWP30P140 U185 ( .A1(n127), .A2(n123), .B1(n125), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140 U186 ( .I(i_data_bus[52]), .ZN(n124) );
  MOAI22D1BWP30P140 U187 ( .A1(n127), .A2(n124), .B1(n125), .B2(i_data_bus[20]), .ZN(N307) );
  INVD1BWP30P140 U188 ( .I(i_data_bus[40]), .ZN(n126) );
  MOAI22D1BWP30P140 U189 ( .A1(n127), .A2(n126), .B1(n9), .B2(i_data_bus[8]), 
        .ZN(N295) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_54 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n8, n9, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(o_data_bus[2]) );
  DFD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(o_data_bus[8]) );
  DFD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(o_data_bus[9]) );
  DFD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  INVD3BWP30P140 U3 ( .I(n29), .ZN(n117) );
  NR2D4BWP30P140 U4 ( .A1(n25), .A2(n24), .ZN(n29) );
  NR2D1BWP30P140 U5 ( .A1(i_cmd[1]), .A2(n103), .ZN(n36) );
  INVD6BWP30P140 U6 ( .I(n59), .ZN(n1) );
  ND2OPTPAD1BWP30P140 U7 ( .A1(i_cmd[0]), .A2(n23), .ZN(n24) );
  AN2D1BWP30P140 U8 ( .A1(i_valid[0]), .A2(n23), .Z(n8) );
  MUX2NOPTD2BWP30P140 U9 ( .I0(i_valid[0]), .I1(i_valid[1]), .S(i_cmd[1]), 
        .ZN(n25) );
  MUX2NOPTD2BWP30P140 U10 ( .I0(i_valid[0]), .I1(i_valid[1]), .S(i_cmd[0]), 
        .ZN(n35) );
  OR2D8BWP30P140 U11 ( .A1(n26), .A2(i_cmd[0]), .Z(n119) );
  CKND2D4BWP30P140 U12 ( .A1(i_valid[0]), .A2(n23), .ZN(n26) );
  INVD2BWP30P140 U13 ( .I(n119), .ZN(n9) );
  INVD8BWP30P140 U14 ( .I(n119), .ZN(n138) );
  INVD1BWP30P140 U15 ( .I(i_cmd[0]), .ZN(n106) );
  ND3OPTPAD2BWP30P140 U16 ( .A1(i_cmd[1]), .A2(i_valid[1]), .A3(n23), .ZN(n108) );
  ND2D1BWP30P140 U17 ( .A1(n22), .A2(i_en), .ZN(n103) );
  ND2D1BWP30P140 U18 ( .A1(n119), .A2(n107), .ZN(N353) );
  IND2D1BWP30P140 U19 ( .A1(n106), .B1(n105), .ZN(n107) );
  NR2D1BWP30P140 U20 ( .A1(n104), .A2(n103), .ZN(n105) );
  INVD1BWP30P140 U21 ( .I(i_valid[1]), .ZN(n104) );
  OAI21D1BWP30P140 U22 ( .A1(n117), .A2(n102), .B(n101), .ZN(N287) );
  OAI21D1BWP30P140 U23 ( .A1(n117), .A2(n100), .B(n99), .ZN(N288) );
  ND2D1BWP30P140 U24 ( .A1(n9), .A2(i_data_bus[1]), .ZN(n99) );
  ND2D1BWP30P140 U25 ( .A1(n96), .A2(i_data_bus[50]), .ZN(n62) );
  ND2D1BWP30P140 U26 ( .A1(n96), .A2(i_data_bus[51]), .ZN(n60) );
  ND2D1BWP30P140 U27 ( .A1(n96), .A2(i_data_bus[52]), .ZN(n57) );
  ND2D1BWP30P140 U28 ( .A1(n96), .A2(i_data_bus[53]), .ZN(n55) );
  ND2D1BWP30P140 U29 ( .A1(n96), .A2(i_data_bus[54]), .ZN(n53) );
  ND2D1BWP30P140 U30 ( .A1(n96), .A2(i_data_bus[55]), .ZN(n51) );
  ND2D1BWP30P140 U31 ( .A1(n96), .A2(i_data_bus[56]), .ZN(n49) );
  ND2D1BWP30P140 U32 ( .A1(n96), .A2(i_data_bus[57]), .ZN(n47) );
  ND2D1BWP30P140 U33 ( .A1(n96), .A2(i_data_bus[58]), .ZN(n45) );
  ND2D1BWP30P140 U34 ( .A1(n96), .A2(i_data_bus[59]), .ZN(n43) );
  ND2D1BWP30P140 U35 ( .A1(n96), .A2(i_data_bus[60]), .ZN(n97) );
  ND2D1BWP30P140 U36 ( .A1(n96), .A2(i_data_bus[61]), .ZN(n41) );
  ND2D1BWP30P140 U37 ( .A1(n96), .A2(i_data_bus[62]), .ZN(n39) );
  ND2D1BWP30P140 U38 ( .A1(n96), .A2(i_data_bus[63]), .ZN(n37) );
  OAI22D1BWP30P140 U39 ( .A1(n140), .A2(n34), .B1(n119), .B2(n65), .ZN(N304)
         );
  OAI22D1BWP30P140 U40 ( .A1(n140), .A2(n33), .B1(n119), .B2(n38), .ZN(N318)
         );
  OAI22D1BWP30P140 U41 ( .A1(n140), .A2(n32), .B1(n119), .B2(n63), .ZN(N305)
         );
  OAI22D1BWP30P140 U42 ( .A1(n140), .A2(n31), .B1(n119), .B2(n40), .ZN(N317)
         );
  OAI22D1BWP30P140 U43 ( .A1(n119), .A2(n86), .B1(n117), .B2(n30), .ZN(N293)
         );
  INR2D4BWP30P140 U44 ( .A1(n36), .B1(n35), .ZN(n59) );
  INVD1BWP30P140 U45 ( .I(n103), .ZN(n23) );
  INVD1BWP30P140 U46 ( .I(rst), .ZN(n22) );
  INVD6BWP30P140 U47 ( .I(n29), .ZN(n140) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[61]), .ZN(n27) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[29]), .ZN(n42) );
  OAI22D1BWP30P140 U50 ( .A1(n140), .A2(n27), .B1(n119), .B2(n42), .ZN(N316)
         );
  INVD1BWP30P140 U51 ( .I(i_data_bus[51]), .ZN(n28) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[19]), .ZN(n61) );
  OAI22D1BWP30P140 U53 ( .A1(n140), .A2(n28), .B1(n119), .B2(n61), .ZN(N306)
         );
  INVD1BWP30P140 U54 ( .I(i_data_bus[6]), .ZN(n86) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[38]), .ZN(n30) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[62]), .ZN(n31) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[30]), .ZN(n40) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[50]), .ZN(n32) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[18]), .ZN(n63) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[63]), .ZN(n33) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[31]), .ZN(n38) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[49]), .ZN(n34) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[17]), .ZN(n65) );
  INVD6BWP30P140 U64 ( .I(n108), .ZN(n96) );
  OAI21D1BWP30P140 U65 ( .A1(n1), .A2(n38), .B(n37), .ZN(N350) );
  OAI21D1BWP30P140 U66 ( .A1(n1), .A2(n40), .B(n39), .ZN(N349) );
  OAI21D1BWP30P140 U67 ( .A1(n1), .A2(n42), .B(n41), .ZN(N348) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[27]), .ZN(n44) );
  OAI21D1BWP30P140 U69 ( .A1(n1), .A2(n44), .B(n43), .ZN(N346) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[26]), .ZN(n46) );
  OAI21D1BWP30P140 U71 ( .A1(n1), .A2(n46), .B(n45), .ZN(N345) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[25]), .ZN(n48) );
  OAI21D1BWP30P140 U73 ( .A1(n1), .A2(n48), .B(n47), .ZN(N344) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[24]), .ZN(n50) );
  OAI21D1BWP30P140 U75 ( .A1(n1), .A2(n50), .B(n49), .ZN(N343) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[23]), .ZN(n52) );
  OAI21D1BWP30P140 U77 ( .A1(n1), .A2(n52), .B(n51), .ZN(N342) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n54) );
  OAI21D1BWP30P140 U79 ( .A1(n1), .A2(n54), .B(n53), .ZN(N341) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[21]), .ZN(n56) );
  OAI21D1BWP30P140 U81 ( .A1(n1), .A2(n56), .B(n55), .ZN(N340) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[20]), .ZN(n58) );
  OAI21D1BWP30P140 U83 ( .A1(n1), .A2(n58), .B(n57), .ZN(N339) );
  OAI21D1BWP30P140 U84 ( .A1(n1), .A2(n61), .B(n60), .ZN(N338) );
  OAI21D1BWP30P140 U85 ( .A1(n1), .A2(n63), .B(n62), .ZN(N337) );
  ND2OPTIBD1BWP30P140 U86 ( .A1(n96), .A2(i_data_bus[49]), .ZN(n64) );
  OAI21D1BWP30P140 U87 ( .A1(n1), .A2(n65), .B(n64), .ZN(N336) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[16]), .ZN(n67) );
  ND2OPTIBD1BWP30P140 U89 ( .A1(n96), .A2(i_data_bus[48]), .ZN(n66) );
  OAI21D1BWP30P140 U90 ( .A1(n1), .A2(n67), .B(n66), .ZN(N335) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[15]), .ZN(n69) );
  ND2OPTIBD1BWP30P140 U92 ( .A1(n96), .A2(i_data_bus[47]), .ZN(n68) );
  OAI21D1BWP30P140 U93 ( .A1(n1), .A2(n69), .B(n68), .ZN(N334) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[14]), .ZN(n71) );
  ND2OPTIBD1BWP30P140 U95 ( .A1(n96), .A2(i_data_bus[46]), .ZN(n70) );
  OAI21D1BWP30P140 U96 ( .A1(n1), .A2(n71), .B(n70), .ZN(N333) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[13]), .ZN(n73) );
  ND2OPTIBD1BWP30P140 U98 ( .A1(n96), .A2(i_data_bus[45]), .ZN(n72) );
  OAI21D1BWP30P140 U99 ( .A1(n1), .A2(n73), .B(n72), .ZN(N332) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[12]), .ZN(n75) );
  ND2OPTIBD1BWP30P140 U101 ( .A1(n96), .A2(i_data_bus[44]), .ZN(n74) );
  OAI21D1BWP30P140 U102 ( .A1(n1), .A2(n75), .B(n74), .ZN(N331) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[11]), .ZN(n77) );
  ND2OPTIBD1BWP30P140 U104 ( .A1(n96), .A2(i_data_bus[43]), .ZN(n76) );
  OAI21D1BWP30P140 U105 ( .A1(n1), .A2(n77), .B(n76), .ZN(N330) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[10]), .ZN(n79) );
  ND2OPTIBD1BWP30P140 U107 ( .A1(n96), .A2(i_data_bus[42]), .ZN(n78) );
  OAI21D1BWP30P140 U108 ( .A1(n1), .A2(n79), .B(n78), .ZN(N329) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[9]), .ZN(n81) );
  ND2OPTIBD1BWP30P140 U110 ( .A1(n96), .A2(i_data_bus[41]), .ZN(n80) );
  OAI21D1BWP30P140 U111 ( .A1(n1), .A2(n81), .B(n80), .ZN(N328) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[8]), .ZN(n83) );
  ND2OPTIBD1BWP30P140 U113 ( .A1(n96), .A2(i_data_bus[40]), .ZN(n82) );
  OAI21D1BWP30P140 U114 ( .A1(n1), .A2(n83), .B(n82), .ZN(N327) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[7]), .ZN(n111) );
  ND2OPTIBD1BWP30P140 U116 ( .A1(n96), .A2(i_data_bus[39]), .ZN(n84) );
  OAI21D1BWP30P140 U117 ( .A1(n1), .A2(n111), .B(n84), .ZN(N326) );
  ND2OPTIBD1BWP30P140 U118 ( .A1(n96), .A2(i_data_bus[38]), .ZN(n85) );
  OAI21D1BWP30P140 U119 ( .A1(n1), .A2(n86), .B(n85), .ZN(N325) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[5]), .ZN(n118) );
  ND2OPTIBD1BWP30P140 U121 ( .A1(n96), .A2(i_data_bus[37]), .ZN(n87) );
  OAI21D1BWP30P140 U122 ( .A1(n1), .A2(n118), .B(n87), .ZN(N324) );
  INVD1BWP30P140 U123 ( .I(i_data_bus[4]), .ZN(n115) );
  ND2OPTIBD1BWP30P140 U124 ( .A1(n96), .A2(i_data_bus[36]), .ZN(n88) );
  OAI21D1BWP30P140 U125 ( .A1(n1), .A2(n115), .B(n88), .ZN(N323) );
  INVD1BWP30P140 U126 ( .I(i_data_bus[3]), .ZN(n113) );
  ND2OPTIBD1BWP30P140 U127 ( .A1(n96), .A2(i_data_bus[35]), .ZN(n89) );
  OAI21D1BWP30P140 U128 ( .A1(n1), .A2(n113), .B(n89), .ZN(N322) );
  INVD1BWP30P140 U129 ( .I(i_data_bus[2]), .ZN(n91) );
  ND2OPTIBD1BWP30P140 U130 ( .A1(n96), .A2(i_data_bus[34]), .ZN(n90) );
  OAI21D1BWP30P140 U131 ( .A1(n1), .A2(n91), .B(n90), .ZN(N321) );
  INVD1BWP30P140 U132 ( .I(i_data_bus[1]), .ZN(n93) );
  ND2OPTIBD1BWP30P140 U133 ( .A1(n96), .A2(i_data_bus[33]), .ZN(n92) );
  OAI21D1BWP30P140 U134 ( .A1(n1), .A2(n93), .B(n92), .ZN(N320) );
  INVD1BWP30P140 U135 ( .I(i_data_bus[0]), .ZN(n95) );
  ND2OPTIBD1BWP30P140 U136 ( .A1(n96), .A2(i_data_bus[32]), .ZN(n94) );
  OAI21D1BWP30P140 U137 ( .A1(n1), .A2(n95), .B(n94), .ZN(N319) );
  INVD1BWP30P140 U138 ( .I(i_data_bus[28]), .ZN(n98) );
  OAI21D1BWP30P140 U139 ( .A1(n1), .A2(n98), .B(n97), .ZN(N347) );
  INVD1BWP30P140 U140 ( .I(i_data_bus[33]), .ZN(n100) );
  INVD1BWP30P140 U141 ( .I(i_data_bus[32]), .ZN(n102) );
  IND2D2BWP30P140 U142 ( .A1(n119), .B1(i_data_bus[0]), .ZN(n101) );
  INVD1BWP30P140 U143 ( .I(n8), .ZN(n109) );
  OAI21D1BWP30P140 U144 ( .A1(n109), .A2(i_cmd[1]), .B(n108), .ZN(N354) );
  INVD1BWP30P140 U145 ( .I(i_data_bus[39]), .ZN(n110) );
  OAI22D1BWP30P140 U146 ( .A1(n119), .A2(n111), .B1(n117), .B2(n110), .ZN(N294) );
  INVD1BWP30P140 U147 ( .I(i_data_bus[35]), .ZN(n112) );
  OAI22D1BWP30P140 U148 ( .A1(n119), .A2(n113), .B1(n117), .B2(n112), .ZN(N290) );
  INVD1BWP30P140 U149 ( .I(i_data_bus[36]), .ZN(n114) );
  OAI22D1BWP30P140 U150 ( .A1(n119), .A2(n115), .B1(n117), .B2(n114), .ZN(N291) );
  INVD1BWP30P140 U151 ( .I(i_data_bus[37]), .ZN(n116) );
  OAI22D1BWP30P140 U152 ( .A1(n119), .A2(n118), .B1(n117), .B2(n116), .ZN(N292) );
  INVD1BWP30P140 U153 ( .I(i_data_bus[60]), .ZN(n120) );
  MOAI22D1BWP30P140 U154 ( .A1(n140), .A2(n120), .B1(n138), .B2(i_data_bus[28]), .ZN(N315) );
  INVD1BWP30P140 U155 ( .I(i_data_bus[48]), .ZN(n121) );
  MOAI22D1BWP30P140 U156 ( .A1(n140), .A2(n121), .B1(n138), .B2(i_data_bus[16]), .ZN(N303) );
  INVD1BWP30P140 U157 ( .I(i_data_bus[34]), .ZN(n122) );
  MOAI22D1BWP30P140 U158 ( .A1(n140), .A2(n122), .B1(n138), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140 U159 ( .I(i_data_bus[59]), .ZN(n123) );
  MOAI22D1BWP30P140 U160 ( .A1(n140), .A2(n123), .B1(n138), .B2(i_data_bus[27]), .ZN(N314) );
  INVD1BWP30P140 U161 ( .I(i_data_bus[47]), .ZN(n124) );
  MOAI22D1BWP30P140 U162 ( .A1(n140), .A2(n124), .B1(n138), .B2(i_data_bus[15]), .ZN(N302) );
  INVD1BWP30P140 U163 ( .I(i_data_bus[58]), .ZN(n125) );
  MOAI22D1BWP30P140 U164 ( .A1(n140), .A2(n125), .B1(n138), .B2(i_data_bus[26]), .ZN(N313) );
  INVD1BWP30P140 U165 ( .I(i_data_bus[46]), .ZN(n126) );
  MOAI22D1BWP30P140 U166 ( .A1(n140), .A2(n126), .B1(n138), .B2(i_data_bus[14]), .ZN(N301) );
  INVD1BWP30P140 U167 ( .I(i_data_bus[57]), .ZN(n127) );
  MOAI22D1BWP30P140 U168 ( .A1(n140), .A2(n127), .B1(n138), .B2(i_data_bus[25]), .ZN(N312) );
  INVD1BWP30P140 U169 ( .I(i_data_bus[45]), .ZN(n128) );
  MOAI22D1BWP30P140 U170 ( .A1(n140), .A2(n128), .B1(n138), .B2(i_data_bus[13]), .ZN(N300) );
  INVD1BWP30P140 U171 ( .I(i_data_bus[56]), .ZN(n129) );
  MOAI22D1BWP30P140 U172 ( .A1(n140), .A2(n129), .B1(n138), .B2(i_data_bus[24]), .ZN(N311) );
  INVD1BWP30P140 U173 ( .I(i_data_bus[44]), .ZN(n130) );
  MOAI22D1BWP30P140 U174 ( .A1(n140), .A2(n130), .B1(n138), .B2(i_data_bus[12]), .ZN(N299) );
  INVD1BWP30P140 U175 ( .I(i_data_bus[55]), .ZN(n131) );
  MOAI22D1BWP30P140 U176 ( .A1(n140), .A2(n131), .B1(n138), .B2(i_data_bus[23]), .ZN(N310) );
  INVD1BWP30P140 U177 ( .I(i_data_bus[43]), .ZN(n132) );
  MOAI22D1BWP30P140 U178 ( .A1(n140), .A2(n132), .B1(n138), .B2(i_data_bus[11]), .ZN(N298) );
  INVD1BWP30P140 U179 ( .I(i_data_bus[54]), .ZN(n133) );
  MOAI22D1BWP30P140 U180 ( .A1(n140), .A2(n133), .B1(n138), .B2(i_data_bus[22]), .ZN(N309) );
  INVD1BWP30P140 U181 ( .I(i_data_bus[42]), .ZN(n134) );
  MOAI22D1BWP30P140 U182 ( .A1(n140), .A2(n134), .B1(n138), .B2(i_data_bus[10]), .ZN(N297) );
  INVD1BWP30P140 U183 ( .I(i_data_bus[53]), .ZN(n135) );
  MOAI22D1BWP30P140 U184 ( .A1(n140), .A2(n135), .B1(n138), .B2(i_data_bus[21]), .ZN(N308) );
  INVD1BWP30P140 U185 ( .I(i_data_bus[41]), .ZN(n136) );
  MOAI22D1BWP30P140 U186 ( .A1(n140), .A2(n136), .B1(n138), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140 U187 ( .I(i_data_bus[52]), .ZN(n137) );
  MOAI22D1BWP30P140 U188 ( .A1(n140), .A2(n137), .B1(n138), .B2(i_data_bus[20]), .ZN(N307) );
  INVD1BWP30P140 U189 ( .I(i_data_bus[40]), .ZN(n139) );
  MOAI22D1BWP30P140 U190 ( .A1(n140), .A2(n139), .B1(n9), .B2(i_data_bus[8]), 
        .ZN(N295) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_55 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n8, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(o_data_bus[2]) );
  DFD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(o_data_bus[8]) );
  DFD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(o_data_bus[9]) );
  DFD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  INVD3BWP30P140 U3 ( .I(n35), .ZN(n124) );
  NR2D4BWP30P140 U4 ( .A1(n31), .A2(n30), .ZN(n35) );
  NR2D1BWP30P140 U5 ( .A1(i_cmd[1]), .A2(n109), .ZN(n42) );
  INVD6BWP30P140 U6 ( .I(n57), .ZN(n1) );
  ND2OPTPAD1BWP30P140 U7 ( .A1(i_cmd[0]), .A2(n29), .ZN(n30) );
  MUX2NOPTD2BWP30P140 U8 ( .I0(i_valid[0]), .I1(i_valid[1]), .S(i_cmd[1]), 
        .ZN(n31) );
  MUX2NOPTD2BWP30P140 U9 ( .I0(i_valid[0]), .I1(i_valid[1]), .S(i_cmd[0]), 
        .ZN(n41) );
  OR2D8BWP30P140 U10 ( .A1(n32), .A2(i_cmd[0]), .Z(n126) );
  CKND2D4BWP30P140 U11 ( .A1(i_valid[0]), .A2(n29), .ZN(n32) );
  INVD1BWP30P140 U12 ( .I(n126), .ZN(n8) );
  INVD8BWP30P140 U13 ( .I(n126), .ZN(n145) );
  INVD1BWP30P140 U14 ( .I(n32), .ZN(n114) );
  INVD1BWP30P140 U15 ( .I(i_cmd[0]), .ZN(n112) );
  ND3OPTPAD2BWP30P140 U16 ( .A1(i_cmd[1]), .A2(i_valid[1]), .A3(n29), .ZN(n115) );
  ND2D1BWP30P140 U17 ( .A1(n28), .A2(i_en), .ZN(n109) );
  ND2D1BWP30P140 U18 ( .A1(n126), .A2(n113), .ZN(N353) );
  IND2D1BWP30P140 U19 ( .A1(n112), .B1(n111), .ZN(n113) );
  NR2D1BWP30P140 U20 ( .A1(n110), .A2(n109), .ZN(n111) );
  INVD1BWP30P140 U21 ( .I(i_valid[1]), .ZN(n110) );
  OAI21D1BWP30P140 U22 ( .A1(n124), .A2(n108), .B(n107), .ZN(N287) );
  OAI21D1BWP30P140 U23 ( .A1(n124), .A2(n106), .B(n105), .ZN(N288) );
  ND2D1BWP30P140 U24 ( .A1(n8), .A2(i_data_bus[1]), .ZN(n105) );
  OAI22D1BWP30P140 U25 ( .A1(n126), .A2(n67), .B1(n124), .B2(n36), .ZN(N292)
         );
  OAI22D1BWP30P140 U26 ( .A1(n147), .A2(n38), .B1(n126), .B2(n83), .ZN(N305)
         );
  OAI22D1BWP30P140 U27 ( .A1(n147), .A2(n37), .B1(n126), .B2(n85), .ZN(N306)
         );
  OAI22D1BWP30P140 U28 ( .A1(n147), .A2(n40), .B1(n126), .B2(n46), .ZN(N317)
         );
  OAI22D1BWP30P140 U29 ( .A1(n147), .A2(n39), .B1(n126), .B2(n44), .ZN(N318)
         );
  ND2D1BWP30P140 U30 ( .A1(n102), .A2(i_data_bus[50]), .ZN(n82) );
  ND2D1BWP30P140 U31 ( .A1(n102), .A2(i_data_bus[51]), .ZN(n84) );
  ND2D1BWP30P140 U32 ( .A1(n102), .A2(i_data_bus[52]), .ZN(n86) );
  ND2D1BWP30P140 U33 ( .A1(n102), .A2(i_data_bus[53]), .ZN(n88) );
  ND2D1BWP30P140 U34 ( .A1(n102), .A2(i_data_bus[54]), .ZN(n103) );
  ND2D1BWP30P140 U35 ( .A1(n102), .A2(i_data_bus[55]), .ZN(n98) );
  ND2D1BWP30P140 U36 ( .A1(n102), .A2(i_data_bus[56]), .ZN(n96) );
  ND2D1BWP30P140 U37 ( .A1(n102), .A2(i_data_bus[57]), .ZN(n55) );
  ND2D1BWP30P140 U38 ( .A1(n102), .A2(i_data_bus[58]), .ZN(n53) );
  ND2D1BWP30P140 U39 ( .A1(n102), .A2(i_data_bus[59]), .ZN(n51) );
  ND2D1BWP30P140 U40 ( .A1(n102), .A2(i_data_bus[60]), .ZN(n49) );
  ND2D1BWP30P140 U41 ( .A1(n102), .A2(i_data_bus[61]), .ZN(n47) );
  ND2D1BWP30P140 U42 ( .A1(n102), .A2(i_data_bus[62]), .ZN(n45) );
  ND2D1BWP30P140 U43 ( .A1(n102), .A2(i_data_bus[63]), .ZN(n43) );
  INR2D4BWP30P140 U44 ( .A1(n42), .B1(n41), .ZN(n57) );
  INVD1BWP30P140 U45 ( .I(n109), .ZN(n29) );
  INVD1BWP30P140 U46 ( .I(rst), .ZN(n28) );
  INVD6BWP30P140 U47 ( .I(n35), .ZN(n147) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[49]), .ZN(n33) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[17]), .ZN(n93) );
  OAI22D1BWP30P140 U50 ( .A1(n147), .A2(n33), .B1(n126), .B2(n93), .ZN(N304)
         );
  INVD1BWP30P140 U51 ( .I(i_data_bus[61]), .ZN(n34) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[29]), .ZN(n48) );
  OAI22D1BWP30P140 U53 ( .A1(n147), .A2(n34), .B1(n126), .B2(n48), .ZN(N316)
         );
  INVD1BWP30P140 U54 ( .I(i_data_bus[5]), .ZN(n67) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[37]), .ZN(n36) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[51]), .ZN(n37) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[19]), .ZN(n85) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[50]), .ZN(n38) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[18]), .ZN(n83) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[63]), .ZN(n39) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[31]), .ZN(n44) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[62]), .ZN(n40) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[30]), .ZN(n46) );
  INVD6BWP30P140 U64 ( .I(n115), .ZN(n102) );
  OAI21D1BWP30P140 U65 ( .A1(n1), .A2(n44), .B(n43), .ZN(N350) );
  OAI21D1BWP30P140 U66 ( .A1(n1), .A2(n46), .B(n45), .ZN(N349) );
  OAI21D1BWP30P140 U67 ( .A1(n1), .A2(n48), .B(n47), .ZN(N348) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[28]), .ZN(n50) );
  OAI21D1BWP30P140 U69 ( .A1(n1), .A2(n50), .B(n49), .ZN(N347) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[27]), .ZN(n52) );
  OAI21D1BWP30P140 U71 ( .A1(n1), .A2(n52), .B(n51), .ZN(N346) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[26]), .ZN(n54) );
  OAI21D1BWP30P140 U73 ( .A1(n1), .A2(n54), .B(n53), .ZN(N345) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[25]), .ZN(n56) );
  OAI21D1BWP30P140 U75 ( .A1(n1), .A2(n56), .B(n55), .ZN(N344) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[0]), .ZN(n59) );
  ND2OPTIBD1BWP30P140 U77 ( .A1(n102), .A2(i_data_bus[32]), .ZN(n58) );
  OAI21D1BWP30P140 U78 ( .A1(n1), .A2(n59), .B(n58), .ZN(N319) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[1]), .ZN(n61) );
  ND2OPTIBD1BWP30P140 U80 ( .A1(n102), .A2(i_data_bus[33]), .ZN(n60) );
  OAI21D1BWP30P140 U81 ( .A1(n1), .A2(n61), .B(n60), .ZN(N320) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[2]), .ZN(n63) );
  ND2OPTIBD1BWP30P140 U83 ( .A1(n102), .A2(i_data_bus[34]), .ZN(n62) );
  OAI21D1BWP30P140 U84 ( .A1(n1), .A2(n63), .B(n62), .ZN(N321) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[3]), .ZN(n125) );
  ND2OPTIBD1BWP30P140 U86 ( .A1(n102), .A2(i_data_bus[35]), .ZN(n64) );
  OAI21D1BWP30P140 U87 ( .A1(n1), .A2(n125), .B(n64), .ZN(N322) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[4]), .ZN(n122) );
  ND2OPTIBD1BWP30P140 U89 ( .A1(n102), .A2(i_data_bus[36]), .ZN(n65) );
  OAI21D1BWP30P140 U90 ( .A1(n1), .A2(n122), .B(n65), .ZN(N323) );
  ND2OPTIBD1BWP30P140 U91 ( .A1(n102), .A2(i_data_bus[37]), .ZN(n66) );
  OAI21D1BWP30P140 U92 ( .A1(n1), .A2(n67), .B(n66), .ZN(N324) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[6]), .ZN(n120) );
  ND2OPTIBD1BWP30P140 U94 ( .A1(n102), .A2(i_data_bus[38]), .ZN(n68) );
  OAI21D1BWP30P140 U95 ( .A1(n1), .A2(n120), .B(n68), .ZN(N325) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[7]), .ZN(n118) );
  ND2OPTIBD1BWP30P140 U97 ( .A1(n102), .A2(i_data_bus[39]), .ZN(n69) );
  OAI21D1BWP30P140 U98 ( .A1(n1), .A2(n118), .B(n69), .ZN(N326) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[8]), .ZN(n71) );
  ND2OPTIBD1BWP30P140 U100 ( .A1(n102), .A2(i_data_bus[40]), .ZN(n70) );
  OAI21D1BWP30P140 U101 ( .A1(n1), .A2(n71), .B(n70), .ZN(N327) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[9]), .ZN(n73) );
  ND2OPTIBD1BWP30P140 U103 ( .A1(n102), .A2(i_data_bus[41]), .ZN(n72) );
  OAI21D1BWP30P140 U104 ( .A1(n1), .A2(n73), .B(n72), .ZN(N328) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[10]), .ZN(n75) );
  ND2OPTIBD1BWP30P140 U106 ( .A1(n102), .A2(i_data_bus[42]), .ZN(n74) );
  OAI21D1BWP30P140 U107 ( .A1(n1), .A2(n75), .B(n74), .ZN(N329) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[11]), .ZN(n77) );
  ND2OPTIBD1BWP30P140 U109 ( .A1(n102), .A2(i_data_bus[43]), .ZN(n76) );
  OAI21D1BWP30P140 U110 ( .A1(n1), .A2(n77), .B(n76), .ZN(N330) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[12]), .ZN(n79) );
  ND2OPTIBD1BWP30P140 U112 ( .A1(n102), .A2(i_data_bus[44]), .ZN(n78) );
  OAI21D1BWP30P140 U113 ( .A1(n1), .A2(n79), .B(n78), .ZN(N331) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[13]), .ZN(n81) );
  ND2OPTIBD1BWP30P140 U115 ( .A1(n102), .A2(i_data_bus[45]), .ZN(n80) );
  OAI21D1BWP30P140 U116 ( .A1(n1), .A2(n81), .B(n80), .ZN(N332) );
  OAI21D1BWP30P140 U117 ( .A1(n1), .A2(n83), .B(n82), .ZN(N337) );
  OAI21D1BWP30P140 U118 ( .A1(n1), .A2(n85), .B(n84), .ZN(N338) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[20]), .ZN(n87) );
  OAI21D1BWP30P140 U120 ( .A1(n1), .A2(n87), .B(n86), .ZN(N339) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[21]), .ZN(n89) );
  OAI21D1BWP30P140 U122 ( .A1(n1), .A2(n89), .B(n88), .ZN(N340) );
  INVD1BWP30P140 U123 ( .I(i_data_bus[16]), .ZN(n91) );
  ND2OPTIBD1BWP30P140 U124 ( .A1(n102), .A2(i_data_bus[48]), .ZN(n90) );
  OAI21D1BWP30P140 U125 ( .A1(n1), .A2(n91), .B(n90), .ZN(N335) );
  ND2OPTIBD1BWP30P140 U126 ( .A1(n102), .A2(i_data_bus[49]), .ZN(n92) );
  OAI21D1BWP30P140 U127 ( .A1(n1), .A2(n93), .B(n92), .ZN(N336) );
  INVD1BWP30P140 U128 ( .I(i_data_bus[15]), .ZN(n95) );
  ND2OPTIBD1BWP30P140 U129 ( .A1(n102), .A2(i_data_bus[47]), .ZN(n94) );
  OAI21D1BWP30P140 U130 ( .A1(n1), .A2(n95), .B(n94), .ZN(N334) );
  INVD1BWP30P140 U131 ( .I(i_data_bus[24]), .ZN(n97) );
  OAI21D1BWP30P140 U132 ( .A1(n1), .A2(n97), .B(n96), .ZN(N343) );
  INVD1BWP30P140 U133 ( .I(i_data_bus[23]), .ZN(n99) );
  OAI21D1BWP30P140 U134 ( .A1(n1), .A2(n99), .B(n98), .ZN(N342) );
  INVD1BWP30P140 U135 ( .I(i_data_bus[14]), .ZN(n101) );
  ND2OPTIBD1BWP30P140 U136 ( .A1(n102), .A2(i_data_bus[46]), .ZN(n100) );
  OAI21D1BWP30P140 U137 ( .A1(n1), .A2(n101), .B(n100), .ZN(N333) );
  INVD1BWP30P140 U138 ( .I(i_data_bus[22]), .ZN(n104) );
  OAI21D1BWP30P140 U139 ( .A1(n1), .A2(n104), .B(n103), .ZN(N341) );
  INVD1BWP30P140 U140 ( .I(i_data_bus[33]), .ZN(n106) );
  INVD1BWP30P140 U141 ( .I(i_data_bus[32]), .ZN(n108) );
  IND2D2BWP30P140 U142 ( .A1(n126), .B1(i_data_bus[0]), .ZN(n107) );
  INVD1BWP30P140 U143 ( .I(n114), .ZN(n116) );
  OAI21D1BWP30P140 U144 ( .A1(n116), .A2(i_cmd[1]), .B(n115), .ZN(N354) );
  INVD1BWP30P140 U145 ( .I(i_data_bus[39]), .ZN(n117) );
  OAI22D1BWP30P140 U146 ( .A1(n126), .A2(n118), .B1(n124), .B2(n117), .ZN(N294) );
  INVD1BWP30P140 U147 ( .I(i_data_bus[38]), .ZN(n119) );
  OAI22D1BWP30P140 U148 ( .A1(n126), .A2(n120), .B1(n124), .B2(n119), .ZN(N293) );
  INVD1BWP30P140 U149 ( .I(i_data_bus[36]), .ZN(n121) );
  OAI22D1BWP30P140 U150 ( .A1(n126), .A2(n122), .B1(n124), .B2(n121), .ZN(N291) );
  INVD1BWP30P140 U151 ( .I(i_data_bus[35]), .ZN(n123) );
  OAI22D1BWP30P140 U152 ( .A1(n126), .A2(n125), .B1(n124), .B2(n123), .ZN(N290) );
  INVD1BWP30P140 U153 ( .I(i_data_bus[60]), .ZN(n127) );
  MOAI22D1BWP30P140 U154 ( .A1(n147), .A2(n127), .B1(n145), .B2(i_data_bus[28]), .ZN(N315) );
  INVD1BWP30P140 U155 ( .I(i_data_bus[48]), .ZN(n128) );
  MOAI22D1BWP30P140 U156 ( .A1(n147), .A2(n128), .B1(n145), .B2(i_data_bus[16]), .ZN(N303) );
  INVD1BWP30P140 U157 ( .I(i_data_bus[34]), .ZN(n129) );
  MOAI22D1BWP30P140 U158 ( .A1(n147), .A2(n129), .B1(n145), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140 U159 ( .I(i_data_bus[59]), .ZN(n130) );
  MOAI22D1BWP30P140 U160 ( .A1(n147), .A2(n130), .B1(n145), .B2(i_data_bus[27]), .ZN(N314) );
  INVD1BWP30P140 U161 ( .I(i_data_bus[47]), .ZN(n131) );
  MOAI22D1BWP30P140 U162 ( .A1(n147), .A2(n131), .B1(n145), .B2(i_data_bus[15]), .ZN(N302) );
  INVD1BWP30P140 U163 ( .I(i_data_bus[58]), .ZN(n132) );
  MOAI22D1BWP30P140 U164 ( .A1(n147), .A2(n132), .B1(n145), .B2(i_data_bus[26]), .ZN(N313) );
  INVD1BWP30P140 U165 ( .I(i_data_bus[46]), .ZN(n133) );
  MOAI22D1BWP30P140 U166 ( .A1(n147), .A2(n133), .B1(n145), .B2(i_data_bus[14]), .ZN(N301) );
  INVD1BWP30P140 U167 ( .I(i_data_bus[57]), .ZN(n134) );
  MOAI22D1BWP30P140 U168 ( .A1(n147), .A2(n134), .B1(n145), .B2(i_data_bus[25]), .ZN(N312) );
  INVD1BWP30P140 U169 ( .I(i_data_bus[45]), .ZN(n135) );
  MOAI22D1BWP30P140 U170 ( .A1(n147), .A2(n135), .B1(n145), .B2(i_data_bus[13]), .ZN(N300) );
  INVD1BWP30P140 U171 ( .I(i_data_bus[56]), .ZN(n136) );
  MOAI22D1BWP30P140 U172 ( .A1(n147), .A2(n136), .B1(n145), .B2(i_data_bus[24]), .ZN(N311) );
  INVD1BWP30P140 U173 ( .I(i_data_bus[44]), .ZN(n137) );
  MOAI22D1BWP30P140 U174 ( .A1(n147), .A2(n137), .B1(n145), .B2(i_data_bus[12]), .ZN(N299) );
  INVD1BWP30P140 U175 ( .I(i_data_bus[55]), .ZN(n138) );
  MOAI22D1BWP30P140 U176 ( .A1(n147), .A2(n138), .B1(n145), .B2(i_data_bus[23]), .ZN(N310) );
  INVD1BWP30P140 U177 ( .I(i_data_bus[43]), .ZN(n139) );
  MOAI22D1BWP30P140 U178 ( .A1(n147), .A2(n139), .B1(n145), .B2(i_data_bus[11]), .ZN(N298) );
  INVD1BWP30P140 U179 ( .I(i_data_bus[54]), .ZN(n140) );
  MOAI22D1BWP30P140 U180 ( .A1(n147), .A2(n140), .B1(n145), .B2(i_data_bus[22]), .ZN(N309) );
  INVD1BWP30P140 U181 ( .I(i_data_bus[42]), .ZN(n141) );
  MOAI22D1BWP30P140 U182 ( .A1(n147), .A2(n141), .B1(n145), .B2(i_data_bus[10]), .ZN(N297) );
  INVD1BWP30P140 U183 ( .I(i_data_bus[53]), .ZN(n142) );
  MOAI22D1BWP30P140 U184 ( .A1(n147), .A2(n142), .B1(n145), .B2(i_data_bus[21]), .ZN(N308) );
  INVD1BWP30P140 U185 ( .I(i_data_bus[41]), .ZN(n143) );
  MOAI22D1BWP30P140 U186 ( .A1(n147), .A2(n143), .B1(n145), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140 U187 ( .I(i_data_bus[52]), .ZN(n144) );
  MOAI22D1BWP30P140 U188 ( .A1(n147), .A2(n144), .B1(n145), .B2(i_data_bus[20]), .ZN(N307) );
  INVD1BWP30P140 U189 ( .I(i_data_bus[40]), .ZN(n146) );
  MOAI22D1BWP30P140 U190 ( .A1(n147), .A2(n146), .B1(n145), .B2(i_data_bus[8]), 
        .ZN(N295) );
endmodule


module benes_simple_seq ( clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, 
        i_en, i_cmd );
  input [15:0] i_valid;
  input [511:0] i_data_bus;
  output [15:0] o_valid;
  output [511:0] o_data_bus;
  input [111:0] i_cmd;
  input clk, rst, i_en;
  wire   n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, connection_0__0__31_,
         connection_0__0__30_, connection_0__0__29_, connection_0__0__28_,
         connection_0__0__27_, connection_0__0__26_, connection_0__0__25_,
         connection_0__0__24_, connection_0__0__23_, connection_0__0__22_,
         connection_0__0__21_, connection_0__0__20_, connection_0__0__19_,
         connection_0__0__18_, connection_0__0__17_, connection_0__0__16_,
         connection_0__0__15_, connection_0__0__14_, connection_0__0__13_,
         connection_0__0__12_, connection_0__0__11_, connection_0__0__10_,
         connection_0__0__9_, connection_0__0__8_, connection_0__0__7_,
         connection_0__0__6_, connection_0__0__5_, connection_0__0__4_,
         connection_0__0__3_, connection_0__0__2_, connection_0__0__1_,
         connection_0__0__0_, connection_0__1__31_, connection_0__1__30_,
         connection_0__1__29_, connection_0__1__28_, connection_0__1__27_,
         connection_0__1__26_, connection_0__1__25_, connection_0__1__24_,
         connection_0__1__23_, connection_0__1__22_, connection_0__1__21_,
         connection_0__1__20_, connection_0__1__19_, connection_0__1__18_,
         connection_0__1__17_, connection_0__1__16_, connection_0__1__15_,
         connection_0__1__14_, connection_0__1__13_, connection_0__1__12_,
         connection_0__1__11_, connection_0__1__10_, connection_0__1__9_,
         connection_0__1__8_, connection_0__1__7_, connection_0__1__6_,
         connection_0__1__5_, connection_0__1__4_, connection_0__1__3_,
         connection_0__1__2_, connection_0__1__1_, connection_0__1__0_,
         connection_0__2__31_, connection_0__2__30_, connection_0__2__29_,
         connection_0__2__28_, connection_0__2__27_, connection_0__2__26_,
         connection_0__2__25_, connection_0__2__24_, connection_0__2__23_,
         connection_0__2__22_, connection_0__2__21_, connection_0__2__20_,
         connection_0__2__19_, connection_0__2__18_, connection_0__2__17_,
         connection_0__2__16_, connection_0__2__15_, connection_0__2__14_,
         connection_0__2__13_, connection_0__2__12_, connection_0__2__11_,
         connection_0__2__10_, connection_0__2__9_, connection_0__2__8_,
         connection_0__2__7_, connection_0__2__6_, connection_0__2__5_,
         connection_0__2__4_, connection_0__2__3_, connection_0__2__2_,
         connection_0__2__1_, connection_0__2__0_, connection_0__3__31_,
         connection_0__3__30_, connection_0__3__29_, connection_0__3__28_,
         connection_0__3__27_, connection_0__3__26_, connection_0__3__25_,
         connection_0__3__24_, connection_0__3__23_, connection_0__3__22_,
         connection_0__3__21_, connection_0__3__20_, connection_0__3__19_,
         connection_0__3__18_, connection_0__3__17_, connection_0__3__16_,
         connection_0__3__15_, connection_0__3__14_, connection_0__3__13_,
         connection_0__3__12_, connection_0__3__11_, connection_0__3__10_,
         connection_0__3__9_, connection_0__3__8_, connection_0__3__7_,
         connection_0__3__6_, connection_0__3__5_, connection_0__3__4_,
         connection_0__3__3_, connection_0__3__2_, connection_0__3__1_,
         connection_0__3__0_, connection_0__4__31_, connection_0__4__30_,
         connection_0__4__29_, connection_0__4__28_, connection_0__4__27_,
         connection_0__4__26_, connection_0__4__25_, connection_0__4__24_,
         connection_0__4__23_, connection_0__4__22_, connection_0__4__21_,
         connection_0__4__20_, connection_0__4__19_, connection_0__4__18_,
         connection_0__4__17_, connection_0__4__16_, connection_0__4__15_,
         connection_0__4__14_, connection_0__4__13_, connection_0__4__12_,
         connection_0__4__11_, connection_0__4__10_, connection_0__4__9_,
         connection_0__4__8_, connection_0__4__7_, connection_0__4__6_,
         connection_0__4__5_, connection_0__4__4_, connection_0__4__3_,
         connection_0__4__2_, connection_0__4__1_, connection_0__4__0_,
         connection_0__5__31_, connection_0__5__30_, connection_0__5__29_,
         connection_0__5__28_, connection_0__5__27_, connection_0__5__26_,
         connection_0__5__25_, connection_0__5__24_, connection_0__5__23_,
         connection_0__5__22_, connection_0__5__21_, connection_0__5__20_,
         connection_0__5__19_, connection_0__5__18_, connection_0__5__17_,
         connection_0__5__16_, connection_0__5__15_, connection_0__5__14_,
         connection_0__5__13_, connection_0__5__12_, connection_0__5__11_,
         connection_0__5__10_, connection_0__5__9_, connection_0__5__8_,
         connection_0__5__7_, connection_0__5__6_, connection_0__5__5_,
         connection_0__5__4_, connection_0__5__3_, connection_0__5__2_,
         connection_0__5__1_, connection_0__5__0_, connection_0__6__31_,
         connection_0__6__30_, connection_0__6__29_, connection_0__6__28_,
         connection_0__6__27_, connection_0__6__26_, connection_0__6__25_,
         connection_0__6__24_, connection_0__6__23_, connection_0__6__22_,
         connection_0__6__21_, connection_0__6__20_, connection_0__6__19_,
         connection_0__6__18_, connection_0__6__17_, connection_0__6__16_,
         connection_0__6__15_, connection_0__6__14_, connection_0__6__13_,
         connection_0__6__12_, connection_0__6__11_, connection_0__6__10_,
         connection_0__6__9_, connection_0__6__8_, connection_0__6__7_,
         connection_0__6__6_, connection_0__6__5_, connection_0__6__4_,
         connection_0__6__3_, connection_0__6__2_, connection_0__6__1_,
         connection_0__6__0_, connection_0__7__31_, connection_0__7__30_,
         connection_0__7__29_, connection_0__7__28_, connection_0__7__27_,
         connection_0__7__26_, connection_0__7__25_, connection_0__7__24_,
         connection_0__7__23_, connection_0__7__22_, connection_0__7__21_,
         connection_0__7__20_, connection_0__7__19_, connection_0__7__18_,
         connection_0__7__17_, connection_0__7__16_, connection_0__7__15_,
         connection_0__7__14_, connection_0__7__13_, connection_0__7__12_,
         connection_0__7__11_, connection_0__7__10_, connection_0__7__9_,
         connection_0__7__8_, connection_0__7__7_, connection_0__7__6_,
         connection_0__7__5_, connection_0__7__4_, connection_0__7__3_,
         connection_0__7__2_, connection_0__7__1_, connection_0__7__0_,
         connection_0__8__31_, connection_0__8__30_, connection_0__8__29_,
         connection_0__8__28_, connection_0__8__27_, connection_0__8__26_,
         connection_0__8__25_, connection_0__8__24_, connection_0__8__23_,
         connection_0__8__22_, connection_0__8__21_, connection_0__8__20_,
         connection_0__8__19_, connection_0__8__18_, connection_0__8__17_,
         connection_0__8__16_, connection_0__8__15_, connection_0__8__14_,
         connection_0__8__13_, connection_0__8__12_, connection_0__8__11_,
         connection_0__8__10_, connection_0__8__9_, connection_0__8__8_,
         connection_0__8__7_, connection_0__8__6_, connection_0__8__5_,
         connection_0__8__4_, connection_0__8__3_, connection_0__8__2_,
         connection_0__8__1_, connection_0__8__0_, connection_0__9__31_,
         connection_0__9__30_, connection_0__9__29_, connection_0__9__28_,
         connection_0__9__27_, connection_0__9__26_, connection_0__9__25_,
         connection_0__9__24_, connection_0__9__23_, connection_0__9__22_,
         connection_0__9__21_, connection_0__9__20_, connection_0__9__19_,
         connection_0__9__18_, connection_0__9__17_, connection_0__9__16_,
         connection_0__9__15_, connection_0__9__14_, connection_0__9__13_,
         connection_0__9__12_, connection_0__9__11_, connection_0__9__10_,
         connection_0__9__9_, connection_0__9__8_, connection_0__9__7_,
         connection_0__9__6_, connection_0__9__5_, connection_0__9__4_,
         connection_0__9__3_, connection_0__9__2_, connection_0__9__1_,
         connection_0__9__0_, connection_0__10__31_, connection_0__10__30_,
         connection_0__10__29_, connection_0__10__28_, connection_0__10__27_,
         connection_0__10__26_, connection_0__10__25_, connection_0__10__24_,
         connection_0__10__23_, connection_0__10__22_, connection_0__10__21_,
         connection_0__10__20_, connection_0__10__19_, connection_0__10__18_,
         connection_0__10__17_, connection_0__10__16_, connection_0__10__15_,
         connection_0__10__14_, connection_0__10__13_, connection_0__10__12_,
         connection_0__10__11_, connection_0__10__10_, connection_0__10__9_,
         connection_0__10__8_, connection_0__10__7_, connection_0__10__6_,
         connection_0__10__5_, connection_0__10__4_, connection_0__10__3_,
         connection_0__10__2_, connection_0__10__1_, connection_0__10__0_,
         connection_0__11__31_, connection_0__11__30_, connection_0__11__29_,
         connection_0__11__28_, connection_0__11__27_, connection_0__11__26_,
         connection_0__11__25_, connection_0__11__24_, connection_0__11__23_,
         connection_0__11__22_, connection_0__11__21_, connection_0__11__20_,
         connection_0__11__19_, connection_0__11__18_, connection_0__11__17_,
         connection_0__11__16_, connection_0__11__15_, connection_0__11__14_,
         connection_0__11__13_, connection_0__11__12_, connection_0__11__11_,
         connection_0__11__10_, connection_0__11__9_, connection_0__11__8_,
         connection_0__11__7_, connection_0__11__6_, connection_0__11__5_,
         connection_0__11__4_, connection_0__11__3_, connection_0__11__2_,
         connection_0__11__1_, connection_0__11__0_, connection_0__12__31_,
         connection_0__12__30_, connection_0__12__29_, connection_0__12__28_,
         connection_0__12__27_, connection_0__12__26_, connection_0__12__25_,
         connection_0__12__24_, connection_0__12__23_, connection_0__12__22_,
         connection_0__12__21_, connection_0__12__20_, connection_0__12__19_,
         connection_0__12__18_, connection_0__12__17_, connection_0__12__16_,
         connection_0__12__15_, connection_0__12__14_, connection_0__12__13_,
         connection_0__12__12_, connection_0__12__11_, connection_0__12__10_,
         connection_0__12__9_, connection_0__12__8_, connection_0__12__7_,
         connection_0__12__6_, connection_0__12__5_, connection_0__12__4_,
         connection_0__12__3_, connection_0__12__2_, connection_0__12__1_,
         connection_0__12__0_, connection_0__13__31_, connection_0__13__30_,
         connection_0__13__29_, connection_0__13__28_, connection_0__13__27_,
         connection_0__13__26_, connection_0__13__25_, connection_0__13__24_,
         connection_0__13__23_, connection_0__13__22_, connection_0__13__21_,
         connection_0__13__20_, connection_0__13__19_, connection_0__13__18_,
         connection_0__13__17_, connection_0__13__16_, connection_0__13__15_,
         connection_0__13__14_, connection_0__13__13_, connection_0__13__12_,
         connection_0__13__11_, connection_0__13__10_, connection_0__13__9_,
         connection_0__13__8_, connection_0__13__7_, connection_0__13__6_,
         connection_0__13__5_, connection_0__13__4_, connection_0__13__3_,
         connection_0__13__2_, connection_0__13__1_, connection_0__13__0_,
         connection_0__14__31_, connection_0__14__30_, connection_0__14__29_,
         connection_0__14__28_, connection_0__14__27_, connection_0__14__26_,
         connection_0__14__25_, connection_0__14__24_, connection_0__14__23_,
         connection_0__14__22_, connection_0__14__21_, connection_0__14__20_,
         connection_0__14__19_, connection_0__14__18_, connection_0__14__17_,
         connection_0__14__16_, connection_0__14__15_, connection_0__14__14_,
         connection_0__14__13_, connection_0__14__12_, connection_0__14__11_,
         connection_0__14__10_, connection_0__14__9_, connection_0__14__8_,
         connection_0__14__7_, connection_0__14__6_, connection_0__14__5_,
         connection_0__14__4_, connection_0__14__3_, connection_0__14__2_,
         connection_0__14__1_, connection_0__14__0_, connection_0__15__31_,
         connection_0__15__30_, connection_0__15__29_, connection_0__15__28_,
         connection_0__15__27_, connection_0__15__26_, connection_0__15__25_,
         connection_0__15__24_, connection_0__15__23_, connection_0__15__22_,
         connection_0__15__21_, connection_0__15__20_, connection_0__15__19_,
         connection_0__15__18_, connection_0__15__17_, connection_0__15__16_,
         connection_0__15__15_, connection_0__15__14_, connection_0__15__13_,
         connection_0__15__12_, connection_0__15__11_, connection_0__15__10_,
         connection_0__15__9_, connection_0__15__8_, connection_0__15__7_,
         connection_0__15__6_, connection_0__15__5_, connection_0__15__4_,
         connection_0__15__3_, connection_0__15__2_, connection_0__15__1_,
         connection_0__15__0_, connection_valid_0__0_, connection_valid_0__1_,
         connection_valid_0__2_, connection_valid_0__3_,
         connection_valid_0__4_, connection_valid_0__5_,
         connection_valid_0__6_, connection_valid_0__7_,
         connection_valid_0__8_, connection_valid_0__9_,
         connection_valid_0__10_, connection_valid_0__11_,
         connection_valid_0__12_, connection_valid_0__13_,
         connection_valid_0__14_, connection_valid_0__15_,
         connection_valid_1__0_, connection_valid_1__1_,
         connection_valid_1__2_, connection_valid_1__3_,
         connection_valid_1__4_, connection_valid_1__5_,
         connection_valid_1__6_, connection_valid_1__7_,
         connection_valid_1__8_, connection_valid_1__9_,
         connection_valid_1__10_, connection_valid_1__11_,
         connection_valid_1__12_, connection_valid_1__13_,
         connection_valid_1__14_, connection_valid_1__15_,
         connection_valid_2__0_, connection_valid_2__1_,
         connection_valid_2__2_, connection_valid_2__3_,
         connection_valid_2__4_, connection_valid_2__5_,
         connection_valid_2__6_, connection_valid_2__7_,
         connection_valid_2__8_, connection_valid_2__9_,
         connection_valid_2__10_, connection_valid_2__11_,
         connection_valid_2__12_, connection_valid_2__13_,
         connection_valid_2__14_, connection_valid_2__15_,
         connection_valid_3__0_, connection_valid_3__1_,
         connection_valid_3__2_, connection_valid_3__3_,
         connection_valid_3__4_, connection_valid_3__5_,
         connection_valid_3__6_, connection_valid_3__7_,
         connection_valid_3__8_, connection_valid_3__9_,
         connection_valid_3__10_, connection_valid_3__11_,
         connection_valid_3__12_, connection_valid_3__13_,
         connection_valid_3__14_, connection_valid_3__15_,
         connection_valid_4__0_, connection_valid_4__1_,
         connection_valid_4__2_, connection_valid_4__3_,
         connection_valid_4__4_, connection_valid_4__5_,
         connection_valid_4__6_, connection_valid_4__7_,
         connection_valid_4__8_, connection_valid_4__9_,
         connection_valid_4__10_, connection_valid_4__11_,
         connection_valid_4__12_, connection_valid_4__13_,
         connection_valid_4__14_, connection_valid_4__15_,
         connection_valid_5__0_, connection_valid_5__1_,
         connection_valid_5__2_, connection_valid_5__3_,
         connection_valid_5__4_, connection_valid_5__5_,
         connection_valid_5__6_, connection_valid_5__7_,
         connection_valid_5__8_, connection_valid_5__9_,
         connection_valid_5__10_, connection_valid_5__11_,
         connection_valid_5__12_, connection_valid_5__13_,
         connection_valid_5__14_, connection_valid_5__15_,
         connection_1__0__31_, connection_1__0__30_, connection_1__0__29_,
         connection_1__0__28_, connection_1__0__27_, connection_1__0__26_,
         connection_1__0__25_, connection_1__0__24_, connection_1__0__23_,
         connection_1__0__22_, connection_1__0__21_, connection_1__0__20_,
         connection_1__0__19_, connection_1__0__18_, connection_1__0__17_,
         connection_1__0__16_, connection_1__0__15_, connection_1__0__14_,
         connection_1__0__13_, connection_1__0__12_, connection_1__0__11_,
         connection_1__0__10_, connection_1__0__9_, connection_1__0__8_,
         connection_1__0__7_, connection_1__0__6_, connection_1__0__5_,
         connection_1__0__4_, connection_1__0__3_, connection_1__0__2_,
         connection_1__0__1_, connection_1__0__0_, connection_1__1__31_,
         connection_1__1__30_, connection_1__1__29_, connection_1__1__28_,
         connection_1__1__27_, connection_1__1__26_, connection_1__1__25_,
         connection_1__1__24_, connection_1__1__23_, connection_1__1__22_,
         connection_1__1__21_, connection_1__1__20_, connection_1__1__19_,
         connection_1__1__18_, connection_1__1__17_, connection_1__1__16_,
         connection_1__1__15_, connection_1__1__14_, connection_1__1__13_,
         connection_1__1__12_, connection_1__1__11_, connection_1__1__10_,
         connection_1__1__9_, connection_1__1__8_, connection_1__1__7_,
         connection_1__1__6_, connection_1__1__5_, connection_1__1__4_,
         connection_1__1__3_, connection_1__1__2_, connection_1__1__1_,
         connection_1__1__0_, connection_1__2__31_, connection_1__2__30_,
         connection_1__2__29_, connection_1__2__28_, connection_1__2__27_,
         connection_1__2__26_, connection_1__2__25_, connection_1__2__24_,
         connection_1__2__23_, connection_1__2__22_, connection_1__2__21_,
         connection_1__2__20_, connection_1__2__19_, connection_1__2__18_,
         connection_1__2__17_, connection_1__2__16_, connection_1__2__15_,
         connection_1__2__14_, connection_1__2__13_, connection_1__2__12_,
         connection_1__2__11_, connection_1__2__10_, connection_1__2__9_,
         connection_1__2__8_, connection_1__2__7_, connection_1__2__6_,
         connection_1__2__5_, connection_1__2__4_, connection_1__2__3_,
         connection_1__2__2_, connection_1__2__1_, connection_1__2__0_,
         connection_1__3__31_, connection_1__3__30_, connection_1__3__29_,
         connection_1__3__28_, connection_1__3__27_, connection_1__3__26_,
         connection_1__3__25_, connection_1__3__24_, connection_1__3__23_,
         connection_1__3__22_, connection_1__3__21_, connection_1__3__20_,
         connection_1__3__19_, connection_1__3__18_, connection_1__3__17_,
         connection_1__3__16_, connection_1__3__15_, connection_1__3__14_,
         connection_1__3__13_, connection_1__3__12_, connection_1__3__11_,
         connection_1__3__10_, connection_1__3__9_, connection_1__3__8_,
         connection_1__3__7_, connection_1__3__6_, connection_1__3__5_,
         connection_1__3__4_, connection_1__3__3_, connection_1__3__2_,
         connection_1__3__1_, connection_1__3__0_, connection_1__4__31_,
         connection_1__4__30_, connection_1__4__29_, connection_1__4__28_,
         connection_1__4__27_, connection_1__4__26_, connection_1__4__25_,
         connection_1__4__24_, connection_1__4__23_, connection_1__4__22_,
         connection_1__4__21_, connection_1__4__20_, connection_1__4__19_,
         connection_1__4__18_, connection_1__4__17_, connection_1__4__16_,
         connection_1__4__15_, connection_1__4__14_, connection_1__4__13_,
         connection_1__4__12_, connection_1__4__11_, connection_1__4__10_,
         connection_1__4__9_, connection_1__4__8_, connection_1__4__7_,
         connection_1__4__6_, connection_1__4__5_, connection_1__4__4_,
         connection_1__4__3_, connection_1__4__2_, connection_1__4__1_,
         connection_1__4__0_, connection_1__5__31_, connection_1__5__30_,
         connection_1__5__29_, connection_1__5__28_, connection_1__5__27_,
         connection_1__5__26_, connection_1__5__25_, connection_1__5__24_,
         connection_1__5__23_, connection_1__5__22_, connection_1__5__21_,
         connection_1__5__20_, connection_1__5__19_, connection_1__5__18_,
         connection_1__5__17_, connection_1__5__16_, connection_1__5__15_,
         connection_1__5__14_, connection_1__5__13_, connection_1__5__12_,
         connection_1__5__11_, connection_1__5__10_, connection_1__5__9_,
         connection_1__5__8_, connection_1__5__7_, connection_1__5__6_,
         connection_1__5__5_, connection_1__5__4_, connection_1__5__3_,
         connection_1__5__2_, connection_1__5__1_, connection_1__5__0_,
         connection_1__6__31_, connection_1__6__30_, connection_1__6__29_,
         connection_1__6__28_, connection_1__6__27_, connection_1__6__26_,
         connection_1__6__25_, connection_1__6__24_, connection_1__6__23_,
         connection_1__6__22_, connection_1__6__21_, connection_1__6__20_,
         connection_1__6__19_, connection_1__6__18_, connection_1__6__17_,
         connection_1__6__16_, connection_1__6__15_, connection_1__6__14_,
         connection_1__6__13_, connection_1__6__12_, connection_1__6__11_,
         connection_1__6__10_, connection_1__6__9_, connection_1__6__8_,
         connection_1__6__7_, connection_1__6__6_, connection_1__6__5_,
         connection_1__6__4_, connection_1__6__3_, connection_1__6__2_,
         connection_1__6__1_, connection_1__6__0_, connection_1__7__31_,
         connection_1__7__30_, connection_1__7__29_, connection_1__7__28_,
         connection_1__7__27_, connection_1__7__26_, connection_1__7__25_,
         connection_1__7__24_, connection_1__7__23_, connection_1__7__22_,
         connection_1__7__21_, connection_1__7__20_, connection_1__7__19_,
         connection_1__7__18_, connection_1__7__17_, connection_1__7__16_,
         connection_1__7__15_, connection_1__7__14_, connection_1__7__13_,
         connection_1__7__12_, connection_1__7__11_, connection_1__7__10_,
         connection_1__7__9_, connection_1__7__8_, connection_1__7__7_,
         connection_1__7__6_, connection_1__7__5_, connection_1__7__4_,
         connection_1__7__3_, connection_1__7__2_, connection_1__7__1_,
         connection_1__7__0_, connection_1__8__31_, connection_1__8__30_,
         connection_1__8__29_, connection_1__8__28_, connection_1__8__27_,
         connection_1__8__26_, connection_1__8__25_, connection_1__8__24_,
         connection_1__8__23_, connection_1__8__22_, connection_1__8__21_,
         connection_1__8__20_, connection_1__8__19_, connection_1__8__18_,
         connection_1__8__17_, connection_1__8__16_, connection_1__8__15_,
         connection_1__8__14_, connection_1__8__13_, connection_1__8__12_,
         connection_1__8__11_, connection_1__8__10_, connection_1__8__9_,
         connection_1__8__8_, connection_1__8__7_, connection_1__8__6_,
         connection_1__8__5_, connection_1__8__4_, connection_1__8__3_,
         connection_1__8__2_, connection_1__8__1_, connection_1__8__0_,
         connection_1__9__31_, connection_1__9__30_, connection_1__9__29_,
         connection_1__9__28_, connection_1__9__27_, connection_1__9__26_,
         connection_1__9__25_, connection_1__9__24_, connection_1__9__23_,
         connection_1__9__22_, connection_1__9__21_, connection_1__9__20_,
         connection_1__9__19_, connection_1__9__18_, connection_1__9__17_,
         connection_1__9__16_, connection_1__9__15_, connection_1__9__14_,
         connection_1__9__13_, connection_1__9__12_, connection_1__9__11_,
         connection_1__9__10_, connection_1__9__9_, connection_1__9__8_,
         connection_1__9__7_, connection_1__9__6_, connection_1__9__5_,
         connection_1__9__4_, connection_1__9__3_, connection_1__9__2_,
         connection_1__9__1_, connection_1__9__0_, connection_1__10__31_,
         connection_1__10__30_, connection_1__10__29_, connection_1__10__28_,
         connection_1__10__27_, connection_1__10__26_, connection_1__10__25_,
         connection_1__10__24_, connection_1__10__23_, connection_1__10__22_,
         connection_1__10__21_, connection_1__10__20_, connection_1__10__19_,
         connection_1__10__18_, connection_1__10__17_, connection_1__10__16_,
         connection_1__10__15_, connection_1__10__14_, connection_1__10__13_,
         connection_1__10__12_, connection_1__10__11_, connection_1__10__10_,
         connection_1__10__9_, connection_1__10__8_, connection_1__10__7_,
         connection_1__10__6_, connection_1__10__5_, connection_1__10__4_,
         connection_1__10__3_, connection_1__10__2_, connection_1__10__1_,
         connection_1__10__0_, connection_1__11__31_, connection_1__11__30_,
         connection_1__11__29_, connection_1__11__28_, connection_1__11__27_,
         connection_1__11__26_, connection_1__11__25_, connection_1__11__24_,
         connection_1__11__23_, connection_1__11__22_, connection_1__11__21_,
         connection_1__11__20_, connection_1__11__19_, connection_1__11__18_,
         connection_1__11__17_, connection_1__11__16_, connection_1__11__15_,
         connection_1__11__14_, connection_1__11__13_, connection_1__11__12_,
         connection_1__11__11_, connection_1__11__10_, connection_1__11__9_,
         connection_1__11__8_, connection_1__11__7_, connection_1__11__6_,
         connection_1__11__5_, connection_1__11__4_, connection_1__11__3_,
         connection_1__11__2_, connection_1__11__1_, connection_1__11__0_,
         connection_1__12__31_, connection_1__12__30_, connection_1__12__29_,
         connection_1__12__28_, connection_1__12__27_, connection_1__12__26_,
         connection_1__12__25_, connection_1__12__24_, connection_1__12__23_,
         connection_1__12__22_, connection_1__12__21_, connection_1__12__20_,
         connection_1__12__19_, connection_1__12__18_, connection_1__12__17_,
         connection_1__12__16_, connection_1__12__15_, connection_1__12__14_,
         connection_1__12__13_, connection_1__12__12_, connection_1__12__11_,
         connection_1__12__10_, connection_1__12__9_, connection_1__12__8_,
         connection_1__12__7_, connection_1__12__6_, connection_1__12__5_,
         connection_1__12__4_, connection_1__12__3_, connection_1__12__2_,
         connection_1__12__1_, connection_1__12__0_, connection_1__13__31_,
         connection_1__13__30_, connection_1__13__29_, connection_1__13__28_,
         connection_1__13__27_, connection_1__13__26_, connection_1__13__25_,
         connection_1__13__24_, connection_1__13__23_, connection_1__13__22_,
         connection_1__13__21_, connection_1__13__20_, connection_1__13__19_,
         connection_1__13__18_, connection_1__13__17_, connection_1__13__16_,
         connection_1__13__15_, connection_1__13__14_, connection_1__13__13_,
         connection_1__13__12_, connection_1__13__11_, connection_1__13__10_,
         connection_1__13__9_, connection_1__13__8_, connection_1__13__7_,
         connection_1__13__6_, connection_1__13__5_, connection_1__13__4_,
         connection_1__13__3_, connection_1__13__2_, connection_1__13__1_,
         connection_1__13__0_, connection_1__14__31_, connection_1__14__30_,
         connection_1__14__29_, connection_1__14__28_, connection_1__14__27_,
         connection_1__14__26_, connection_1__14__25_, connection_1__14__24_,
         connection_1__14__23_, connection_1__14__22_, connection_1__14__21_,
         connection_1__14__20_, connection_1__14__19_, connection_1__14__18_,
         connection_1__14__17_, connection_1__14__16_, connection_1__14__15_,
         connection_1__14__14_, connection_1__14__13_, connection_1__14__12_,
         connection_1__14__11_, connection_1__14__10_, connection_1__14__9_,
         connection_1__14__8_, connection_1__14__7_, connection_1__14__6_,
         connection_1__14__5_, connection_1__14__4_, connection_1__14__3_,
         connection_1__14__2_, connection_1__14__1_, connection_1__14__0_,
         connection_1__15__31_, connection_1__15__30_, connection_1__15__29_,
         connection_1__15__28_, connection_1__15__27_, connection_1__15__26_,
         connection_1__15__25_, connection_1__15__24_, connection_1__15__23_,
         connection_1__15__22_, connection_1__15__21_, connection_1__15__20_,
         connection_1__15__19_, connection_1__15__18_, connection_1__15__17_,
         connection_1__15__16_, connection_1__15__15_, connection_1__15__14_,
         connection_1__15__13_, connection_1__15__12_, connection_1__15__11_,
         connection_1__15__10_, connection_1__15__9_, connection_1__15__8_,
         connection_1__15__7_, connection_1__15__6_, connection_1__15__5_,
         connection_1__15__4_, connection_1__15__3_, connection_1__15__2_,
         connection_1__15__1_, connection_1__15__0_, connection_2__0__31_,
         connection_2__0__30_, connection_2__0__29_, connection_2__0__28_,
         connection_2__0__27_, connection_2__0__26_, connection_2__0__25_,
         connection_2__0__24_, connection_2__0__23_, connection_2__0__22_,
         connection_2__0__21_, connection_2__0__20_, connection_2__0__19_,
         connection_2__0__18_, connection_2__0__17_, connection_2__0__16_,
         connection_2__0__15_, connection_2__0__14_, connection_2__0__13_,
         connection_2__0__12_, connection_2__0__11_, connection_2__0__10_,
         connection_2__0__9_, connection_2__0__8_, connection_2__0__7_,
         connection_2__0__6_, connection_2__0__5_, connection_2__0__4_,
         connection_2__0__3_, connection_2__0__2_, connection_2__0__1_,
         connection_2__0__0_, connection_2__1__31_, connection_2__1__30_,
         connection_2__1__29_, connection_2__1__28_, connection_2__1__27_,
         connection_2__1__26_, connection_2__1__25_, connection_2__1__24_,
         connection_2__1__23_, connection_2__1__22_, connection_2__1__21_,
         connection_2__1__20_, connection_2__1__19_, connection_2__1__18_,
         connection_2__1__17_, connection_2__1__16_, connection_2__1__15_,
         connection_2__1__14_, connection_2__1__13_, connection_2__1__12_,
         connection_2__1__11_, connection_2__1__10_, connection_2__1__9_,
         connection_2__1__8_, connection_2__1__7_, connection_2__1__6_,
         connection_2__1__5_, connection_2__1__4_, connection_2__1__3_,
         connection_2__1__2_, connection_2__1__1_, connection_2__1__0_,
         connection_2__2__31_, connection_2__2__30_, connection_2__2__29_,
         connection_2__2__28_, connection_2__2__27_, connection_2__2__26_,
         connection_2__2__25_, connection_2__2__24_, connection_2__2__23_,
         connection_2__2__22_, connection_2__2__21_, connection_2__2__20_,
         connection_2__2__19_, connection_2__2__18_, connection_2__2__17_,
         connection_2__2__16_, connection_2__2__15_, connection_2__2__14_,
         connection_2__2__13_, connection_2__2__12_, connection_2__2__11_,
         connection_2__2__10_, connection_2__2__9_, connection_2__2__8_,
         connection_2__2__7_, connection_2__2__6_, connection_2__2__5_,
         connection_2__2__4_, connection_2__2__3_, connection_2__2__2_,
         connection_2__2__1_, connection_2__2__0_, connection_2__3__31_,
         connection_2__3__30_, connection_2__3__29_, connection_2__3__28_,
         connection_2__3__27_, connection_2__3__26_, connection_2__3__25_,
         connection_2__3__24_, connection_2__3__23_, connection_2__3__22_,
         connection_2__3__21_, connection_2__3__20_, connection_2__3__19_,
         connection_2__3__18_, connection_2__3__17_, connection_2__3__16_,
         connection_2__3__15_, connection_2__3__14_, connection_2__3__13_,
         connection_2__3__12_, connection_2__3__11_, connection_2__3__10_,
         connection_2__3__9_, connection_2__3__8_, connection_2__3__7_,
         connection_2__3__6_, connection_2__3__5_, connection_2__3__4_,
         connection_2__3__3_, connection_2__3__2_, connection_2__3__1_,
         connection_2__3__0_, connection_2__4__31_, connection_2__4__30_,
         connection_2__4__29_, connection_2__4__28_, connection_2__4__27_,
         connection_2__4__26_, connection_2__4__25_, connection_2__4__24_,
         connection_2__4__23_, connection_2__4__22_, connection_2__4__21_,
         connection_2__4__20_, connection_2__4__19_, connection_2__4__18_,
         connection_2__4__17_, connection_2__4__16_, connection_2__4__15_,
         connection_2__4__14_, connection_2__4__13_, connection_2__4__12_,
         connection_2__4__11_, connection_2__4__10_, connection_2__4__9_,
         connection_2__4__8_, connection_2__4__7_, connection_2__4__6_,
         connection_2__4__5_, connection_2__4__4_, connection_2__4__3_,
         connection_2__4__2_, connection_2__4__1_, connection_2__4__0_,
         connection_2__5__31_, connection_2__5__30_, connection_2__5__29_,
         connection_2__5__28_, connection_2__5__27_, connection_2__5__26_,
         connection_2__5__25_, connection_2__5__24_, connection_2__5__23_,
         connection_2__5__22_, connection_2__5__21_, connection_2__5__20_,
         connection_2__5__19_, connection_2__5__18_, connection_2__5__17_,
         connection_2__5__16_, connection_2__5__15_, connection_2__5__14_,
         connection_2__5__13_, connection_2__5__12_, connection_2__5__11_,
         connection_2__5__10_, connection_2__5__9_, connection_2__5__8_,
         connection_2__5__7_, connection_2__5__6_, connection_2__5__5_,
         connection_2__5__4_, connection_2__5__3_, connection_2__5__2_,
         connection_2__5__1_, connection_2__5__0_, connection_2__6__31_,
         connection_2__6__30_, connection_2__6__29_, connection_2__6__28_,
         connection_2__6__27_, connection_2__6__26_, connection_2__6__25_,
         connection_2__6__24_, connection_2__6__23_, connection_2__6__22_,
         connection_2__6__21_, connection_2__6__20_, connection_2__6__19_,
         connection_2__6__18_, connection_2__6__17_, connection_2__6__16_,
         connection_2__6__15_, connection_2__6__14_, connection_2__6__13_,
         connection_2__6__12_, connection_2__6__11_, connection_2__6__10_,
         connection_2__6__9_, connection_2__6__8_, connection_2__6__7_,
         connection_2__6__6_, connection_2__6__5_, connection_2__6__4_,
         connection_2__6__3_, connection_2__6__2_, connection_2__6__1_,
         connection_2__6__0_, connection_2__7__31_, connection_2__7__30_,
         connection_2__7__29_, connection_2__7__28_, connection_2__7__27_,
         connection_2__7__26_, connection_2__7__25_, connection_2__7__24_,
         connection_2__7__23_, connection_2__7__22_, connection_2__7__21_,
         connection_2__7__20_, connection_2__7__19_, connection_2__7__18_,
         connection_2__7__17_, connection_2__7__16_, connection_2__7__15_,
         connection_2__7__14_, connection_2__7__13_, connection_2__7__12_,
         connection_2__7__11_, connection_2__7__10_, connection_2__7__9_,
         connection_2__7__8_, connection_2__7__7_, connection_2__7__6_,
         connection_2__7__5_, connection_2__7__4_, connection_2__7__3_,
         connection_2__7__2_, connection_2__7__1_, connection_2__7__0_,
         connection_2__8__31_, connection_2__8__30_, connection_2__8__29_,
         connection_2__8__28_, connection_2__8__27_, connection_2__8__26_,
         connection_2__8__25_, connection_2__8__24_, connection_2__8__23_,
         connection_2__8__22_, connection_2__8__21_, connection_2__8__20_,
         connection_2__8__19_, connection_2__8__18_, connection_2__8__17_,
         connection_2__8__16_, connection_2__8__15_, connection_2__8__14_,
         connection_2__8__13_, connection_2__8__12_, connection_2__8__11_,
         connection_2__8__10_, connection_2__8__9_, connection_2__8__8_,
         connection_2__8__7_, connection_2__8__6_, connection_2__8__5_,
         connection_2__8__4_, connection_2__8__3_, connection_2__8__2_,
         connection_2__8__1_, connection_2__8__0_, connection_2__9__31_,
         connection_2__9__30_, connection_2__9__29_, connection_2__9__28_,
         connection_2__9__27_, connection_2__9__26_, connection_2__9__25_,
         connection_2__9__24_, connection_2__9__23_, connection_2__9__22_,
         connection_2__9__21_, connection_2__9__20_, connection_2__9__19_,
         connection_2__9__18_, connection_2__9__17_, connection_2__9__16_,
         connection_2__9__15_, connection_2__9__14_, connection_2__9__13_,
         connection_2__9__12_, connection_2__9__11_, connection_2__9__10_,
         connection_2__9__9_, connection_2__9__8_, connection_2__9__7_,
         connection_2__9__6_, connection_2__9__5_, connection_2__9__4_,
         connection_2__9__3_, connection_2__9__2_, connection_2__9__1_,
         connection_2__9__0_, connection_2__10__31_, connection_2__10__30_,
         connection_2__10__29_, connection_2__10__28_, connection_2__10__27_,
         connection_2__10__26_, connection_2__10__25_, connection_2__10__24_,
         connection_2__10__23_, connection_2__10__22_, connection_2__10__21_,
         connection_2__10__20_, connection_2__10__19_, connection_2__10__18_,
         connection_2__10__17_, connection_2__10__16_, connection_2__10__15_,
         connection_2__10__14_, connection_2__10__13_, connection_2__10__12_,
         connection_2__10__11_, connection_2__10__10_, connection_2__10__9_,
         connection_2__10__8_, connection_2__10__7_, connection_2__10__6_,
         connection_2__10__5_, connection_2__10__4_, connection_2__10__3_,
         connection_2__10__2_, connection_2__10__1_, connection_2__10__0_,
         connection_2__11__31_, connection_2__11__30_, connection_2__11__29_,
         connection_2__11__28_, connection_2__11__27_, connection_2__11__26_,
         connection_2__11__25_, connection_2__11__24_, connection_2__11__23_,
         connection_2__11__22_, connection_2__11__21_, connection_2__11__20_,
         connection_2__11__19_, connection_2__11__18_, connection_2__11__17_,
         connection_2__11__16_, connection_2__11__15_, connection_2__11__14_,
         connection_2__11__13_, connection_2__11__12_, connection_2__11__11_,
         connection_2__11__10_, connection_2__11__9_, connection_2__11__8_,
         connection_2__11__7_, connection_2__11__6_, connection_2__11__5_,
         connection_2__11__4_, connection_2__11__3_, connection_2__11__2_,
         connection_2__11__1_, connection_2__11__0_, connection_2__12__31_,
         connection_2__12__30_, connection_2__12__29_, connection_2__12__28_,
         connection_2__12__27_, connection_2__12__26_, connection_2__12__25_,
         connection_2__12__24_, connection_2__12__23_, connection_2__12__22_,
         connection_2__12__21_, connection_2__12__20_, connection_2__12__19_,
         connection_2__12__18_, connection_2__12__17_, connection_2__12__16_,
         connection_2__12__15_, connection_2__12__14_, connection_2__12__13_,
         connection_2__12__12_, connection_2__12__11_, connection_2__12__10_,
         connection_2__12__9_, connection_2__12__8_, connection_2__12__7_,
         connection_2__12__6_, connection_2__12__5_, connection_2__12__4_,
         connection_2__12__3_, connection_2__12__2_, connection_2__12__1_,
         connection_2__12__0_, connection_2__13__31_, connection_2__13__30_,
         connection_2__13__29_, connection_2__13__28_, connection_2__13__27_,
         connection_2__13__26_, connection_2__13__25_, connection_2__13__24_,
         connection_2__13__23_, connection_2__13__22_, connection_2__13__21_,
         connection_2__13__20_, connection_2__13__19_, connection_2__13__18_,
         connection_2__13__17_, connection_2__13__16_, connection_2__13__15_,
         connection_2__13__14_, connection_2__13__13_, connection_2__13__12_,
         connection_2__13__11_, connection_2__13__10_, connection_2__13__9_,
         connection_2__13__8_, connection_2__13__7_, connection_2__13__6_,
         connection_2__13__5_, connection_2__13__4_, connection_2__13__3_,
         connection_2__13__2_, connection_2__13__1_, connection_2__13__0_,
         connection_2__14__31_, connection_2__14__30_, connection_2__14__29_,
         connection_2__14__28_, connection_2__14__27_, connection_2__14__26_,
         connection_2__14__25_, connection_2__14__24_, connection_2__14__23_,
         connection_2__14__22_, connection_2__14__21_, connection_2__14__20_,
         connection_2__14__19_, connection_2__14__18_, connection_2__14__17_,
         connection_2__14__16_, connection_2__14__15_, connection_2__14__14_,
         connection_2__14__13_, connection_2__14__12_, connection_2__14__11_,
         connection_2__14__10_, connection_2__14__9_, connection_2__14__8_,
         connection_2__14__7_, connection_2__14__6_, connection_2__14__5_,
         connection_2__14__4_, connection_2__14__3_, connection_2__14__2_,
         connection_2__14__1_, connection_2__14__0_, connection_2__15__31_,
         connection_2__15__30_, connection_2__15__29_, connection_2__15__28_,
         connection_2__15__27_, connection_2__15__26_, connection_2__15__25_,
         connection_2__15__24_, connection_2__15__23_, connection_2__15__22_,
         connection_2__15__21_, connection_2__15__20_, connection_2__15__19_,
         connection_2__15__18_, connection_2__15__17_, connection_2__15__16_,
         connection_2__15__15_, connection_2__15__14_, connection_2__15__13_,
         connection_2__15__12_, connection_2__15__11_, connection_2__15__10_,
         connection_2__15__9_, connection_2__15__8_, connection_2__15__7_,
         connection_2__15__6_, connection_2__15__5_, connection_2__15__4_,
         connection_2__15__3_, connection_2__15__2_, connection_2__15__1_,
         connection_2__15__0_, connection_3__0__31_, connection_3__0__30_,
         connection_3__0__29_, connection_3__0__28_, connection_3__0__27_,
         connection_3__0__26_, connection_3__0__25_, connection_3__0__24_,
         connection_3__0__23_, connection_3__0__22_, connection_3__0__21_,
         connection_3__0__20_, connection_3__0__19_, connection_3__0__18_,
         connection_3__0__17_, connection_3__0__16_, connection_3__0__15_,
         connection_3__0__14_, connection_3__0__13_, connection_3__0__12_,
         connection_3__0__11_, connection_3__0__10_, connection_3__0__9_,
         connection_3__0__8_, connection_3__0__7_, connection_3__0__6_,
         connection_3__0__5_, connection_3__0__4_, connection_3__0__3_,
         connection_3__0__2_, connection_3__0__1_, connection_3__0__0_,
         connection_3__1__31_, connection_3__1__30_, connection_3__1__29_,
         connection_3__1__28_, connection_3__1__27_, connection_3__1__26_,
         connection_3__1__25_, connection_3__1__24_, connection_3__1__23_,
         connection_3__1__22_, connection_3__1__21_, connection_3__1__20_,
         connection_3__1__19_, connection_3__1__18_, connection_3__1__17_,
         connection_3__1__16_, connection_3__1__15_, connection_3__1__14_,
         connection_3__1__13_, connection_3__1__12_, connection_3__1__11_,
         connection_3__1__10_, connection_3__1__9_, connection_3__1__8_,
         connection_3__1__7_, connection_3__1__6_, connection_3__1__5_,
         connection_3__1__4_, connection_3__1__3_, connection_3__1__2_,
         connection_3__1__1_, connection_3__1__0_, connection_3__2__31_,
         connection_3__2__30_, connection_3__2__29_, connection_3__2__28_,
         connection_3__2__27_, connection_3__2__26_, connection_3__2__25_,
         connection_3__2__24_, connection_3__2__23_, connection_3__2__22_,
         connection_3__2__21_, connection_3__2__20_, connection_3__2__19_,
         connection_3__2__18_, connection_3__2__17_, connection_3__2__16_,
         connection_3__2__15_, connection_3__2__14_, connection_3__2__13_,
         connection_3__2__12_, connection_3__2__11_, connection_3__2__10_,
         connection_3__2__9_, connection_3__2__8_, connection_3__2__7_,
         connection_3__2__6_, connection_3__2__5_, connection_3__2__4_,
         connection_3__2__3_, connection_3__2__2_, connection_3__2__1_,
         connection_3__2__0_, connection_3__3__31_, connection_3__3__30_,
         connection_3__3__29_, connection_3__3__28_, connection_3__3__27_,
         connection_3__3__26_, connection_3__3__25_, connection_3__3__24_,
         connection_3__3__23_, connection_3__3__22_, connection_3__3__21_,
         connection_3__3__20_, connection_3__3__19_, connection_3__3__18_,
         connection_3__3__17_, connection_3__3__16_, connection_3__3__15_,
         connection_3__3__14_, connection_3__3__13_, connection_3__3__12_,
         connection_3__3__11_, connection_3__3__10_, connection_3__3__9_,
         connection_3__3__8_, connection_3__3__7_, connection_3__3__6_,
         connection_3__3__5_, connection_3__3__4_, connection_3__3__3_,
         connection_3__3__2_, connection_3__3__1_, connection_3__3__0_,
         connection_3__4__31_, connection_3__4__30_, connection_3__4__29_,
         connection_3__4__28_, connection_3__4__27_, connection_3__4__26_,
         connection_3__4__25_, connection_3__4__24_, connection_3__4__23_,
         connection_3__4__22_, connection_3__4__21_, connection_3__4__20_,
         connection_3__4__19_, connection_3__4__18_, connection_3__4__17_,
         connection_3__4__16_, connection_3__4__15_, connection_3__4__14_,
         connection_3__4__13_, connection_3__4__12_, connection_3__4__11_,
         connection_3__4__10_, connection_3__4__9_, connection_3__4__8_,
         connection_3__4__7_, connection_3__4__6_, connection_3__4__5_,
         connection_3__4__4_, connection_3__4__3_, connection_3__4__2_,
         connection_3__4__1_, connection_3__4__0_, connection_3__5__31_,
         connection_3__5__30_, connection_3__5__29_, connection_3__5__28_,
         connection_3__5__27_, connection_3__5__26_, connection_3__5__25_,
         connection_3__5__24_, connection_3__5__23_, connection_3__5__22_,
         connection_3__5__21_, connection_3__5__20_, connection_3__5__19_,
         connection_3__5__18_, connection_3__5__17_, connection_3__5__16_,
         connection_3__5__15_, connection_3__5__14_, connection_3__5__13_,
         connection_3__5__12_, connection_3__5__11_, connection_3__5__10_,
         connection_3__5__9_, connection_3__5__8_, connection_3__5__7_,
         connection_3__5__6_, connection_3__5__5_, connection_3__5__4_,
         connection_3__5__3_, connection_3__5__2_, connection_3__5__1_,
         connection_3__5__0_, connection_3__6__31_, connection_3__6__30_,
         connection_3__6__29_, connection_3__6__28_, connection_3__6__27_,
         connection_3__6__26_, connection_3__6__25_, connection_3__6__24_,
         connection_3__6__23_, connection_3__6__22_, connection_3__6__21_,
         connection_3__6__20_, connection_3__6__19_, connection_3__6__18_,
         connection_3__6__17_, connection_3__6__16_, connection_3__6__15_,
         connection_3__6__14_, connection_3__6__13_, connection_3__6__12_,
         connection_3__6__11_, connection_3__6__10_, connection_3__6__9_,
         connection_3__6__8_, connection_3__6__7_, connection_3__6__6_,
         connection_3__6__5_, connection_3__6__4_, connection_3__6__3_,
         connection_3__6__2_, connection_3__6__1_, connection_3__6__0_,
         connection_3__7__31_, connection_3__7__30_, connection_3__7__29_,
         connection_3__7__28_, connection_3__7__27_, connection_3__7__26_,
         connection_3__7__25_, connection_3__7__24_, connection_3__7__23_,
         connection_3__7__22_, connection_3__7__21_, connection_3__7__20_,
         connection_3__7__19_, connection_3__7__18_, connection_3__7__17_,
         connection_3__7__16_, connection_3__7__15_, connection_3__7__14_,
         connection_3__7__13_, connection_3__7__12_, connection_3__7__11_,
         connection_3__7__10_, connection_3__7__9_, connection_3__7__8_,
         connection_3__7__7_, connection_3__7__6_, connection_3__7__5_,
         connection_3__7__4_, connection_3__7__3_, connection_3__7__2_,
         connection_3__7__1_, connection_3__7__0_, connection_3__8__31_,
         connection_3__8__30_, connection_3__8__29_, connection_3__8__28_,
         connection_3__8__27_, connection_3__8__26_, connection_3__8__25_,
         connection_3__8__24_, connection_3__8__23_, connection_3__8__22_,
         connection_3__8__21_, connection_3__8__20_, connection_3__8__19_,
         connection_3__8__18_, connection_3__8__17_, connection_3__8__16_,
         connection_3__8__15_, connection_3__8__14_, connection_3__8__13_,
         connection_3__8__12_, connection_3__8__11_, connection_3__8__10_,
         connection_3__8__9_, connection_3__8__8_, connection_3__8__7_,
         connection_3__8__6_, connection_3__8__5_, connection_3__8__4_,
         connection_3__8__3_, connection_3__8__2_, connection_3__8__1_,
         connection_3__8__0_, connection_3__9__31_, connection_3__9__30_,
         connection_3__9__29_, connection_3__9__28_, connection_3__9__27_,
         connection_3__9__26_, connection_3__9__25_, connection_3__9__24_,
         connection_3__9__23_, connection_3__9__22_, connection_3__9__21_,
         connection_3__9__20_, connection_3__9__19_, connection_3__9__18_,
         connection_3__9__17_, connection_3__9__16_, connection_3__9__15_,
         connection_3__9__14_, connection_3__9__13_, connection_3__9__12_,
         connection_3__9__11_, connection_3__9__10_, connection_3__9__9_,
         connection_3__9__8_, connection_3__9__7_, connection_3__9__6_,
         connection_3__9__5_, connection_3__9__4_, connection_3__9__3_,
         connection_3__9__2_, connection_3__9__1_, connection_3__9__0_,
         connection_3__10__31_, connection_3__10__30_, connection_3__10__29_,
         connection_3__10__28_, connection_3__10__27_, connection_3__10__26_,
         connection_3__10__25_, connection_3__10__24_, connection_3__10__23_,
         connection_3__10__22_, connection_3__10__21_, connection_3__10__20_,
         connection_3__10__19_, connection_3__10__18_, connection_3__10__17_,
         connection_3__10__16_, connection_3__10__15_, connection_3__10__14_,
         connection_3__10__13_, connection_3__10__12_, connection_3__10__11_,
         connection_3__10__10_, connection_3__10__9_, connection_3__10__8_,
         connection_3__10__7_, connection_3__10__6_, connection_3__10__5_,
         connection_3__10__4_, connection_3__10__3_, connection_3__10__2_,
         connection_3__10__1_, connection_3__10__0_, connection_3__11__31_,
         connection_3__11__30_, connection_3__11__29_, connection_3__11__28_,
         connection_3__11__27_, connection_3__11__26_, connection_3__11__25_,
         connection_3__11__24_, connection_3__11__23_, connection_3__11__22_,
         connection_3__11__21_, connection_3__11__20_, connection_3__11__19_,
         connection_3__11__18_, connection_3__11__17_, connection_3__11__16_,
         connection_3__11__15_, connection_3__11__14_, connection_3__11__13_,
         connection_3__11__12_, connection_3__11__11_, connection_3__11__10_,
         connection_3__11__9_, connection_3__11__8_, connection_3__11__7_,
         connection_3__11__6_, connection_3__11__5_, connection_3__11__4_,
         connection_3__11__3_, connection_3__11__2_, connection_3__11__1_,
         connection_3__11__0_, connection_3__12__31_, connection_3__12__30_,
         connection_3__12__29_, connection_3__12__28_, connection_3__12__27_,
         connection_3__12__26_, connection_3__12__25_, connection_3__12__24_,
         connection_3__12__23_, connection_3__12__22_, connection_3__12__21_,
         connection_3__12__20_, connection_3__12__19_, connection_3__12__18_,
         connection_3__12__17_, connection_3__12__16_, connection_3__12__15_,
         connection_3__12__14_, connection_3__12__13_, connection_3__12__12_,
         connection_3__12__11_, connection_3__12__10_, connection_3__12__9_,
         connection_3__12__8_, connection_3__12__7_, connection_3__12__6_,
         connection_3__12__5_, connection_3__12__4_, connection_3__12__3_,
         connection_3__12__2_, connection_3__12__1_, connection_3__12__0_,
         connection_3__13__31_, connection_3__13__30_, connection_3__13__29_,
         connection_3__13__28_, connection_3__13__27_, connection_3__13__26_,
         connection_3__13__25_, connection_3__13__24_, connection_3__13__23_,
         connection_3__13__22_, connection_3__13__21_, connection_3__13__20_,
         connection_3__13__19_, connection_3__13__18_, connection_3__13__17_,
         connection_3__13__16_, connection_3__13__15_, connection_3__13__14_,
         connection_3__13__13_, connection_3__13__12_, connection_3__13__11_,
         connection_3__13__10_, connection_3__13__9_, connection_3__13__8_,
         connection_3__13__7_, connection_3__13__6_, connection_3__13__5_,
         connection_3__13__4_, connection_3__13__3_, connection_3__13__2_,
         connection_3__13__1_, connection_3__13__0_, connection_3__14__31_,
         connection_3__14__30_, connection_3__14__29_, connection_3__14__28_,
         connection_3__14__27_, connection_3__14__26_, connection_3__14__25_,
         connection_3__14__24_, connection_3__14__23_, connection_3__14__22_,
         connection_3__14__21_, connection_3__14__20_, connection_3__14__19_,
         connection_3__14__18_, connection_3__14__17_, connection_3__14__16_,
         connection_3__14__15_, connection_3__14__14_, connection_3__14__13_,
         connection_3__14__12_, connection_3__14__11_, connection_3__14__10_,
         connection_3__14__9_, connection_3__14__8_, connection_3__14__7_,
         connection_3__14__6_, connection_3__14__5_, connection_3__14__4_,
         connection_3__14__3_, connection_3__14__2_, connection_3__14__1_,
         connection_3__14__0_, connection_3__15__31_, connection_3__15__30_,
         connection_3__15__29_, connection_3__15__28_, connection_3__15__27_,
         connection_3__15__26_, connection_3__15__25_, connection_3__15__24_,
         connection_3__15__23_, connection_3__15__22_, connection_3__15__21_,
         connection_3__15__20_, connection_3__15__19_, connection_3__15__18_,
         connection_3__15__17_, connection_3__15__16_, connection_3__15__15_,
         connection_3__15__14_, connection_3__15__13_, connection_3__15__12_,
         connection_3__15__11_, connection_3__15__10_, connection_3__15__9_,
         connection_3__15__8_, connection_3__15__7_, connection_3__15__6_,
         connection_3__15__5_, connection_3__15__4_, connection_3__15__3_,
         connection_3__15__2_, connection_3__15__1_, connection_3__15__0_,
         connection_4__0__31_, connection_4__0__30_, connection_4__0__29_,
         connection_4__0__28_, connection_4__0__27_, connection_4__0__26_,
         connection_4__0__25_, connection_4__0__24_, connection_4__0__23_,
         connection_4__0__22_, connection_4__0__21_, connection_4__0__20_,
         connection_4__0__19_, connection_4__0__18_, connection_4__0__17_,
         connection_4__0__16_, connection_4__0__15_, connection_4__0__14_,
         connection_4__0__13_, connection_4__0__12_, connection_4__0__11_,
         connection_4__0__10_, connection_4__0__9_, connection_4__0__8_,
         connection_4__0__7_, connection_4__0__6_, connection_4__0__5_,
         connection_4__0__4_, connection_4__0__3_, connection_4__0__2_,
         connection_4__0__1_, connection_4__0__0_, connection_4__1__31_,
         connection_4__1__30_, connection_4__1__29_, connection_4__1__28_,
         connection_4__1__27_, connection_4__1__26_, connection_4__1__25_,
         connection_4__1__24_, connection_4__1__23_, connection_4__1__22_,
         connection_4__1__21_, connection_4__1__20_, connection_4__1__19_,
         connection_4__1__18_, connection_4__1__17_, connection_4__1__16_,
         connection_4__1__15_, connection_4__1__14_, connection_4__1__13_,
         connection_4__1__12_, connection_4__1__11_, connection_4__1__10_,
         connection_4__1__9_, connection_4__1__8_, connection_4__1__7_,
         connection_4__1__6_, connection_4__1__5_, connection_4__1__4_,
         connection_4__1__3_, connection_4__1__2_, connection_4__1__1_,
         connection_4__1__0_, connection_4__2__31_, connection_4__2__30_,
         connection_4__2__29_, connection_4__2__28_, connection_4__2__27_,
         connection_4__2__26_, connection_4__2__25_, connection_4__2__24_,
         connection_4__2__23_, connection_4__2__22_, connection_4__2__21_,
         connection_4__2__20_, connection_4__2__19_, connection_4__2__18_,
         connection_4__2__17_, connection_4__2__16_, connection_4__2__15_,
         connection_4__2__14_, connection_4__2__13_, connection_4__2__12_,
         connection_4__2__11_, connection_4__2__10_, connection_4__2__9_,
         connection_4__2__8_, connection_4__2__7_, connection_4__2__6_,
         connection_4__2__5_, connection_4__2__4_, connection_4__2__3_,
         connection_4__2__2_, connection_4__2__1_, connection_4__2__0_,
         connection_4__3__31_, connection_4__3__30_, connection_4__3__29_,
         connection_4__3__28_, connection_4__3__27_, connection_4__3__26_,
         connection_4__3__25_, connection_4__3__24_, connection_4__3__23_,
         connection_4__3__22_, connection_4__3__21_, connection_4__3__20_,
         connection_4__3__19_, connection_4__3__18_, connection_4__3__17_,
         connection_4__3__16_, connection_4__3__15_, connection_4__3__14_,
         connection_4__3__13_, connection_4__3__12_, connection_4__3__11_,
         connection_4__3__10_, connection_4__3__9_, connection_4__3__8_,
         connection_4__3__7_, connection_4__3__6_, connection_4__3__5_,
         connection_4__3__4_, connection_4__3__3_, connection_4__3__2_,
         connection_4__3__1_, connection_4__3__0_, connection_4__4__31_,
         connection_4__4__30_, connection_4__4__29_, connection_4__4__28_,
         connection_4__4__27_, connection_4__4__26_, connection_4__4__25_,
         connection_4__4__24_, connection_4__4__23_, connection_4__4__22_,
         connection_4__4__21_, connection_4__4__20_, connection_4__4__19_,
         connection_4__4__18_, connection_4__4__17_, connection_4__4__16_,
         connection_4__4__15_, connection_4__4__14_, connection_4__4__13_,
         connection_4__4__12_, connection_4__4__11_, connection_4__4__10_,
         connection_4__4__9_, connection_4__4__8_, connection_4__4__7_,
         connection_4__4__6_, connection_4__4__5_, connection_4__4__4_,
         connection_4__4__3_, connection_4__4__2_, connection_4__4__1_,
         connection_4__4__0_, connection_4__5__31_, connection_4__5__30_,
         connection_4__5__29_, connection_4__5__28_, connection_4__5__27_,
         connection_4__5__26_, connection_4__5__25_, connection_4__5__24_,
         connection_4__5__23_, connection_4__5__22_, connection_4__5__21_,
         connection_4__5__20_, connection_4__5__19_, connection_4__5__18_,
         connection_4__5__17_, connection_4__5__16_, connection_4__5__15_,
         connection_4__5__14_, connection_4__5__13_, connection_4__5__12_,
         connection_4__5__11_, connection_4__5__10_, connection_4__5__9_,
         connection_4__5__8_, connection_4__5__7_, connection_4__5__6_,
         connection_4__5__5_, connection_4__5__4_, connection_4__5__3_,
         connection_4__5__2_, connection_4__5__1_, connection_4__5__0_,
         connection_4__6__31_, connection_4__6__30_, connection_4__6__29_,
         connection_4__6__28_, connection_4__6__27_, connection_4__6__26_,
         connection_4__6__25_, connection_4__6__24_, connection_4__6__23_,
         connection_4__6__22_, connection_4__6__21_, connection_4__6__20_,
         connection_4__6__19_, connection_4__6__18_, connection_4__6__17_,
         connection_4__6__16_, connection_4__6__15_, connection_4__6__14_,
         connection_4__6__13_, connection_4__6__12_, connection_4__6__11_,
         connection_4__6__10_, connection_4__6__9_, connection_4__6__8_,
         connection_4__6__7_, connection_4__6__6_, connection_4__6__5_,
         connection_4__6__4_, connection_4__6__3_, connection_4__6__2_,
         connection_4__6__1_, connection_4__6__0_, connection_4__7__31_,
         connection_4__7__30_, connection_4__7__29_, connection_4__7__28_,
         connection_4__7__27_, connection_4__7__26_, connection_4__7__25_,
         connection_4__7__24_, connection_4__7__23_, connection_4__7__22_,
         connection_4__7__21_, connection_4__7__20_, connection_4__7__19_,
         connection_4__7__18_, connection_4__7__17_, connection_4__7__16_,
         connection_4__7__15_, connection_4__7__14_, connection_4__7__13_,
         connection_4__7__12_, connection_4__7__11_, connection_4__7__10_,
         connection_4__7__9_, connection_4__7__8_, connection_4__7__7_,
         connection_4__7__6_, connection_4__7__5_, connection_4__7__4_,
         connection_4__7__3_, connection_4__7__2_, connection_4__7__1_,
         connection_4__7__0_, connection_4__8__31_, connection_4__8__30_,
         connection_4__8__29_, connection_4__8__28_, connection_4__8__27_,
         connection_4__8__26_, connection_4__8__25_, connection_4__8__24_,
         connection_4__8__23_, connection_4__8__22_, connection_4__8__21_,
         connection_4__8__20_, connection_4__8__19_, connection_4__8__18_,
         connection_4__8__17_, connection_4__8__16_, connection_4__8__15_,
         connection_4__8__14_, connection_4__8__13_, connection_4__8__12_,
         connection_4__8__11_, connection_4__8__10_, connection_4__8__9_,
         connection_4__8__8_, connection_4__8__7_, connection_4__8__6_,
         connection_4__8__5_, connection_4__8__4_, connection_4__8__3_,
         connection_4__8__2_, connection_4__8__1_, connection_4__8__0_,
         connection_4__9__31_, connection_4__9__30_, connection_4__9__29_,
         connection_4__9__28_, connection_4__9__27_, connection_4__9__26_,
         connection_4__9__25_, connection_4__9__24_, connection_4__9__23_,
         connection_4__9__22_, connection_4__9__21_, connection_4__9__20_,
         connection_4__9__19_, connection_4__9__18_, connection_4__9__17_,
         connection_4__9__16_, connection_4__9__15_, connection_4__9__14_,
         connection_4__9__13_, connection_4__9__12_, connection_4__9__11_,
         connection_4__9__10_, connection_4__9__9_, connection_4__9__8_,
         connection_4__9__7_, connection_4__9__6_, connection_4__9__5_,
         connection_4__9__4_, connection_4__9__3_, connection_4__9__2_,
         connection_4__9__1_, connection_4__9__0_, connection_4__10__31_,
         connection_4__10__30_, connection_4__10__29_, connection_4__10__28_,
         connection_4__10__27_, connection_4__10__26_, connection_4__10__25_,
         connection_4__10__24_, connection_4__10__23_, connection_4__10__22_,
         connection_4__10__21_, connection_4__10__20_, connection_4__10__19_,
         connection_4__10__18_, connection_4__10__17_, connection_4__10__16_,
         connection_4__10__15_, connection_4__10__14_, connection_4__10__13_,
         connection_4__10__12_, connection_4__10__11_, connection_4__10__10_,
         connection_4__10__9_, connection_4__10__8_, connection_4__10__7_,
         connection_4__10__6_, connection_4__10__5_, connection_4__10__4_,
         connection_4__10__3_, connection_4__10__2_, connection_4__10__1_,
         connection_4__10__0_, connection_4__11__31_, connection_4__11__30_,
         connection_4__11__29_, connection_4__11__28_, connection_4__11__27_,
         connection_4__11__26_, connection_4__11__25_, connection_4__11__24_,
         connection_4__11__23_, connection_4__11__22_, connection_4__11__21_,
         connection_4__11__20_, connection_4__11__19_, connection_4__11__18_,
         connection_4__11__17_, connection_4__11__16_, connection_4__11__15_,
         connection_4__11__14_, connection_4__11__13_, connection_4__11__12_,
         connection_4__11__11_, connection_4__11__10_, connection_4__11__9_,
         connection_4__11__8_, connection_4__11__7_, connection_4__11__6_,
         connection_4__11__5_, connection_4__11__4_, connection_4__11__3_,
         connection_4__11__2_, connection_4__11__1_, connection_4__11__0_,
         connection_4__12__31_, connection_4__12__30_, connection_4__12__29_,
         connection_4__12__28_, connection_4__12__27_, connection_4__12__26_,
         connection_4__12__25_, connection_4__12__24_, connection_4__12__23_,
         connection_4__12__22_, connection_4__12__21_, connection_4__12__20_,
         connection_4__12__19_, connection_4__12__18_, connection_4__12__17_,
         connection_4__12__16_, connection_4__12__15_, connection_4__12__14_,
         connection_4__12__13_, connection_4__12__12_, connection_4__12__11_,
         connection_4__12__10_, connection_4__12__9_, connection_4__12__8_,
         connection_4__12__7_, connection_4__12__6_, connection_4__12__5_,
         connection_4__12__4_, connection_4__12__3_, connection_4__12__2_,
         connection_4__12__1_, connection_4__12__0_, connection_4__13__31_,
         connection_4__13__30_, connection_4__13__29_, connection_4__13__28_,
         connection_4__13__27_, connection_4__13__26_, connection_4__13__25_,
         connection_4__13__24_, connection_4__13__23_, connection_4__13__22_,
         connection_4__13__21_, connection_4__13__20_, connection_4__13__19_,
         connection_4__13__18_, connection_4__13__17_, connection_4__13__16_,
         connection_4__13__15_, connection_4__13__14_, connection_4__13__13_,
         connection_4__13__12_, connection_4__13__11_, connection_4__13__10_,
         connection_4__13__9_, connection_4__13__8_, connection_4__13__7_,
         connection_4__13__6_, connection_4__13__5_, connection_4__13__4_,
         connection_4__13__3_, connection_4__13__2_, connection_4__13__1_,
         connection_4__13__0_, connection_4__14__31_, connection_4__14__30_,
         connection_4__14__29_, connection_4__14__28_, connection_4__14__27_,
         connection_4__14__26_, connection_4__14__25_, connection_4__14__24_,
         connection_4__14__23_, connection_4__14__22_, connection_4__14__21_,
         connection_4__14__20_, connection_4__14__19_, connection_4__14__18_,
         connection_4__14__17_, connection_4__14__16_, connection_4__14__15_,
         connection_4__14__14_, connection_4__14__13_, connection_4__14__12_,
         connection_4__14__11_, connection_4__14__10_, connection_4__14__9_,
         connection_4__14__8_, connection_4__14__7_, connection_4__14__6_,
         connection_4__14__5_, connection_4__14__4_, connection_4__14__3_,
         connection_4__14__2_, connection_4__14__1_, connection_4__14__0_,
         connection_4__15__31_, connection_4__15__30_, connection_4__15__29_,
         connection_4__15__28_, connection_4__15__27_, connection_4__15__26_,
         connection_4__15__25_, connection_4__15__24_, connection_4__15__23_,
         connection_4__15__22_, connection_4__15__21_, connection_4__15__20_,
         connection_4__15__19_, connection_4__15__18_, connection_4__15__17_,
         connection_4__15__16_, connection_4__15__15_, connection_4__15__14_,
         connection_4__15__13_, connection_4__15__12_, connection_4__15__11_,
         connection_4__15__10_, connection_4__15__9_, connection_4__15__8_,
         connection_4__15__7_, connection_4__15__6_, connection_4__15__5_,
         connection_4__15__4_, connection_4__15__3_, connection_4__15__2_,
         connection_4__15__1_, connection_4__15__0_, connection_5__0__31_,
         connection_5__0__30_, connection_5__0__29_, connection_5__0__28_,
         connection_5__0__27_, connection_5__0__26_, connection_5__0__25_,
         connection_5__0__24_, connection_5__0__23_, connection_5__0__22_,
         connection_5__0__21_, connection_5__0__20_, connection_5__0__19_,
         connection_5__0__18_, connection_5__0__17_, connection_5__0__16_,
         connection_5__0__15_, connection_5__0__14_, connection_5__0__13_,
         connection_5__0__12_, connection_5__0__11_, connection_5__0__10_,
         connection_5__0__9_, connection_5__0__8_, connection_5__0__7_,
         connection_5__0__6_, connection_5__0__5_, connection_5__0__4_,
         connection_5__0__3_, connection_5__0__2_, connection_5__0__1_,
         connection_5__0__0_, connection_5__1__31_, connection_5__1__30_,
         connection_5__1__29_, connection_5__1__28_, connection_5__1__27_,
         connection_5__1__26_, connection_5__1__25_, connection_5__1__24_,
         connection_5__1__23_, connection_5__1__22_, connection_5__1__21_,
         connection_5__1__20_, connection_5__1__19_, connection_5__1__18_,
         connection_5__1__17_, connection_5__1__16_, connection_5__1__15_,
         connection_5__1__14_, connection_5__1__13_, connection_5__1__12_,
         connection_5__1__11_, connection_5__1__10_, connection_5__1__9_,
         connection_5__1__8_, connection_5__1__7_, connection_5__1__6_,
         connection_5__1__5_, connection_5__1__4_, connection_5__1__3_,
         connection_5__1__2_, connection_5__1__1_, connection_5__1__0_,
         connection_5__2__31_, connection_5__2__30_, connection_5__2__29_,
         connection_5__2__28_, connection_5__2__27_, connection_5__2__26_,
         connection_5__2__25_, connection_5__2__24_, connection_5__2__23_,
         connection_5__2__22_, connection_5__2__21_, connection_5__2__20_,
         connection_5__2__19_, connection_5__2__18_, connection_5__2__17_,
         connection_5__2__16_, connection_5__2__15_, connection_5__2__14_,
         connection_5__2__13_, connection_5__2__12_, connection_5__2__11_,
         connection_5__2__10_, connection_5__2__9_, connection_5__2__8_,
         connection_5__2__7_, connection_5__2__6_, connection_5__2__5_,
         connection_5__2__4_, connection_5__2__3_, connection_5__2__2_,
         connection_5__2__1_, connection_5__2__0_, connection_5__3__31_,
         connection_5__3__30_, connection_5__3__29_, connection_5__3__28_,
         connection_5__3__27_, connection_5__3__26_, connection_5__3__25_,
         connection_5__3__24_, connection_5__3__23_, connection_5__3__22_,
         connection_5__3__21_, connection_5__3__20_, connection_5__3__19_,
         connection_5__3__18_, connection_5__3__17_, connection_5__3__16_,
         connection_5__3__15_, connection_5__3__14_, connection_5__3__13_,
         connection_5__3__12_, connection_5__3__11_, connection_5__3__10_,
         connection_5__3__9_, connection_5__3__8_, connection_5__3__7_,
         connection_5__3__6_, connection_5__3__5_, connection_5__3__4_,
         connection_5__3__3_, connection_5__3__2_, connection_5__3__1_,
         connection_5__3__0_, connection_5__4__31_, connection_5__4__30_,
         connection_5__4__29_, connection_5__4__28_, connection_5__4__27_,
         connection_5__4__26_, connection_5__4__25_, connection_5__4__24_,
         connection_5__4__23_, connection_5__4__22_, connection_5__4__21_,
         connection_5__4__20_, connection_5__4__19_, connection_5__4__18_,
         connection_5__4__17_, connection_5__4__16_, connection_5__4__15_,
         connection_5__4__14_, connection_5__4__13_, connection_5__4__12_,
         connection_5__4__11_, connection_5__4__10_, connection_5__4__9_,
         connection_5__4__8_, connection_5__4__7_, connection_5__4__6_,
         connection_5__4__5_, connection_5__4__4_, connection_5__4__3_,
         connection_5__4__2_, connection_5__4__1_, connection_5__4__0_,
         connection_5__5__31_, connection_5__5__30_, connection_5__5__29_,
         connection_5__5__28_, connection_5__5__27_, connection_5__5__26_,
         connection_5__5__25_, connection_5__5__24_, connection_5__5__23_,
         connection_5__5__22_, connection_5__5__21_, connection_5__5__20_,
         connection_5__5__19_, connection_5__5__18_, connection_5__5__17_,
         connection_5__5__16_, connection_5__5__15_, connection_5__5__14_,
         connection_5__5__13_, connection_5__5__12_, connection_5__5__11_,
         connection_5__5__10_, connection_5__5__9_, connection_5__5__8_,
         connection_5__5__7_, connection_5__5__6_, connection_5__5__5_,
         connection_5__5__4_, connection_5__5__3_, connection_5__5__2_,
         connection_5__5__1_, connection_5__5__0_, connection_5__6__31_,
         connection_5__6__30_, connection_5__6__29_, connection_5__6__28_,
         connection_5__6__27_, connection_5__6__26_, connection_5__6__25_,
         connection_5__6__24_, connection_5__6__23_, connection_5__6__22_,
         connection_5__6__21_, connection_5__6__20_, connection_5__6__19_,
         connection_5__6__18_, connection_5__6__17_, connection_5__6__16_,
         connection_5__6__15_, connection_5__6__14_, connection_5__6__13_,
         connection_5__6__12_, connection_5__6__11_, connection_5__6__10_,
         connection_5__6__9_, connection_5__6__8_, connection_5__6__7_,
         connection_5__6__6_, connection_5__6__5_, connection_5__6__4_,
         connection_5__6__3_, connection_5__6__2_, connection_5__6__1_,
         connection_5__6__0_, connection_5__7__31_, connection_5__7__30_,
         connection_5__7__29_, connection_5__7__28_, connection_5__7__27_,
         connection_5__7__26_, connection_5__7__25_, connection_5__7__24_,
         connection_5__7__23_, connection_5__7__22_, connection_5__7__21_,
         connection_5__7__20_, connection_5__7__19_, connection_5__7__18_,
         connection_5__7__17_, connection_5__7__16_, connection_5__7__15_,
         connection_5__7__14_, connection_5__7__13_, connection_5__7__12_,
         connection_5__7__11_, connection_5__7__10_, connection_5__7__9_,
         connection_5__7__8_, connection_5__7__7_, connection_5__7__6_,
         connection_5__7__5_, connection_5__7__4_, connection_5__7__3_,
         connection_5__7__2_, connection_5__7__1_, connection_5__7__0_,
         connection_5__8__31_, connection_5__8__30_, connection_5__8__29_,
         connection_5__8__28_, connection_5__8__27_, connection_5__8__26_,
         connection_5__8__25_, connection_5__8__24_, connection_5__8__23_,
         connection_5__8__22_, connection_5__8__21_, connection_5__8__20_,
         connection_5__8__19_, connection_5__8__18_, connection_5__8__17_,
         connection_5__8__16_, connection_5__8__15_, connection_5__8__14_,
         connection_5__8__13_, connection_5__8__12_, connection_5__8__11_,
         connection_5__8__10_, connection_5__8__9_, connection_5__8__8_,
         connection_5__8__7_, connection_5__8__6_, connection_5__8__5_,
         connection_5__8__4_, connection_5__8__3_, connection_5__8__2_,
         connection_5__8__1_, connection_5__8__0_, connection_5__9__31_,
         connection_5__9__30_, connection_5__9__29_, connection_5__9__28_,
         connection_5__9__27_, connection_5__9__26_, connection_5__9__25_,
         connection_5__9__24_, connection_5__9__23_, connection_5__9__22_,
         connection_5__9__21_, connection_5__9__20_, connection_5__9__19_,
         connection_5__9__18_, connection_5__9__17_, connection_5__9__16_,
         connection_5__9__15_, connection_5__9__14_, connection_5__9__13_,
         connection_5__9__12_, connection_5__9__11_, connection_5__9__10_,
         connection_5__9__9_, connection_5__9__8_, connection_5__9__7_,
         connection_5__9__6_, connection_5__9__5_, connection_5__9__4_,
         connection_5__9__3_, connection_5__9__2_, connection_5__9__1_,
         connection_5__9__0_, connection_5__10__31_, connection_5__10__30_,
         connection_5__10__29_, connection_5__10__28_, connection_5__10__27_,
         connection_5__10__26_, connection_5__10__25_, connection_5__10__24_,
         connection_5__10__23_, connection_5__10__22_, connection_5__10__21_,
         connection_5__10__20_, connection_5__10__19_, connection_5__10__18_,
         connection_5__10__17_, connection_5__10__16_, connection_5__10__15_,
         connection_5__10__14_, connection_5__10__13_, connection_5__10__12_,
         connection_5__10__11_, connection_5__10__10_, connection_5__10__9_,
         connection_5__10__8_, connection_5__10__7_, connection_5__10__6_,
         connection_5__10__5_, connection_5__10__4_, connection_5__10__3_,
         connection_5__10__2_, connection_5__10__1_, connection_5__10__0_,
         connection_5__11__31_, connection_5__11__30_, connection_5__11__29_,
         connection_5__11__28_, connection_5__11__27_, connection_5__11__26_,
         connection_5__11__25_, connection_5__11__24_, connection_5__11__23_,
         connection_5__11__22_, connection_5__11__21_, connection_5__11__20_,
         connection_5__11__19_, connection_5__11__18_, connection_5__11__17_,
         connection_5__11__16_, connection_5__11__15_, connection_5__11__14_,
         connection_5__11__13_, connection_5__11__12_, connection_5__11__11_,
         connection_5__11__10_, connection_5__11__9_, connection_5__11__8_,
         connection_5__11__7_, connection_5__11__6_, connection_5__11__5_,
         connection_5__11__4_, connection_5__11__3_, connection_5__11__2_,
         connection_5__11__1_, connection_5__11__0_, connection_5__12__31_,
         connection_5__12__30_, connection_5__12__29_, connection_5__12__28_,
         connection_5__12__27_, connection_5__12__26_, connection_5__12__25_,
         connection_5__12__24_, connection_5__12__23_, connection_5__12__22_,
         connection_5__12__21_, connection_5__12__20_, connection_5__12__19_,
         connection_5__12__18_, connection_5__12__17_, connection_5__12__16_,
         connection_5__12__15_, connection_5__12__14_, connection_5__12__13_,
         connection_5__12__12_, connection_5__12__11_, connection_5__12__10_,
         connection_5__12__9_, connection_5__12__8_, connection_5__12__7_,
         connection_5__12__6_, connection_5__12__5_, connection_5__12__4_,
         connection_5__12__3_, connection_5__12__2_, connection_5__12__1_,
         connection_5__12__0_, connection_5__13__31_, connection_5__13__30_,
         connection_5__13__29_, connection_5__13__28_, connection_5__13__27_,
         connection_5__13__26_, connection_5__13__25_, connection_5__13__24_,
         connection_5__13__23_, connection_5__13__22_, connection_5__13__21_,
         connection_5__13__20_, connection_5__13__19_, connection_5__13__18_,
         connection_5__13__17_, connection_5__13__16_, connection_5__13__15_,
         connection_5__13__14_, connection_5__13__13_, connection_5__13__12_,
         connection_5__13__11_, connection_5__13__10_, connection_5__13__9_,
         connection_5__13__8_, connection_5__13__7_, connection_5__13__6_,
         connection_5__13__5_, connection_5__13__4_, connection_5__13__3_,
         connection_5__13__2_, connection_5__13__1_, connection_5__13__0_,
         connection_5__14__31_, connection_5__14__30_, connection_5__14__29_,
         connection_5__14__28_, connection_5__14__27_, connection_5__14__26_,
         connection_5__14__25_, connection_5__14__24_, connection_5__14__23_,
         connection_5__14__22_, connection_5__14__21_, connection_5__14__20_,
         connection_5__14__19_, connection_5__14__18_, connection_5__14__17_,
         connection_5__14__16_, connection_5__14__15_, connection_5__14__14_,
         connection_5__14__13_, connection_5__14__12_, connection_5__14__11_,
         connection_5__14__10_, connection_5__14__9_, connection_5__14__8_,
         connection_5__14__7_, connection_5__14__6_, connection_5__14__5_,
         connection_5__14__4_, connection_5__14__3_, connection_5__14__2_,
         connection_5__14__1_, connection_5__14__0_, connection_5__15__31_,
         connection_5__15__30_, connection_5__15__29_, connection_5__15__28_,
         connection_5__15__27_, connection_5__15__26_, connection_5__15__25_,
         connection_5__15__24_, connection_5__15__23_, connection_5__15__22_,
         connection_5__15__21_, connection_5__15__20_, connection_5__15__19_,
         connection_5__15__18_, connection_5__15__17_, connection_5__15__16_,
         connection_5__15__15_, connection_5__15__14_, connection_5__15__13_,
         connection_5__15__12_, connection_5__15__11_, connection_5__15__10_,
         connection_5__15__9_, connection_5__15__8_, connection_5__15__7_,
         connection_5__15__6_, connection_5__15__5_, connection_5__15__4_,
         connection_5__15__3_, connection_5__15__2_, connection_5__15__1_,
         connection_5__15__0_, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30;
  wire   [95:0] cmd_pipeline_stage_0__pipeline_i_cmd_reg;
  wire   [79:0] cmd_pipeline_stage_1__pipeline_i_cmd_reg;
  wire   [63:0] cmd_pipeline_stage_2__pipeline_i_cmd_reg;
  wire   [47:0] cmd_pipeline_stage_3__pipeline_i_cmd_reg;
  wire   [31:0] cmd_pipeline_stage_4__pipeline_i_cmd_reg;
  wire   [15:0] cmd_pipeline_stage_5__pipeline_i_cmd_reg;

  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_0 first_stage_switch_0__first_stage ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[1:0]), .i_data_bus(
        i_data_bus[63:0]), .o_valid({connection_valid_0__1_, 
        connection_valid_0__0_}), .o_data_bus({connection_0__1__31_, 
        connection_0__1__30_, connection_0__1__29_, connection_0__1__28_, 
        connection_0__1__27_, connection_0__1__26_, connection_0__1__25_, 
        connection_0__1__24_, connection_0__1__23_, connection_0__1__22_, 
        connection_0__1__21_, connection_0__1__20_, connection_0__1__19_, 
        connection_0__1__18_, connection_0__1__17_, connection_0__1__16_, 
        connection_0__1__15_, connection_0__1__14_, connection_0__1__13_, 
        connection_0__1__12_, connection_0__1__11_, connection_0__1__10_, 
        connection_0__1__9_, connection_0__1__8_, connection_0__1__7_, 
        connection_0__1__6_, connection_0__1__5_, connection_0__1__4_, 
        connection_0__1__3_, connection_0__1__2_, connection_0__1__1_, 
        connection_0__1__0_, connection_0__0__31_, connection_0__0__30_, 
        connection_0__0__29_, connection_0__0__28_, connection_0__0__27_, 
        connection_0__0__26_, connection_0__0__25_, connection_0__0__24_, 
        connection_0__0__23_, connection_0__0__22_, connection_0__0__21_, 
        connection_0__0__20_, connection_0__0__19_, connection_0__0__18_, 
        connection_0__0__17_, connection_0__0__16_, connection_0__0__15_, 
        connection_0__0__14_, connection_0__0__13_, connection_0__0__12_, 
        connection_0__0__11_, connection_0__0__10_, connection_0__0__9_, 
        connection_0__0__8_, connection_0__0__7_, connection_0__0__6_, 
        connection_0__0__5_, connection_0__0__4_, connection_0__0__3_, 
        connection_0__0__2_, connection_0__0__1_, connection_0__0__0_}), 
        .i_en(i_en), .i_cmd(i_cmd[1:0]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_55 first_stage_switch_1__first_stage ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[3:2]), .i_data_bus(
        i_data_bus[127:64]), .o_valid({connection_valid_0__3_, 
        connection_valid_0__2_}), .o_data_bus({connection_0__3__31_, 
        connection_0__3__30_, connection_0__3__29_, connection_0__3__28_, 
        connection_0__3__27_, connection_0__3__26_, connection_0__3__25_, 
        connection_0__3__24_, connection_0__3__23_, connection_0__3__22_, 
        connection_0__3__21_, connection_0__3__20_, connection_0__3__19_, 
        connection_0__3__18_, connection_0__3__17_, connection_0__3__16_, 
        connection_0__3__15_, connection_0__3__14_, connection_0__3__13_, 
        connection_0__3__12_, connection_0__3__11_, connection_0__3__10_, 
        connection_0__3__9_, connection_0__3__8_, connection_0__3__7_, 
        connection_0__3__6_, connection_0__3__5_, connection_0__3__4_, 
        connection_0__3__3_, connection_0__3__2_, connection_0__3__1_, 
        connection_0__3__0_, connection_0__2__31_, connection_0__2__30_, 
        connection_0__2__29_, connection_0__2__28_, connection_0__2__27_, 
        connection_0__2__26_, connection_0__2__25_, connection_0__2__24_, 
        connection_0__2__23_, connection_0__2__22_, connection_0__2__21_, 
        connection_0__2__20_, connection_0__2__19_, connection_0__2__18_, 
        connection_0__2__17_, connection_0__2__16_, connection_0__2__15_, 
        connection_0__2__14_, connection_0__2__13_, connection_0__2__12_, 
        connection_0__2__11_, connection_0__2__10_, connection_0__2__9_, 
        connection_0__2__8_, connection_0__2__7_, connection_0__2__6_, 
        connection_0__2__5_, connection_0__2__4_, connection_0__2__3_, 
        connection_0__2__2_, connection_0__2__1_, connection_0__2__0_}), 
        .i_en(i_en), .i_cmd(i_cmd[3:2]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_54 first_stage_switch_2__first_stage ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[5:4]), .i_data_bus(
        i_data_bus[191:128]), .o_valid({connection_valid_0__5_, 
        connection_valid_0__4_}), .o_data_bus({connection_0__5__31_, 
        connection_0__5__30_, connection_0__5__29_, connection_0__5__28_, 
        connection_0__5__27_, connection_0__5__26_, connection_0__5__25_, 
        connection_0__5__24_, connection_0__5__23_, connection_0__5__22_, 
        connection_0__5__21_, connection_0__5__20_, connection_0__5__19_, 
        connection_0__5__18_, connection_0__5__17_, connection_0__5__16_, 
        connection_0__5__15_, connection_0__5__14_, connection_0__5__13_, 
        connection_0__5__12_, connection_0__5__11_, connection_0__5__10_, 
        connection_0__5__9_, connection_0__5__8_, connection_0__5__7_, 
        connection_0__5__6_, connection_0__5__5_, connection_0__5__4_, 
        connection_0__5__3_, connection_0__5__2_, connection_0__5__1_, 
        connection_0__5__0_, connection_0__4__31_, connection_0__4__30_, 
        connection_0__4__29_, connection_0__4__28_, connection_0__4__27_, 
        connection_0__4__26_, connection_0__4__25_, connection_0__4__24_, 
        connection_0__4__23_, connection_0__4__22_, connection_0__4__21_, 
        connection_0__4__20_, connection_0__4__19_, connection_0__4__18_, 
        connection_0__4__17_, connection_0__4__16_, connection_0__4__15_, 
        connection_0__4__14_, connection_0__4__13_, connection_0__4__12_, 
        connection_0__4__11_, connection_0__4__10_, connection_0__4__9_, 
        connection_0__4__8_, connection_0__4__7_, connection_0__4__6_, 
        connection_0__4__5_, connection_0__4__4_, connection_0__4__3_, 
        connection_0__4__2_, connection_0__4__1_, connection_0__4__0_}), 
        .i_en(i_en), .i_cmd(i_cmd[5:4]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_53 first_stage_switch_3__first_stage ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[7:6]), .i_data_bus(
        i_data_bus[255:192]), .o_valid({connection_valid_0__7_, 
        connection_valid_0__6_}), .o_data_bus({connection_0__7__31_, 
        connection_0__7__30_, connection_0__7__29_, connection_0__7__28_, 
        connection_0__7__27_, connection_0__7__26_, connection_0__7__25_, 
        connection_0__7__24_, connection_0__7__23_, connection_0__7__22_, 
        connection_0__7__21_, connection_0__7__20_, connection_0__7__19_, 
        connection_0__7__18_, connection_0__7__17_, connection_0__7__16_, 
        connection_0__7__15_, connection_0__7__14_, connection_0__7__13_, 
        connection_0__7__12_, connection_0__7__11_, connection_0__7__10_, 
        connection_0__7__9_, connection_0__7__8_, connection_0__7__7_, 
        connection_0__7__6_, connection_0__7__5_, connection_0__7__4_, 
        connection_0__7__3_, connection_0__7__2_, connection_0__7__1_, 
        connection_0__7__0_, connection_0__6__31_, connection_0__6__30_, 
        connection_0__6__29_, connection_0__6__28_, connection_0__6__27_, 
        connection_0__6__26_, connection_0__6__25_, connection_0__6__24_, 
        connection_0__6__23_, connection_0__6__22_, connection_0__6__21_, 
        connection_0__6__20_, connection_0__6__19_, connection_0__6__18_, 
        connection_0__6__17_, connection_0__6__16_, connection_0__6__15_, 
        connection_0__6__14_, connection_0__6__13_, connection_0__6__12_, 
        connection_0__6__11_, connection_0__6__10_, connection_0__6__9_, 
        connection_0__6__8_, connection_0__6__7_, connection_0__6__6_, 
        connection_0__6__5_, connection_0__6__4_, connection_0__6__3_, 
        connection_0__6__2_, connection_0__6__1_, connection_0__6__0_}), 
        .i_en(i_en), .i_cmd(i_cmd[7:6]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_52 first_stage_switch_4__first_stage ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[9:8]), .i_data_bus(
        i_data_bus[319:256]), .o_valid({connection_valid_0__9_, 
        connection_valid_0__8_}), .o_data_bus({connection_0__9__31_, 
        connection_0__9__30_, connection_0__9__29_, connection_0__9__28_, 
        connection_0__9__27_, connection_0__9__26_, connection_0__9__25_, 
        connection_0__9__24_, connection_0__9__23_, connection_0__9__22_, 
        connection_0__9__21_, connection_0__9__20_, connection_0__9__19_, 
        connection_0__9__18_, connection_0__9__17_, connection_0__9__16_, 
        connection_0__9__15_, connection_0__9__14_, connection_0__9__13_, 
        connection_0__9__12_, connection_0__9__11_, connection_0__9__10_, 
        connection_0__9__9_, connection_0__9__8_, connection_0__9__7_, 
        connection_0__9__6_, connection_0__9__5_, connection_0__9__4_, 
        connection_0__9__3_, connection_0__9__2_, connection_0__9__1_, 
        connection_0__9__0_, connection_0__8__31_, connection_0__8__30_, 
        connection_0__8__29_, connection_0__8__28_, connection_0__8__27_, 
        connection_0__8__26_, connection_0__8__25_, connection_0__8__24_, 
        connection_0__8__23_, connection_0__8__22_, connection_0__8__21_, 
        connection_0__8__20_, connection_0__8__19_, connection_0__8__18_, 
        connection_0__8__17_, connection_0__8__16_, connection_0__8__15_, 
        connection_0__8__14_, connection_0__8__13_, connection_0__8__12_, 
        connection_0__8__11_, connection_0__8__10_, connection_0__8__9_, 
        connection_0__8__8_, connection_0__8__7_, connection_0__8__6_, 
        connection_0__8__5_, connection_0__8__4_, connection_0__8__3_, 
        connection_0__8__2_, connection_0__8__1_, connection_0__8__0_}), 
        .i_en(i_en), .i_cmd(i_cmd[9:8]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_51 first_stage_switch_5__first_stage ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[11:10]), .i_data_bus(
        i_data_bus[383:320]), .o_valid({connection_valid_0__11_, 
        connection_valid_0__10_}), .o_data_bus({connection_0__11__31_, 
        connection_0__11__30_, connection_0__11__29_, connection_0__11__28_, 
        connection_0__11__27_, connection_0__11__26_, connection_0__11__25_, 
        connection_0__11__24_, connection_0__11__23_, connection_0__11__22_, 
        connection_0__11__21_, connection_0__11__20_, connection_0__11__19_, 
        connection_0__11__18_, connection_0__11__17_, connection_0__11__16_, 
        connection_0__11__15_, connection_0__11__14_, connection_0__11__13_, 
        connection_0__11__12_, connection_0__11__11_, connection_0__11__10_, 
        connection_0__11__9_, connection_0__11__8_, connection_0__11__7_, 
        connection_0__11__6_, connection_0__11__5_, connection_0__11__4_, 
        connection_0__11__3_, connection_0__11__2_, connection_0__11__1_, 
        connection_0__11__0_, connection_0__10__31_, connection_0__10__30_, 
        connection_0__10__29_, connection_0__10__28_, connection_0__10__27_, 
        connection_0__10__26_, connection_0__10__25_, connection_0__10__24_, 
        connection_0__10__23_, connection_0__10__22_, connection_0__10__21_, 
        connection_0__10__20_, connection_0__10__19_, connection_0__10__18_, 
        connection_0__10__17_, connection_0__10__16_, connection_0__10__15_, 
        connection_0__10__14_, connection_0__10__13_, connection_0__10__12_, 
        connection_0__10__11_, connection_0__10__10_, connection_0__10__9_, 
        connection_0__10__8_, connection_0__10__7_, connection_0__10__6_, 
        connection_0__10__5_, connection_0__10__4_, connection_0__10__3_, 
        connection_0__10__2_, connection_0__10__1_, connection_0__10__0_}), 
        .i_en(i_en), .i_cmd(i_cmd[11:10]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_50 first_stage_switch_6__first_stage ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[13:12]), .i_data_bus(
        i_data_bus[447:384]), .o_valid({connection_valid_0__13_, 
        connection_valid_0__12_}), .o_data_bus({connection_0__13__31_, 
        connection_0__13__30_, connection_0__13__29_, connection_0__13__28_, 
        connection_0__13__27_, connection_0__13__26_, connection_0__13__25_, 
        connection_0__13__24_, connection_0__13__23_, connection_0__13__22_, 
        connection_0__13__21_, connection_0__13__20_, connection_0__13__19_, 
        connection_0__13__18_, connection_0__13__17_, connection_0__13__16_, 
        connection_0__13__15_, connection_0__13__14_, connection_0__13__13_, 
        connection_0__13__12_, connection_0__13__11_, connection_0__13__10_, 
        connection_0__13__9_, connection_0__13__8_, connection_0__13__7_, 
        connection_0__13__6_, connection_0__13__5_, connection_0__13__4_, 
        connection_0__13__3_, connection_0__13__2_, connection_0__13__1_, 
        connection_0__13__0_, connection_0__12__31_, connection_0__12__30_, 
        connection_0__12__29_, connection_0__12__28_, connection_0__12__27_, 
        connection_0__12__26_, connection_0__12__25_, connection_0__12__24_, 
        connection_0__12__23_, connection_0__12__22_, connection_0__12__21_, 
        connection_0__12__20_, connection_0__12__19_, connection_0__12__18_, 
        connection_0__12__17_, connection_0__12__16_, connection_0__12__15_, 
        connection_0__12__14_, connection_0__12__13_, connection_0__12__12_, 
        connection_0__12__11_, connection_0__12__10_, connection_0__12__9_, 
        connection_0__12__8_, connection_0__12__7_, connection_0__12__6_, 
        connection_0__12__5_, connection_0__12__4_, connection_0__12__3_, 
        connection_0__12__2_, connection_0__12__1_, connection_0__12__0_}), 
        .i_en(i_en), .i_cmd(i_cmd[13:12]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_49 first_stage_switch_7__first_stage ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[15:14]), .i_data_bus(
        i_data_bus[511:448]), .o_valid({connection_valid_0__15_, 
        connection_valid_0__14_}), .o_data_bus({connection_0__15__31_, 
        connection_0__15__30_, connection_0__15__29_, connection_0__15__28_, 
        connection_0__15__27_, connection_0__15__26_, connection_0__15__25_, 
        connection_0__15__24_, connection_0__15__23_, connection_0__15__22_, 
        connection_0__15__21_, connection_0__15__20_, connection_0__15__19_, 
        connection_0__15__18_, connection_0__15__17_, connection_0__15__16_, 
        connection_0__15__15_, connection_0__15__14_, connection_0__15__13_, 
        connection_0__15__12_, connection_0__15__11_, connection_0__15__10_, 
        connection_0__15__9_, connection_0__15__8_, connection_0__15__7_, 
        connection_0__15__6_, connection_0__15__5_, connection_0__15__4_, 
        connection_0__15__3_, connection_0__15__2_, connection_0__15__1_, 
        connection_0__15__0_, connection_0__14__31_, connection_0__14__30_, 
        connection_0__14__29_, connection_0__14__28_, connection_0__14__27_, 
        connection_0__14__26_, connection_0__14__25_, connection_0__14__24_, 
        connection_0__14__23_, connection_0__14__22_, connection_0__14__21_, 
        connection_0__14__20_, connection_0__14__19_, connection_0__14__18_, 
        connection_0__14__17_, connection_0__14__16_, connection_0__14__15_, 
        connection_0__14__14_, connection_0__14__13_, connection_0__14__12_, 
        connection_0__14__11_, connection_0__14__10_, connection_0__14__9_, 
        connection_0__14__8_, connection_0__14__7_, connection_0__14__6_, 
        connection_0__14__5_, connection_0__14__4_, connection_0__14__3_, 
        connection_0__14__2_, connection_0__14__1_, connection_0__14__0_}), 
        .i_en(i_en), .i_cmd(i_cmd[15:14]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_48 first_half_stages_0__group_first_half_0__switch_first_half_0__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__2_, 
        connection_valid_0__0_}), .i_data_bus({connection_0__2__31_, 
        connection_0__2__30_, connection_0__2__29_, connection_0__2__28_, 
        connection_0__2__27_, connection_0__2__26_, connection_0__2__25_, 
        connection_0__2__24_, connection_0__2__23_, connection_0__2__22_, 
        connection_0__2__21_, connection_0__2__20_, connection_0__2__19_, 
        connection_0__2__18_, connection_0__2__17_, connection_0__2__16_, 
        connection_0__2__15_, connection_0__2__14_, connection_0__2__13_, 
        connection_0__2__12_, connection_0__2__11_, connection_0__2__10_, 
        connection_0__2__9_, connection_0__2__8_, connection_0__2__7_, 
        connection_0__2__6_, connection_0__2__5_, connection_0__2__4_, 
        connection_0__2__3_, connection_0__2__2_, connection_0__2__1_, 
        connection_0__2__0_, connection_0__0__31_, connection_0__0__30_, 
        connection_0__0__29_, connection_0__0__28_, connection_0__0__27_, 
        connection_0__0__26_, connection_0__0__25_, connection_0__0__24_, 
        connection_0__0__23_, connection_0__0__22_, connection_0__0__21_, 
        connection_0__0__20_, connection_0__0__19_, connection_0__0__18_, 
        connection_0__0__17_, connection_0__0__16_, connection_0__0__15_, 
        connection_0__0__14_, connection_0__0__13_, connection_0__0__12_, 
        connection_0__0__11_, connection_0__0__10_, connection_0__0__9_, 
        connection_0__0__8_, connection_0__0__7_, connection_0__0__6_, 
        connection_0__0__5_, connection_0__0__4_, connection_0__0__3_, 
        connection_0__0__2_, connection_0__0__1_, connection_0__0__0_}), 
        .o_valid({connection_valid_1__1_, connection_valid_1__0_}), 
        .o_data_bus({connection_1__1__31_, connection_1__1__30_, 
        connection_1__1__29_, connection_1__1__28_, connection_1__1__27_, 
        connection_1__1__26_, connection_1__1__25_, connection_1__1__24_, 
        connection_1__1__23_, connection_1__1__22_, connection_1__1__21_, 
        connection_1__1__20_, connection_1__1__19_, connection_1__1__18_, 
        connection_1__1__17_, connection_1__1__16_, connection_1__1__15_, 
        connection_1__1__14_, connection_1__1__13_, connection_1__1__12_, 
        connection_1__1__11_, connection_1__1__10_, connection_1__1__9_, 
        connection_1__1__8_, connection_1__1__7_, connection_1__1__6_, 
        connection_1__1__5_, connection_1__1__4_, connection_1__1__3_, 
        connection_1__1__2_, connection_1__1__1_, connection_1__1__0_, 
        connection_1__0__31_, connection_1__0__30_, connection_1__0__29_, 
        connection_1__0__28_, connection_1__0__27_, connection_1__0__26_, 
        connection_1__0__25_, connection_1__0__24_, connection_1__0__23_, 
        connection_1__0__22_, connection_1__0__21_, connection_1__0__20_, 
        connection_1__0__19_, connection_1__0__18_, connection_1__0__17_, 
        connection_1__0__16_, connection_1__0__15_, connection_1__0__14_, 
        connection_1__0__13_, connection_1__0__12_, connection_1__0__11_, 
        connection_1__0__10_, connection_1__0__9_, connection_1__0__8_, 
        connection_1__0__7_, connection_1__0__6_, connection_1__0__5_, 
        connection_1__0__4_, connection_1__0__3_, connection_1__0__2_, 
        connection_1__0__1_, connection_1__0__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[95:94]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_47 first_half_stages_0__group_first_half_0__switch_first_half_1__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__6_, 
        connection_valid_0__4_}), .i_data_bus({connection_0__6__31_, 
        connection_0__6__30_, connection_0__6__29_, connection_0__6__28_, 
        connection_0__6__27_, connection_0__6__26_, connection_0__6__25_, 
        connection_0__6__24_, connection_0__6__23_, connection_0__6__22_, 
        connection_0__6__21_, connection_0__6__20_, connection_0__6__19_, 
        connection_0__6__18_, connection_0__6__17_, connection_0__6__16_, 
        connection_0__6__15_, connection_0__6__14_, connection_0__6__13_, 
        connection_0__6__12_, connection_0__6__11_, connection_0__6__10_, 
        connection_0__6__9_, connection_0__6__8_, connection_0__6__7_, 
        connection_0__6__6_, connection_0__6__5_, connection_0__6__4_, 
        connection_0__6__3_, connection_0__6__2_, connection_0__6__1_, 
        connection_0__6__0_, connection_0__4__31_, connection_0__4__30_, 
        connection_0__4__29_, connection_0__4__28_, connection_0__4__27_, 
        connection_0__4__26_, connection_0__4__25_, connection_0__4__24_, 
        connection_0__4__23_, connection_0__4__22_, connection_0__4__21_, 
        connection_0__4__20_, connection_0__4__19_, connection_0__4__18_, 
        connection_0__4__17_, connection_0__4__16_, connection_0__4__15_, 
        connection_0__4__14_, connection_0__4__13_, connection_0__4__12_, 
        connection_0__4__11_, connection_0__4__10_, connection_0__4__9_, 
        connection_0__4__8_, connection_0__4__7_, connection_0__4__6_, 
        connection_0__4__5_, connection_0__4__4_, connection_0__4__3_, 
        connection_0__4__2_, connection_0__4__1_, connection_0__4__0_}), 
        .o_valid({connection_valid_1__3_, connection_valid_1__2_}), 
        .o_data_bus({connection_1__3__31_, connection_1__3__30_, 
        connection_1__3__29_, connection_1__3__28_, connection_1__3__27_, 
        connection_1__3__26_, connection_1__3__25_, connection_1__3__24_, 
        connection_1__3__23_, connection_1__3__22_, connection_1__3__21_, 
        connection_1__3__20_, connection_1__3__19_, connection_1__3__18_, 
        connection_1__3__17_, connection_1__3__16_, connection_1__3__15_, 
        connection_1__3__14_, connection_1__3__13_, connection_1__3__12_, 
        connection_1__3__11_, connection_1__3__10_, connection_1__3__9_, 
        connection_1__3__8_, connection_1__3__7_, connection_1__3__6_, 
        connection_1__3__5_, connection_1__3__4_, connection_1__3__3_, 
        connection_1__3__2_, connection_1__3__1_, connection_1__3__0_, 
        connection_1__2__31_, connection_1__2__30_, connection_1__2__29_, 
        connection_1__2__28_, connection_1__2__27_, connection_1__2__26_, 
        connection_1__2__25_, connection_1__2__24_, connection_1__2__23_, 
        connection_1__2__22_, connection_1__2__21_, connection_1__2__20_, 
        connection_1__2__19_, connection_1__2__18_, connection_1__2__17_, 
        connection_1__2__16_, connection_1__2__15_, connection_1__2__14_, 
        connection_1__2__13_, connection_1__2__12_, connection_1__2__11_, 
        connection_1__2__10_, connection_1__2__9_, connection_1__2__8_, 
        connection_1__2__7_, connection_1__2__6_, connection_1__2__5_, 
        connection_1__2__4_, connection_1__2__3_, connection_1__2__2_, 
        connection_1__2__1_, connection_1__2__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[93:92]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_46 first_half_stages_0__group_first_half_0__switch_first_half_2__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__10_, 
        connection_valid_0__8_}), .i_data_bus({connection_0__10__31_, 
        connection_0__10__30_, connection_0__10__29_, connection_0__10__28_, 
        connection_0__10__27_, connection_0__10__26_, connection_0__10__25_, 
        connection_0__10__24_, connection_0__10__23_, connection_0__10__22_, 
        connection_0__10__21_, connection_0__10__20_, connection_0__10__19_, 
        connection_0__10__18_, connection_0__10__17_, connection_0__10__16_, 
        connection_0__10__15_, connection_0__10__14_, connection_0__10__13_, 
        connection_0__10__12_, connection_0__10__11_, connection_0__10__10_, 
        connection_0__10__9_, connection_0__10__8_, connection_0__10__7_, 
        connection_0__10__6_, connection_0__10__5_, connection_0__10__4_, 
        connection_0__10__3_, connection_0__10__2_, connection_0__10__1_, 
        connection_0__10__0_, connection_0__8__31_, connection_0__8__30_, 
        connection_0__8__29_, connection_0__8__28_, connection_0__8__27_, 
        connection_0__8__26_, connection_0__8__25_, connection_0__8__24_, 
        connection_0__8__23_, connection_0__8__22_, connection_0__8__21_, 
        connection_0__8__20_, connection_0__8__19_, connection_0__8__18_, 
        connection_0__8__17_, connection_0__8__16_, connection_0__8__15_, 
        connection_0__8__14_, connection_0__8__13_, connection_0__8__12_, 
        connection_0__8__11_, connection_0__8__10_, connection_0__8__9_, 
        connection_0__8__8_, connection_0__8__7_, connection_0__8__6_, 
        connection_0__8__5_, connection_0__8__4_, connection_0__8__3_, 
        connection_0__8__2_, connection_0__8__1_, connection_0__8__0_}), 
        .o_valid({connection_valid_1__5_, connection_valid_1__4_}), 
        .o_data_bus({connection_1__5__31_, connection_1__5__30_, 
        connection_1__5__29_, connection_1__5__28_, connection_1__5__27_, 
        connection_1__5__26_, connection_1__5__25_, connection_1__5__24_, 
        connection_1__5__23_, connection_1__5__22_, connection_1__5__21_, 
        connection_1__5__20_, connection_1__5__19_, connection_1__5__18_, 
        connection_1__5__17_, connection_1__5__16_, connection_1__5__15_, 
        connection_1__5__14_, connection_1__5__13_, connection_1__5__12_, 
        connection_1__5__11_, connection_1__5__10_, connection_1__5__9_, 
        connection_1__5__8_, connection_1__5__7_, connection_1__5__6_, 
        connection_1__5__5_, connection_1__5__4_, connection_1__5__3_, 
        connection_1__5__2_, connection_1__5__1_, connection_1__5__0_, 
        connection_1__4__31_, connection_1__4__30_, connection_1__4__29_, 
        connection_1__4__28_, connection_1__4__27_, connection_1__4__26_, 
        connection_1__4__25_, connection_1__4__24_, connection_1__4__23_, 
        connection_1__4__22_, connection_1__4__21_, connection_1__4__20_, 
        connection_1__4__19_, connection_1__4__18_, connection_1__4__17_, 
        connection_1__4__16_, connection_1__4__15_, connection_1__4__14_, 
        connection_1__4__13_, connection_1__4__12_, connection_1__4__11_, 
        connection_1__4__10_, connection_1__4__9_, connection_1__4__8_, 
        connection_1__4__7_, connection_1__4__6_, connection_1__4__5_, 
        connection_1__4__4_, connection_1__4__3_, connection_1__4__2_, 
        connection_1__4__1_, connection_1__4__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[91:90]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_45 first_half_stages_0__group_first_half_0__switch_first_half_3__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__14_, 
        connection_valid_0__12_}), .i_data_bus({connection_0__14__31_, 
        connection_0__14__30_, connection_0__14__29_, connection_0__14__28_, 
        connection_0__14__27_, connection_0__14__26_, connection_0__14__25_, 
        connection_0__14__24_, connection_0__14__23_, connection_0__14__22_, 
        connection_0__14__21_, connection_0__14__20_, connection_0__14__19_, 
        connection_0__14__18_, connection_0__14__17_, connection_0__14__16_, 
        connection_0__14__15_, connection_0__14__14_, connection_0__14__13_, 
        connection_0__14__12_, connection_0__14__11_, connection_0__14__10_, 
        connection_0__14__9_, connection_0__14__8_, connection_0__14__7_, 
        connection_0__14__6_, connection_0__14__5_, connection_0__14__4_, 
        connection_0__14__3_, connection_0__14__2_, connection_0__14__1_, 
        connection_0__14__0_, connection_0__12__31_, connection_0__12__30_, 
        connection_0__12__29_, connection_0__12__28_, connection_0__12__27_, 
        connection_0__12__26_, connection_0__12__25_, connection_0__12__24_, 
        connection_0__12__23_, connection_0__12__22_, connection_0__12__21_, 
        connection_0__12__20_, connection_0__12__19_, connection_0__12__18_, 
        connection_0__12__17_, connection_0__12__16_, connection_0__12__15_, 
        connection_0__12__14_, connection_0__12__13_, connection_0__12__12_, 
        connection_0__12__11_, connection_0__12__10_, connection_0__12__9_, 
        connection_0__12__8_, connection_0__12__7_, connection_0__12__6_, 
        connection_0__12__5_, connection_0__12__4_, connection_0__12__3_, 
        connection_0__12__2_, connection_0__12__1_, connection_0__12__0_}), 
        .o_valid({connection_valid_1__7_, connection_valid_1__6_}), 
        .o_data_bus({connection_1__7__31_, connection_1__7__30_, 
        connection_1__7__29_, connection_1__7__28_, connection_1__7__27_, 
        connection_1__7__26_, connection_1__7__25_, connection_1__7__24_, 
        connection_1__7__23_, connection_1__7__22_, connection_1__7__21_, 
        connection_1__7__20_, connection_1__7__19_, connection_1__7__18_, 
        connection_1__7__17_, connection_1__7__16_, connection_1__7__15_, 
        connection_1__7__14_, connection_1__7__13_, connection_1__7__12_, 
        connection_1__7__11_, connection_1__7__10_, connection_1__7__9_, 
        connection_1__7__8_, connection_1__7__7_, connection_1__7__6_, 
        connection_1__7__5_, connection_1__7__4_, connection_1__7__3_, 
        connection_1__7__2_, connection_1__7__1_, connection_1__7__0_, 
        connection_1__6__31_, connection_1__6__30_, connection_1__6__29_, 
        connection_1__6__28_, connection_1__6__27_, connection_1__6__26_, 
        connection_1__6__25_, connection_1__6__24_, connection_1__6__23_, 
        connection_1__6__22_, connection_1__6__21_, connection_1__6__20_, 
        connection_1__6__19_, connection_1__6__18_, connection_1__6__17_, 
        connection_1__6__16_, connection_1__6__15_, connection_1__6__14_, 
        connection_1__6__13_, connection_1__6__12_, connection_1__6__11_, 
        connection_1__6__10_, connection_1__6__9_, connection_1__6__8_, 
        connection_1__6__7_, connection_1__6__6_, connection_1__6__5_, 
        connection_1__6__4_, connection_1__6__3_, connection_1__6__2_, 
        connection_1__6__1_, connection_1__6__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[89:88]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_44 first_half_stages_0__group_first_half_0__switch_first_half_4__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__3_, 
        connection_valid_0__1_}), .i_data_bus({connection_0__3__31_, 
        connection_0__3__30_, connection_0__3__29_, connection_0__3__28_, 
        connection_0__3__27_, connection_0__3__26_, connection_0__3__25_, 
        connection_0__3__24_, connection_0__3__23_, connection_0__3__22_, 
        connection_0__3__21_, connection_0__3__20_, connection_0__3__19_, 
        connection_0__3__18_, connection_0__3__17_, connection_0__3__16_, 
        connection_0__3__15_, connection_0__3__14_, connection_0__3__13_, 
        connection_0__3__12_, connection_0__3__11_, connection_0__3__10_, 
        connection_0__3__9_, connection_0__3__8_, connection_0__3__7_, 
        connection_0__3__6_, connection_0__3__5_, connection_0__3__4_, 
        connection_0__3__3_, connection_0__3__2_, connection_0__3__1_, 
        connection_0__3__0_, connection_0__1__31_, connection_0__1__30_, 
        connection_0__1__29_, connection_0__1__28_, connection_0__1__27_, 
        connection_0__1__26_, connection_0__1__25_, connection_0__1__24_, 
        connection_0__1__23_, connection_0__1__22_, connection_0__1__21_, 
        connection_0__1__20_, connection_0__1__19_, connection_0__1__18_, 
        connection_0__1__17_, connection_0__1__16_, connection_0__1__15_, 
        connection_0__1__14_, connection_0__1__13_, connection_0__1__12_, 
        connection_0__1__11_, connection_0__1__10_, connection_0__1__9_, 
        connection_0__1__8_, connection_0__1__7_, connection_0__1__6_, 
        connection_0__1__5_, connection_0__1__4_, connection_0__1__3_, 
        connection_0__1__2_, connection_0__1__1_, connection_0__1__0_}), 
        .o_valid({connection_valid_1__9_, connection_valid_1__8_}), 
        .o_data_bus({connection_1__9__31_, connection_1__9__30_, 
        connection_1__9__29_, connection_1__9__28_, connection_1__9__27_, 
        connection_1__9__26_, connection_1__9__25_, connection_1__9__24_, 
        connection_1__9__23_, connection_1__9__22_, connection_1__9__21_, 
        connection_1__9__20_, connection_1__9__19_, connection_1__9__18_, 
        connection_1__9__17_, connection_1__9__16_, connection_1__9__15_, 
        connection_1__9__14_, connection_1__9__13_, connection_1__9__12_, 
        connection_1__9__11_, connection_1__9__10_, connection_1__9__9_, 
        connection_1__9__8_, connection_1__9__7_, connection_1__9__6_, 
        connection_1__9__5_, connection_1__9__4_, connection_1__9__3_, 
        connection_1__9__2_, connection_1__9__1_, connection_1__9__0_, 
        connection_1__8__31_, connection_1__8__30_, connection_1__8__29_, 
        connection_1__8__28_, connection_1__8__27_, connection_1__8__26_, 
        connection_1__8__25_, connection_1__8__24_, connection_1__8__23_, 
        connection_1__8__22_, connection_1__8__21_, connection_1__8__20_, 
        connection_1__8__19_, connection_1__8__18_, connection_1__8__17_, 
        connection_1__8__16_, connection_1__8__15_, connection_1__8__14_, 
        connection_1__8__13_, connection_1__8__12_, connection_1__8__11_, 
        connection_1__8__10_, connection_1__8__9_, connection_1__8__8_, 
        connection_1__8__7_, connection_1__8__6_, connection_1__8__5_, 
        connection_1__8__4_, connection_1__8__3_, connection_1__8__2_, 
        connection_1__8__1_, connection_1__8__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[87:86]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_43 first_half_stages_0__group_first_half_0__switch_first_half_5__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__7_, 
        connection_valid_0__5_}), .i_data_bus({connection_0__7__31_, 
        connection_0__7__30_, connection_0__7__29_, connection_0__7__28_, 
        connection_0__7__27_, connection_0__7__26_, connection_0__7__25_, 
        connection_0__7__24_, connection_0__7__23_, connection_0__7__22_, 
        connection_0__7__21_, connection_0__7__20_, connection_0__7__19_, 
        connection_0__7__18_, connection_0__7__17_, connection_0__7__16_, 
        connection_0__7__15_, connection_0__7__14_, connection_0__7__13_, 
        connection_0__7__12_, connection_0__7__11_, connection_0__7__10_, 
        connection_0__7__9_, connection_0__7__8_, connection_0__7__7_, 
        connection_0__7__6_, connection_0__7__5_, connection_0__7__4_, 
        connection_0__7__3_, connection_0__7__2_, connection_0__7__1_, 
        connection_0__7__0_, connection_0__5__31_, connection_0__5__30_, 
        connection_0__5__29_, connection_0__5__28_, connection_0__5__27_, 
        connection_0__5__26_, connection_0__5__25_, connection_0__5__24_, 
        connection_0__5__23_, connection_0__5__22_, connection_0__5__21_, 
        connection_0__5__20_, connection_0__5__19_, connection_0__5__18_, 
        connection_0__5__17_, connection_0__5__16_, connection_0__5__15_, 
        connection_0__5__14_, connection_0__5__13_, connection_0__5__12_, 
        connection_0__5__11_, connection_0__5__10_, connection_0__5__9_, 
        connection_0__5__8_, connection_0__5__7_, connection_0__5__6_, 
        connection_0__5__5_, connection_0__5__4_, connection_0__5__3_, 
        connection_0__5__2_, connection_0__5__1_, connection_0__5__0_}), 
        .o_valid({connection_valid_1__11_, connection_valid_1__10_}), 
        .o_data_bus({connection_1__11__31_, connection_1__11__30_, 
        connection_1__11__29_, connection_1__11__28_, connection_1__11__27_, 
        connection_1__11__26_, connection_1__11__25_, connection_1__11__24_, 
        connection_1__11__23_, connection_1__11__22_, connection_1__11__21_, 
        connection_1__11__20_, connection_1__11__19_, connection_1__11__18_, 
        connection_1__11__17_, connection_1__11__16_, connection_1__11__15_, 
        connection_1__11__14_, connection_1__11__13_, connection_1__11__12_, 
        connection_1__11__11_, connection_1__11__10_, connection_1__11__9_, 
        connection_1__11__8_, connection_1__11__7_, connection_1__11__6_, 
        connection_1__11__5_, connection_1__11__4_, connection_1__11__3_, 
        connection_1__11__2_, connection_1__11__1_, connection_1__11__0_, 
        connection_1__10__31_, connection_1__10__30_, connection_1__10__29_, 
        connection_1__10__28_, connection_1__10__27_, connection_1__10__26_, 
        connection_1__10__25_, connection_1__10__24_, connection_1__10__23_, 
        connection_1__10__22_, connection_1__10__21_, connection_1__10__20_, 
        connection_1__10__19_, connection_1__10__18_, connection_1__10__17_, 
        connection_1__10__16_, connection_1__10__15_, connection_1__10__14_, 
        connection_1__10__13_, connection_1__10__12_, connection_1__10__11_, 
        connection_1__10__10_, connection_1__10__9_, connection_1__10__8_, 
        connection_1__10__7_, connection_1__10__6_, connection_1__10__5_, 
        connection_1__10__4_, connection_1__10__3_, connection_1__10__2_, 
        connection_1__10__1_, connection_1__10__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[85:84]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_42 first_half_stages_0__group_first_half_0__switch_first_half_6__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__11_, 
        connection_valid_0__9_}), .i_data_bus({connection_0__11__31_, 
        connection_0__11__30_, connection_0__11__29_, connection_0__11__28_, 
        connection_0__11__27_, connection_0__11__26_, connection_0__11__25_, 
        connection_0__11__24_, connection_0__11__23_, connection_0__11__22_, 
        connection_0__11__21_, connection_0__11__20_, connection_0__11__19_, 
        connection_0__11__18_, connection_0__11__17_, connection_0__11__16_, 
        connection_0__11__15_, connection_0__11__14_, connection_0__11__13_, 
        connection_0__11__12_, connection_0__11__11_, connection_0__11__10_, 
        connection_0__11__9_, connection_0__11__8_, connection_0__11__7_, 
        connection_0__11__6_, connection_0__11__5_, connection_0__11__4_, 
        connection_0__11__3_, connection_0__11__2_, connection_0__11__1_, 
        connection_0__11__0_, connection_0__9__31_, connection_0__9__30_, 
        connection_0__9__29_, connection_0__9__28_, connection_0__9__27_, 
        connection_0__9__26_, connection_0__9__25_, connection_0__9__24_, 
        connection_0__9__23_, connection_0__9__22_, connection_0__9__21_, 
        connection_0__9__20_, connection_0__9__19_, connection_0__9__18_, 
        connection_0__9__17_, connection_0__9__16_, connection_0__9__15_, 
        connection_0__9__14_, connection_0__9__13_, connection_0__9__12_, 
        connection_0__9__11_, connection_0__9__10_, connection_0__9__9_, 
        connection_0__9__8_, connection_0__9__7_, connection_0__9__6_, 
        connection_0__9__5_, connection_0__9__4_, connection_0__9__3_, 
        connection_0__9__2_, connection_0__9__1_, connection_0__9__0_}), 
        .o_valid({connection_valid_1__13_, connection_valid_1__12_}), 
        .o_data_bus({connection_1__13__31_, connection_1__13__30_, 
        connection_1__13__29_, connection_1__13__28_, connection_1__13__27_, 
        connection_1__13__26_, connection_1__13__25_, connection_1__13__24_, 
        connection_1__13__23_, connection_1__13__22_, connection_1__13__21_, 
        connection_1__13__20_, connection_1__13__19_, connection_1__13__18_, 
        connection_1__13__17_, connection_1__13__16_, connection_1__13__15_, 
        connection_1__13__14_, connection_1__13__13_, connection_1__13__12_, 
        connection_1__13__11_, connection_1__13__10_, connection_1__13__9_, 
        connection_1__13__8_, connection_1__13__7_, connection_1__13__6_, 
        connection_1__13__5_, connection_1__13__4_, connection_1__13__3_, 
        connection_1__13__2_, connection_1__13__1_, connection_1__13__0_, 
        connection_1__12__31_, connection_1__12__30_, connection_1__12__29_, 
        connection_1__12__28_, connection_1__12__27_, connection_1__12__26_, 
        connection_1__12__25_, connection_1__12__24_, connection_1__12__23_, 
        connection_1__12__22_, connection_1__12__21_, connection_1__12__20_, 
        connection_1__12__19_, connection_1__12__18_, connection_1__12__17_, 
        connection_1__12__16_, connection_1__12__15_, connection_1__12__14_, 
        connection_1__12__13_, connection_1__12__12_, connection_1__12__11_, 
        connection_1__12__10_, connection_1__12__9_, connection_1__12__8_, 
        connection_1__12__7_, connection_1__12__6_, connection_1__12__5_, 
        connection_1__12__4_, connection_1__12__3_, connection_1__12__2_, 
        connection_1__12__1_, connection_1__12__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[83:82]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_41 first_half_stages_0__group_first_half_0__switch_first_half_7__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__15_, 
        connection_valid_0__13_}), .i_data_bus({connection_0__15__31_, 
        connection_0__15__30_, connection_0__15__29_, connection_0__15__28_, 
        connection_0__15__27_, connection_0__15__26_, connection_0__15__25_, 
        connection_0__15__24_, connection_0__15__23_, connection_0__15__22_, 
        connection_0__15__21_, connection_0__15__20_, connection_0__15__19_, 
        connection_0__15__18_, connection_0__15__17_, connection_0__15__16_, 
        connection_0__15__15_, connection_0__15__14_, connection_0__15__13_, 
        connection_0__15__12_, connection_0__15__11_, connection_0__15__10_, 
        connection_0__15__9_, connection_0__15__8_, connection_0__15__7_, 
        connection_0__15__6_, connection_0__15__5_, connection_0__15__4_, 
        connection_0__15__3_, connection_0__15__2_, connection_0__15__1_, 
        connection_0__15__0_, connection_0__13__31_, connection_0__13__30_, 
        connection_0__13__29_, connection_0__13__28_, connection_0__13__27_, 
        connection_0__13__26_, connection_0__13__25_, connection_0__13__24_, 
        connection_0__13__23_, connection_0__13__22_, connection_0__13__21_, 
        connection_0__13__20_, connection_0__13__19_, connection_0__13__18_, 
        connection_0__13__17_, connection_0__13__16_, connection_0__13__15_, 
        connection_0__13__14_, connection_0__13__13_, connection_0__13__12_, 
        connection_0__13__11_, connection_0__13__10_, connection_0__13__9_, 
        connection_0__13__8_, connection_0__13__7_, connection_0__13__6_, 
        connection_0__13__5_, connection_0__13__4_, connection_0__13__3_, 
        connection_0__13__2_, connection_0__13__1_, connection_0__13__0_}), 
        .o_valid({connection_valid_1__15_, connection_valid_1__14_}), 
        .o_data_bus({connection_1__15__31_, connection_1__15__30_, 
        connection_1__15__29_, connection_1__15__28_, connection_1__15__27_, 
        connection_1__15__26_, connection_1__15__25_, connection_1__15__24_, 
        connection_1__15__23_, connection_1__15__22_, connection_1__15__21_, 
        connection_1__15__20_, connection_1__15__19_, connection_1__15__18_, 
        connection_1__15__17_, connection_1__15__16_, connection_1__15__15_, 
        connection_1__15__14_, connection_1__15__13_, connection_1__15__12_, 
        connection_1__15__11_, connection_1__15__10_, connection_1__15__9_, 
        connection_1__15__8_, connection_1__15__7_, connection_1__15__6_, 
        connection_1__15__5_, connection_1__15__4_, connection_1__15__3_, 
        connection_1__15__2_, connection_1__15__1_, connection_1__15__0_, 
        connection_1__14__31_, connection_1__14__30_, connection_1__14__29_, 
        connection_1__14__28_, connection_1__14__27_, connection_1__14__26_, 
        connection_1__14__25_, connection_1__14__24_, connection_1__14__23_, 
        connection_1__14__22_, connection_1__14__21_, connection_1__14__20_, 
        connection_1__14__19_, connection_1__14__18_, connection_1__14__17_, 
        connection_1__14__16_, connection_1__14__15_, connection_1__14__14_, 
        connection_1__14__13_, connection_1__14__12_, connection_1__14__11_, 
        connection_1__14__10_, connection_1__14__9_, connection_1__14__8_, 
        connection_1__14__7_, connection_1__14__6_, connection_1__14__5_, 
        connection_1__14__4_, connection_1__14__3_, connection_1__14__2_, 
        connection_1__14__1_, connection_1__14__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[81:80]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_40 first_half_stages_1__group_first_half_0__switch_first_half_0__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_1__2_, 
        connection_valid_1__0_}), .i_data_bus({connection_1__2__31_, 
        connection_1__2__30_, connection_1__2__29_, connection_1__2__28_, 
        connection_1__2__27_, connection_1__2__26_, connection_1__2__25_, 
        connection_1__2__24_, connection_1__2__23_, connection_1__2__22_, 
        connection_1__2__21_, connection_1__2__20_, connection_1__2__19_, 
        connection_1__2__18_, connection_1__2__17_, connection_1__2__16_, 
        connection_1__2__15_, connection_1__2__14_, connection_1__2__13_, 
        connection_1__2__12_, connection_1__2__11_, connection_1__2__10_, 
        connection_1__2__9_, connection_1__2__8_, connection_1__2__7_, 
        connection_1__2__6_, connection_1__2__5_, connection_1__2__4_, 
        connection_1__2__3_, connection_1__2__2_, connection_1__2__1_, 
        connection_1__2__0_, connection_1__0__31_, connection_1__0__30_, 
        connection_1__0__29_, connection_1__0__28_, connection_1__0__27_, 
        connection_1__0__26_, connection_1__0__25_, connection_1__0__24_, 
        connection_1__0__23_, connection_1__0__22_, connection_1__0__21_, 
        connection_1__0__20_, connection_1__0__19_, connection_1__0__18_, 
        connection_1__0__17_, connection_1__0__16_, connection_1__0__15_, 
        connection_1__0__14_, connection_1__0__13_, connection_1__0__12_, 
        connection_1__0__11_, connection_1__0__10_, connection_1__0__9_, 
        connection_1__0__8_, connection_1__0__7_, connection_1__0__6_, 
        connection_1__0__5_, connection_1__0__4_, connection_1__0__3_, 
        connection_1__0__2_, connection_1__0__1_, connection_1__0__0_}), 
        .o_valid({connection_valid_2__1_, connection_valid_2__0_}), 
        .o_data_bus({connection_2__1__31_, connection_2__1__30_, 
        connection_2__1__29_, connection_2__1__28_, connection_2__1__27_, 
        connection_2__1__26_, connection_2__1__25_, connection_2__1__24_, 
        connection_2__1__23_, connection_2__1__22_, connection_2__1__21_, 
        connection_2__1__20_, connection_2__1__19_, connection_2__1__18_, 
        connection_2__1__17_, connection_2__1__16_, connection_2__1__15_, 
        connection_2__1__14_, connection_2__1__13_, connection_2__1__12_, 
        connection_2__1__11_, connection_2__1__10_, connection_2__1__9_, 
        connection_2__1__8_, connection_2__1__7_, connection_2__1__6_, 
        connection_2__1__5_, connection_2__1__4_, connection_2__1__3_, 
        connection_2__1__2_, connection_2__1__1_, connection_2__1__0_, 
        connection_2__0__31_, connection_2__0__30_, connection_2__0__29_, 
        connection_2__0__28_, connection_2__0__27_, connection_2__0__26_, 
        connection_2__0__25_, connection_2__0__24_, connection_2__0__23_, 
        connection_2__0__22_, connection_2__0__21_, connection_2__0__20_, 
        connection_2__0__19_, connection_2__0__18_, connection_2__0__17_, 
        connection_2__0__16_, connection_2__0__15_, connection_2__0__14_, 
        connection_2__0__13_, connection_2__0__12_, connection_2__0__11_, 
        connection_2__0__10_, connection_2__0__9_, connection_2__0__8_, 
        connection_2__0__7_, connection_2__0__6_, connection_2__0__5_, 
        connection_2__0__4_, connection_2__0__3_, connection_2__0__2_, 
        connection_2__0__1_, connection_2__0__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[79:78]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_39 first_half_stages_1__group_first_half_0__switch_first_half_1__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_1__6_, 
        connection_valid_1__4_}), .i_data_bus({connection_1__6__31_, 
        connection_1__6__30_, connection_1__6__29_, connection_1__6__28_, 
        connection_1__6__27_, connection_1__6__26_, connection_1__6__25_, 
        connection_1__6__24_, connection_1__6__23_, connection_1__6__22_, 
        connection_1__6__21_, connection_1__6__20_, connection_1__6__19_, 
        connection_1__6__18_, connection_1__6__17_, connection_1__6__16_, 
        connection_1__6__15_, connection_1__6__14_, connection_1__6__13_, 
        connection_1__6__12_, connection_1__6__11_, connection_1__6__10_, 
        connection_1__6__9_, connection_1__6__8_, connection_1__6__7_, 
        connection_1__6__6_, connection_1__6__5_, connection_1__6__4_, 
        connection_1__6__3_, connection_1__6__2_, connection_1__6__1_, 
        connection_1__6__0_, connection_1__4__31_, connection_1__4__30_, 
        connection_1__4__29_, connection_1__4__28_, connection_1__4__27_, 
        connection_1__4__26_, connection_1__4__25_, connection_1__4__24_, 
        connection_1__4__23_, connection_1__4__22_, connection_1__4__21_, 
        connection_1__4__20_, connection_1__4__19_, connection_1__4__18_, 
        connection_1__4__17_, connection_1__4__16_, connection_1__4__15_, 
        connection_1__4__14_, connection_1__4__13_, connection_1__4__12_, 
        connection_1__4__11_, connection_1__4__10_, connection_1__4__9_, 
        connection_1__4__8_, connection_1__4__7_, connection_1__4__6_, 
        connection_1__4__5_, connection_1__4__4_, connection_1__4__3_, 
        connection_1__4__2_, connection_1__4__1_, connection_1__4__0_}), 
        .o_valid({connection_valid_2__3_, connection_valid_2__2_}), 
        .o_data_bus({connection_2__3__31_, connection_2__3__30_, 
        connection_2__3__29_, connection_2__3__28_, connection_2__3__27_, 
        connection_2__3__26_, connection_2__3__25_, connection_2__3__24_, 
        connection_2__3__23_, connection_2__3__22_, connection_2__3__21_, 
        connection_2__3__20_, connection_2__3__19_, connection_2__3__18_, 
        connection_2__3__17_, connection_2__3__16_, connection_2__3__15_, 
        connection_2__3__14_, connection_2__3__13_, connection_2__3__12_, 
        connection_2__3__11_, connection_2__3__10_, connection_2__3__9_, 
        connection_2__3__8_, connection_2__3__7_, connection_2__3__6_, 
        connection_2__3__5_, connection_2__3__4_, connection_2__3__3_, 
        connection_2__3__2_, connection_2__3__1_, connection_2__3__0_, 
        connection_2__2__31_, connection_2__2__30_, connection_2__2__29_, 
        connection_2__2__28_, connection_2__2__27_, connection_2__2__26_, 
        connection_2__2__25_, connection_2__2__24_, connection_2__2__23_, 
        connection_2__2__22_, connection_2__2__21_, connection_2__2__20_, 
        connection_2__2__19_, connection_2__2__18_, connection_2__2__17_, 
        connection_2__2__16_, connection_2__2__15_, connection_2__2__14_, 
        connection_2__2__13_, connection_2__2__12_, connection_2__2__11_, 
        connection_2__2__10_, connection_2__2__9_, connection_2__2__8_, 
        connection_2__2__7_, connection_2__2__6_, connection_2__2__5_, 
        connection_2__2__4_, connection_2__2__3_, connection_2__2__2_, 
        connection_2__2__1_, connection_2__2__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[77:76]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_38 first_half_stages_1__group_first_half_0__switch_first_half_2__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_1__3_, 
        connection_valid_1__1_}), .i_data_bus({connection_1__3__31_, 
        connection_1__3__30_, connection_1__3__29_, connection_1__3__28_, 
        connection_1__3__27_, connection_1__3__26_, connection_1__3__25_, 
        connection_1__3__24_, connection_1__3__23_, connection_1__3__22_, 
        connection_1__3__21_, connection_1__3__20_, connection_1__3__19_, 
        connection_1__3__18_, connection_1__3__17_, connection_1__3__16_, 
        connection_1__3__15_, connection_1__3__14_, connection_1__3__13_, 
        connection_1__3__12_, connection_1__3__11_, connection_1__3__10_, 
        connection_1__3__9_, connection_1__3__8_, connection_1__3__7_, 
        connection_1__3__6_, connection_1__3__5_, connection_1__3__4_, 
        connection_1__3__3_, connection_1__3__2_, connection_1__3__1_, 
        connection_1__3__0_, connection_1__1__31_, connection_1__1__30_, 
        connection_1__1__29_, connection_1__1__28_, connection_1__1__27_, 
        connection_1__1__26_, connection_1__1__25_, connection_1__1__24_, 
        connection_1__1__23_, connection_1__1__22_, connection_1__1__21_, 
        connection_1__1__20_, connection_1__1__19_, connection_1__1__18_, 
        connection_1__1__17_, connection_1__1__16_, connection_1__1__15_, 
        connection_1__1__14_, connection_1__1__13_, connection_1__1__12_, 
        connection_1__1__11_, connection_1__1__10_, connection_1__1__9_, 
        connection_1__1__8_, connection_1__1__7_, connection_1__1__6_, 
        connection_1__1__5_, connection_1__1__4_, connection_1__1__3_, 
        connection_1__1__2_, connection_1__1__1_, connection_1__1__0_}), 
        .o_valid({connection_valid_2__5_, connection_valid_2__4_}), 
        .o_data_bus({connection_2__5__31_, connection_2__5__30_, 
        connection_2__5__29_, connection_2__5__28_, connection_2__5__27_, 
        connection_2__5__26_, connection_2__5__25_, connection_2__5__24_, 
        connection_2__5__23_, connection_2__5__22_, connection_2__5__21_, 
        connection_2__5__20_, connection_2__5__19_, connection_2__5__18_, 
        connection_2__5__17_, connection_2__5__16_, connection_2__5__15_, 
        connection_2__5__14_, connection_2__5__13_, connection_2__5__12_, 
        connection_2__5__11_, connection_2__5__10_, connection_2__5__9_, 
        connection_2__5__8_, connection_2__5__7_, connection_2__5__6_, 
        connection_2__5__5_, connection_2__5__4_, connection_2__5__3_, 
        connection_2__5__2_, connection_2__5__1_, connection_2__5__0_, 
        connection_2__4__31_, connection_2__4__30_, connection_2__4__29_, 
        connection_2__4__28_, connection_2__4__27_, connection_2__4__26_, 
        connection_2__4__25_, connection_2__4__24_, connection_2__4__23_, 
        connection_2__4__22_, connection_2__4__21_, connection_2__4__20_, 
        connection_2__4__19_, connection_2__4__18_, connection_2__4__17_, 
        connection_2__4__16_, connection_2__4__15_, connection_2__4__14_, 
        connection_2__4__13_, connection_2__4__12_, connection_2__4__11_, 
        connection_2__4__10_, connection_2__4__9_, connection_2__4__8_, 
        connection_2__4__7_, connection_2__4__6_, connection_2__4__5_, 
        connection_2__4__4_, connection_2__4__3_, connection_2__4__2_, 
        connection_2__4__1_, connection_2__4__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[75:74]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_37 first_half_stages_1__group_first_half_0__switch_first_half_3__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_1__7_, 
        connection_valid_1__5_}), .i_data_bus({connection_1__7__31_, 
        connection_1__7__30_, connection_1__7__29_, connection_1__7__28_, 
        connection_1__7__27_, connection_1__7__26_, connection_1__7__25_, 
        connection_1__7__24_, connection_1__7__23_, connection_1__7__22_, 
        connection_1__7__21_, connection_1__7__20_, connection_1__7__19_, 
        connection_1__7__18_, connection_1__7__17_, connection_1__7__16_, 
        connection_1__7__15_, connection_1__7__14_, connection_1__7__13_, 
        connection_1__7__12_, connection_1__7__11_, connection_1__7__10_, 
        connection_1__7__9_, connection_1__7__8_, connection_1__7__7_, 
        connection_1__7__6_, connection_1__7__5_, connection_1__7__4_, 
        connection_1__7__3_, connection_1__7__2_, connection_1__7__1_, 
        connection_1__7__0_, connection_1__5__31_, connection_1__5__30_, 
        connection_1__5__29_, connection_1__5__28_, connection_1__5__27_, 
        connection_1__5__26_, connection_1__5__25_, connection_1__5__24_, 
        connection_1__5__23_, connection_1__5__22_, connection_1__5__21_, 
        connection_1__5__20_, connection_1__5__19_, connection_1__5__18_, 
        connection_1__5__17_, connection_1__5__16_, connection_1__5__15_, 
        connection_1__5__14_, connection_1__5__13_, connection_1__5__12_, 
        connection_1__5__11_, connection_1__5__10_, connection_1__5__9_, 
        connection_1__5__8_, connection_1__5__7_, connection_1__5__6_, 
        connection_1__5__5_, connection_1__5__4_, connection_1__5__3_, 
        connection_1__5__2_, connection_1__5__1_, connection_1__5__0_}), 
        .o_valid({connection_valid_2__7_, connection_valid_2__6_}), 
        .o_data_bus({connection_2__7__31_, connection_2__7__30_, 
        connection_2__7__29_, connection_2__7__28_, connection_2__7__27_, 
        connection_2__7__26_, connection_2__7__25_, connection_2__7__24_, 
        connection_2__7__23_, connection_2__7__22_, connection_2__7__21_, 
        connection_2__7__20_, connection_2__7__19_, connection_2__7__18_, 
        connection_2__7__17_, connection_2__7__16_, connection_2__7__15_, 
        connection_2__7__14_, connection_2__7__13_, connection_2__7__12_, 
        connection_2__7__11_, connection_2__7__10_, connection_2__7__9_, 
        connection_2__7__8_, connection_2__7__7_, connection_2__7__6_, 
        connection_2__7__5_, connection_2__7__4_, connection_2__7__3_, 
        connection_2__7__2_, connection_2__7__1_, connection_2__7__0_, 
        connection_2__6__31_, connection_2__6__30_, connection_2__6__29_, 
        connection_2__6__28_, connection_2__6__27_, connection_2__6__26_, 
        connection_2__6__25_, connection_2__6__24_, connection_2__6__23_, 
        connection_2__6__22_, connection_2__6__21_, connection_2__6__20_, 
        connection_2__6__19_, connection_2__6__18_, connection_2__6__17_, 
        connection_2__6__16_, connection_2__6__15_, connection_2__6__14_, 
        connection_2__6__13_, connection_2__6__12_, connection_2__6__11_, 
        connection_2__6__10_, connection_2__6__9_, connection_2__6__8_, 
        connection_2__6__7_, connection_2__6__6_, connection_2__6__5_, 
        connection_2__6__4_, connection_2__6__3_, connection_2__6__2_, 
        connection_2__6__1_, connection_2__6__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[73:72]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_36 first_half_stages_1__group_first_half_1__switch_first_half_0__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_1__10_, 
        connection_valid_1__8_}), .i_data_bus({connection_1__10__31_, 
        connection_1__10__30_, connection_1__10__29_, connection_1__10__28_, 
        connection_1__10__27_, connection_1__10__26_, connection_1__10__25_, 
        connection_1__10__24_, connection_1__10__23_, connection_1__10__22_, 
        connection_1__10__21_, connection_1__10__20_, connection_1__10__19_, 
        connection_1__10__18_, connection_1__10__17_, connection_1__10__16_, 
        connection_1__10__15_, connection_1__10__14_, connection_1__10__13_, 
        connection_1__10__12_, connection_1__10__11_, connection_1__10__10_, 
        connection_1__10__9_, connection_1__10__8_, connection_1__10__7_, 
        connection_1__10__6_, connection_1__10__5_, connection_1__10__4_, 
        connection_1__10__3_, connection_1__10__2_, connection_1__10__1_, 
        connection_1__10__0_, connection_1__8__31_, connection_1__8__30_, 
        connection_1__8__29_, connection_1__8__28_, connection_1__8__27_, 
        connection_1__8__26_, connection_1__8__25_, connection_1__8__24_, 
        connection_1__8__23_, connection_1__8__22_, connection_1__8__21_, 
        connection_1__8__20_, connection_1__8__19_, connection_1__8__18_, 
        connection_1__8__17_, connection_1__8__16_, connection_1__8__15_, 
        connection_1__8__14_, connection_1__8__13_, connection_1__8__12_, 
        connection_1__8__11_, connection_1__8__10_, connection_1__8__9_, 
        connection_1__8__8_, connection_1__8__7_, connection_1__8__6_, 
        connection_1__8__5_, connection_1__8__4_, connection_1__8__3_, 
        connection_1__8__2_, connection_1__8__1_, connection_1__8__0_}), 
        .o_valid({connection_valid_2__9_, connection_valid_2__8_}), 
        .o_data_bus({connection_2__9__31_, connection_2__9__30_, 
        connection_2__9__29_, connection_2__9__28_, connection_2__9__27_, 
        connection_2__9__26_, connection_2__9__25_, connection_2__9__24_, 
        connection_2__9__23_, connection_2__9__22_, connection_2__9__21_, 
        connection_2__9__20_, connection_2__9__19_, connection_2__9__18_, 
        connection_2__9__17_, connection_2__9__16_, connection_2__9__15_, 
        connection_2__9__14_, connection_2__9__13_, connection_2__9__12_, 
        connection_2__9__11_, connection_2__9__10_, connection_2__9__9_, 
        connection_2__9__8_, connection_2__9__7_, connection_2__9__6_, 
        connection_2__9__5_, connection_2__9__4_, connection_2__9__3_, 
        connection_2__9__2_, connection_2__9__1_, connection_2__9__0_, 
        connection_2__8__31_, connection_2__8__30_, connection_2__8__29_, 
        connection_2__8__28_, connection_2__8__27_, connection_2__8__26_, 
        connection_2__8__25_, connection_2__8__24_, connection_2__8__23_, 
        connection_2__8__22_, connection_2__8__21_, connection_2__8__20_, 
        connection_2__8__19_, connection_2__8__18_, connection_2__8__17_, 
        connection_2__8__16_, connection_2__8__15_, connection_2__8__14_, 
        connection_2__8__13_, connection_2__8__12_, connection_2__8__11_, 
        connection_2__8__10_, connection_2__8__9_, connection_2__8__8_, 
        connection_2__8__7_, connection_2__8__6_, connection_2__8__5_, 
        connection_2__8__4_, connection_2__8__3_, connection_2__8__2_, 
        connection_2__8__1_, connection_2__8__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[71:70]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_35 first_half_stages_1__group_first_half_1__switch_first_half_1__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_1__14_, 
        connection_valid_1__12_}), .i_data_bus({connection_1__14__31_, 
        connection_1__14__30_, connection_1__14__29_, connection_1__14__28_, 
        connection_1__14__27_, connection_1__14__26_, connection_1__14__25_, 
        connection_1__14__24_, connection_1__14__23_, connection_1__14__22_, 
        connection_1__14__21_, connection_1__14__20_, connection_1__14__19_, 
        connection_1__14__18_, connection_1__14__17_, connection_1__14__16_, 
        connection_1__14__15_, connection_1__14__14_, connection_1__14__13_, 
        connection_1__14__12_, connection_1__14__11_, connection_1__14__10_, 
        connection_1__14__9_, connection_1__14__8_, connection_1__14__7_, 
        connection_1__14__6_, connection_1__14__5_, connection_1__14__4_, 
        connection_1__14__3_, connection_1__14__2_, connection_1__14__1_, 
        connection_1__14__0_, connection_1__12__31_, connection_1__12__30_, 
        connection_1__12__29_, connection_1__12__28_, connection_1__12__27_, 
        connection_1__12__26_, connection_1__12__25_, connection_1__12__24_, 
        connection_1__12__23_, connection_1__12__22_, connection_1__12__21_, 
        connection_1__12__20_, connection_1__12__19_, connection_1__12__18_, 
        connection_1__12__17_, connection_1__12__16_, connection_1__12__15_, 
        connection_1__12__14_, connection_1__12__13_, connection_1__12__12_, 
        connection_1__12__11_, connection_1__12__10_, connection_1__12__9_, 
        connection_1__12__8_, connection_1__12__7_, connection_1__12__6_, 
        connection_1__12__5_, connection_1__12__4_, connection_1__12__3_, 
        connection_1__12__2_, connection_1__12__1_, connection_1__12__0_}), 
        .o_valid({connection_valid_2__11_, connection_valid_2__10_}), 
        .o_data_bus({connection_2__11__31_, connection_2__11__30_, 
        connection_2__11__29_, connection_2__11__28_, connection_2__11__27_, 
        connection_2__11__26_, connection_2__11__25_, connection_2__11__24_, 
        connection_2__11__23_, connection_2__11__22_, connection_2__11__21_, 
        connection_2__11__20_, connection_2__11__19_, connection_2__11__18_, 
        connection_2__11__17_, connection_2__11__16_, connection_2__11__15_, 
        connection_2__11__14_, connection_2__11__13_, connection_2__11__12_, 
        connection_2__11__11_, connection_2__11__10_, connection_2__11__9_, 
        connection_2__11__8_, connection_2__11__7_, connection_2__11__6_, 
        connection_2__11__5_, connection_2__11__4_, connection_2__11__3_, 
        connection_2__11__2_, connection_2__11__1_, connection_2__11__0_, 
        connection_2__10__31_, connection_2__10__30_, connection_2__10__29_, 
        connection_2__10__28_, connection_2__10__27_, connection_2__10__26_, 
        connection_2__10__25_, connection_2__10__24_, connection_2__10__23_, 
        connection_2__10__22_, connection_2__10__21_, connection_2__10__20_, 
        connection_2__10__19_, connection_2__10__18_, connection_2__10__17_, 
        connection_2__10__16_, connection_2__10__15_, connection_2__10__14_, 
        connection_2__10__13_, connection_2__10__12_, connection_2__10__11_, 
        connection_2__10__10_, connection_2__10__9_, connection_2__10__8_, 
        connection_2__10__7_, connection_2__10__6_, connection_2__10__5_, 
        connection_2__10__4_, connection_2__10__3_, connection_2__10__2_, 
        connection_2__10__1_, connection_2__10__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[69:68]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_34 first_half_stages_1__group_first_half_1__switch_first_half_2__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_1__11_, 
        connection_valid_1__9_}), .i_data_bus({connection_1__11__31_, 
        connection_1__11__30_, connection_1__11__29_, connection_1__11__28_, 
        connection_1__11__27_, connection_1__11__26_, connection_1__11__25_, 
        connection_1__11__24_, connection_1__11__23_, connection_1__11__22_, 
        connection_1__11__21_, connection_1__11__20_, connection_1__11__19_, 
        connection_1__11__18_, connection_1__11__17_, connection_1__11__16_, 
        connection_1__11__15_, connection_1__11__14_, connection_1__11__13_, 
        connection_1__11__12_, connection_1__11__11_, connection_1__11__10_, 
        connection_1__11__9_, connection_1__11__8_, connection_1__11__7_, 
        connection_1__11__6_, connection_1__11__5_, connection_1__11__4_, 
        connection_1__11__3_, connection_1__11__2_, connection_1__11__1_, 
        connection_1__11__0_, connection_1__9__31_, connection_1__9__30_, 
        connection_1__9__29_, connection_1__9__28_, connection_1__9__27_, 
        connection_1__9__26_, connection_1__9__25_, connection_1__9__24_, 
        connection_1__9__23_, connection_1__9__22_, connection_1__9__21_, 
        connection_1__9__20_, connection_1__9__19_, connection_1__9__18_, 
        connection_1__9__17_, connection_1__9__16_, connection_1__9__15_, 
        connection_1__9__14_, connection_1__9__13_, connection_1__9__12_, 
        connection_1__9__11_, connection_1__9__10_, connection_1__9__9_, 
        connection_1__9__8_, connection_1__9__7_, connection_1__9__6_, 
        connection_1__9__5_, connection_1__9__4_, connection_1__9__3_, 
        connection_1__9__2_, connection_1__9__1_, connection_1__9__0_}), 
        .o_valid({connection_valid_2__13_, connection_valid_2__12_}), 
        .o_data_bus({connection_2__13__31_, connection_2__13__30_, 
        connection_2__13__29_, connection_2__13__28_, connection_2__13__27_, 
        connection_2__13__26_, connection_2__13__25_, connection_2__13__24_, 
        connection_2__13__23_, connection_2__13__22_, connection_2__13__21_, 
        connection_2__13__20_, connection_2__13__19_, connection_2__13__18_, 
        connection_2__13__17_, connection_2__13__16_, connection_2__13__15_, 
        connection_2__13__14_, connection_2__13__13_, connection_2__13__12_, 
        connection_2__13__11_, connection_2__13__10_, connection_2__13__9_, 
        connection_2__13__8_, connection_2__13__7_, connection_2__13__6_, 
        connection_2__13__5_, connection_2__13__4_, connection_2__13__3_, 
        connection_2__13__2_, connection_2__13__1_, connection_2__13__0_, 
        connection_2__12__31_, connection_2__12__30_, connection_2__12__29_, 
        connection_2__12__28_, connection_2__12__27_, connection_2__12__26_, 
        connection_2__12__25_, connection_2__12__24_, connection_2__12__23_, 
        connection_2__12__22_, connection_2__12__21_, connection_2__12__20_, 
        connection_2__12__19_, connection_2__12__18_, connection_2__12__17_, 
        connection_2__12__16_, connection_2__12__15_, connection_2__12__14_, 
        connection_2__12__13_, connection_2__12__12_, connection_2__12__11_, 
        connection_2__12__10_, connection_2__12__9_, connection_2__12__8_, 
        connection_2__12__7_, connection_2__12__6_, connection_2__12__5_, 
        connection_2__12__4_, connection_2__12__3_, connection_2__12__2_, 
        connection_2__12__1_, connection_2__12__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[67:66]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_33 first_half_stages_1__group_first_half_1__switch_first_half_3__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_1__15_, 
        connection_valid_1__13_}), .i_data_bus({connection_1__15__31_, 
        connection_1__15__30_, connection_1__15__29_, connection_1__15__28_, 
        connection_1__15__27_, connection_1__15__26_, connection_1__15__25_, 
        connection_1__15__24_, connection_1__15__23_, connection_1__15__22_, 
        connection_1__15__21_, connection_1__15__20_, connection_1__15__19_, 
        connection_1__15__18_, connection_1__15__17_, connection_1__15__16_, 
        connection_1__15__15_, connection_1__15__14_, connection_1__15__13_, 
        connection_1__15__12_, connection_1__15__11_, connection_1__15__10_, 
        connection_1__15__9_, connection_1__15__8_, connection_1__15__7_, 
        connection_1__15__6_, connection_1__15__5_, connection_1__15__4_, 
        connection_1__15__3_, connection_1__15__2_, connection_1__15__1_, 
        connection_1__15__0_, connection_1__13__31_, connection_1__13__30_, 
        connection_1__13__29_, connection_1__13__28_, connection_1__13__27_, 
        connection_1__13__26_, connection_1__13__25_, connection_1__13__24_, 
        connection_1__13__23_, connection_1__13__22_, connection_1__13__21_, 
        connection_1__13__20_, connection_1__13__19_, connection_1__13__18_, 
        connection_1__13__17_, connection_1__13__16_, connection_1__13__15_, 
        connection_1__13__14_, connection_1__13__13_, connection_1__13__12_, 
        connection_1__13__11_, connection_1__13__10_, connection_1__13__9_, 
        connection_1__13__8_, connection_1__13__7_, connection_1__13__6_, 
        connection_1__13__5_, connection_1__13__4_, connection_1__13__3_, 
        connection_1__13__2_, connection_1__13__1_, connection_1__13__0_}), 
        .o_valid({connection_valid_2__15_, connection_valid_2__14_}), 
        .o_data_bus({connection_2__15__31_, connection_2__15__30_, 
        connection_2__15__29_, connection_2__15__28_, connection_2__15__27_, 
        connection_2__15__26_, connection_2__15__25_, connection_2__15__24_, 
        connection_2__15__23_, connection_2__15__22_, connection_2__15__21_, 
        connection_2__15__20_, connection_2__15__19_, connection_2__15__18_, 
        connection_2__15__17_, connection_2__15__16_, connection_2__15__15_, 
        connection_2__15__14_, connection_2__15__13_, connection_2__15__12_, 
        connection_2__15__11_, connection_2__15__10_, connection_2__15__9_, 
        connection_2__15__8_, connection_2__15__7_, connection_2__15__6_, 
        connection_2__15__5_, connection_2__15__4_, connection_2__15__3_, 
        connection_2__15__2_, connection_2__15__1_, connection_2__15__0_, 
        connection_2__14__31_, connection_2__14__30_, connection_2__14__29_, 
        connection_2__14__28_, connection_2__14__27_, connection_2__14__26_, 
        connection_2__14__25_, connection_2__14__24_, connection_2__14__23_, 
        connection_2__14__22_, connection_2__14__21_, connection_2__14__20_, 
        connection_2__14__19_, connection_2__14__18_, connection_2__14__17_, 
        connection_2__14__16_, connection_2__14__15_, connection_2__14__14_, 
        connection_2__14__13_, connection_2__14__12_, connection_2__14__11_, 
        connection_2__14__10_, connection_2__14__9_, connection_2__14__8_, 
        connection_2__14__7_, connection_2__14__6_, connection_2__14__5_, 
        connection_2__14__4_, connection_2__14__3_, connection_2__14__2_, 
        connection_2__14__1_, connection_2__14__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[65:64]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_32 first_half_stages_2__group_first_half_0__switch_first_half_0__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__2_, 
        connection_valid_2__0_}), .i_data_bus({connection_2__2__31_, 
        connection_2__2__30_, connection_2__2__29_, connection_2__2__28_, 
        connection_2__2__27_, connection_2__2__26_, connection_2__2__25_, 
        connection_2__2__24_, connection_2__2__23_, connection_2__2__22_, 
        connection_2__2__21_, connection_2__2__20_, connection_2__2__19_, 
        connection_2__2__18_, connection_2__2__17_, connection_2__2__16_, 
        connection_2__2__15_, connection_2__2__14_, connection_2__2__13_, 
        connection_2__2__12_, connection_2__2__11_, connection_2__2__10_, 
        connection_2__2__9_, connection_2__2__8_, connection_2__2__7_, 
        connection_2__2__6_, connection_2__2__5_, connection_2__2__4_, 
        connection_2__2__3_, connection_2__2__2_, connection_2__2__1_, 
        connection_2__2__0_, connection_2__0__31_, connection_2__0__30_, 
        connection_2__0__29_, connection_2__0__28_, connection_2__0__27_, 
        connection_2__0__26_, connection_2__0__25_, connection_2__0__24_, 
        connection_2__0__23_, connection_2__0__22_, connection_2__0__21_, 
        connection_2__0__20_, connection_2__0__19_, connection_2__0__18_, 
        connection_2__0__17_, connection_2__0__16_, connection_2__0__15_, 
        connection_2__0__14_, connection_2__0__13_, connection_2__0__12_, 
        connection_2__0__11_, connection_2__0__10_, connection_2__0__9_, 
        connection_2__0__8_, connection_2__0__7_, connection_2__0__6_, 
        connection_2__0__5_, connection_2__0__4_, connection_2__0__3_, 
        connection_2__0__2_, connection_2__0__1_, connection_2__0__0_}), 
        .o_valid({connection_valid_3__1_, connection_valid_3__0_}), 
        .o_data_bus({connection_3__1__31_, connection_3__1__30_, 
        connection_3__1__29_, connection_3__1__28_, connection_3__1__27_, 
        connection_3__1__26_, connection_3__1__25_, connection_3__1__24_, 
        connection_3__1__23_, connection_3__1__22_, connection_3__1__21_, 
        connection_3__1__20_, connection_3__1__19_, connection_3__1__18_, 
        connection_3__1__17_, connection_3__1__16_, connection_3__1__15_, 
        connection_3__1__14_, connection_3__1__13_, connection_3__1__12_, 
        connection_3__1__11_, connection_3__1__10_, connection_3__1__9_, 
        connection_3__1__8_, connection_3__1__7_, connection_3__1__6_, 
        connection_3__1__5_, connection_3__1__4_, connection_3__1__3_, 
        connection_3__1__2_, connection_3__1__1_, connection_3__1__0_, 
        connection_3__0__31_, connection_3__0__30_, connection_3__0__29_, 
        connection_3__0__28_, connection_3__0__27_, connection_3__0__26_, 
        connection_3__0__25_, connection_3__0__24_, connection_3__0__23_, 
        connection_3__0__22_, connection_3__0__21_, connection_3__0__20_, 
        connection_3__0__19_, connection_3__0__18_, connection_3__0__17_, 
        connection_3__0__16_, connection_3__0__15_, connection_3__0__14_, 
        connection_3__0__13_, connection_3__0__12_, connection_3__0__11_, 
        connection_3__0__10_, connection_3__0__9_, connection_3__0__8_, 
        connection_3__0__7_, connection_3__0__6_, connection_3__0__5_, 
        connection_3__0__4_, connection_3__0__3_, connection_3__0__2_, 
        connection_3__0__1_, connection_3__0__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[63:62]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_31 first_half_stages_2__group_first_half_0__switch_first_half_1__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__3_, 
        connection_valid_2__1_}), .i_data_bus({connection_2__3__31_, 
        connection_2__3__30_, connection_2__3__29_, connection_2__3__28_, 
        connection_2__3__27_, connection_2__3__26_, connection_2__3__25_, 
        connection_2__3__24_, connection_2__3__23_, connection_2__3__22_, 
        connection_2__3__21_, connection_2__3__20_, connection_2__3__19_, 
        connection_2__3__18_, connection_2__3__17_, connection_2__3__16_, 
        connection_2__3__15_, connection_2__3__14_, connection_2__3__13_, 
        connection_2__3__12_, connection_2__3__11_, connection_2__3__10_, 
        connection_2__3__9_, connection_2__3__8_, connection_2__3__7_, 
        connection_2__3__6_, connection_2__3__5_, connection_2__3__4_, 
        connection_2__3__3_, connection_2__3__2_, connection_2__3__1_, 
        connection_2__3__0_, connection_2__1__31_, connection_2__1__30_, 
        connection_2__1__29_, connection_2__1__28_, connection_2__1__27_, 
        connection_2__1__26_, connection_2__1__25_, connection_2__1__24_, 
        connection_2__1__23_, connection_2__1__22_, connection_2__1__21_, 
        connection_2__1__20_, connection_2__1__19_, connection_2__1__18_, 
        connection_2__1__17_, connection_2__1__16_, connection_2__1__15_, 
        connection_2__1__14_, connection_2__1__13_, connection_2__1__12_, 
        connection_2__1__11_, connection_2__1__10_, connection_2__1__9_, 
        connection_2__1__8_, connection_2__1__7_, connection_2__1__6_, 
        connection_2__1__5_, connection_2__1__4_, connection_2__1__3_, 
        connection_2__1__2_, connection_2__1__1_, connection_2__1__0_}), 
        .o_valid({connection_valid_3__3_, connection_valid_3__2_}), 
        .o_data_bus({connection_3__3__31_, connection_3__3__30_, 
        connection_3__3__29_, connection_3__3__28_, connection_3__3__27_, 
        connection_3__3__26_, connection_3__3__25_, connection_3__3__24_, 
        connection_3__3__23_, connection_3__3__22_, connection_3__3__21_, 
        connection_3__3__20_, connection_3__3__19_, connection_3__3__18_, 
        connection_3__3__17_, connection_3__3__16_, connection_3__3__15_, 
        connection_3__3__14_, connection_3__3__13_, connection_3__3__12_, 
        connection_3__3__11_, connection_3__3__10_, connection_3__3__9_, 
        connection_3__3__8_, connection_3__3__7_, connection_3__3__6_, 
        connection_3__3__5_, connection_3__3__4_, connection_3__3__3_, 
        connection_3__3__2_, connection_3__3__1_, connection_3__3__0_, 
        connection_3__2__31_, connection_3__2__30_, connection_3__2__29_, 
        connection_3__2__28_, connection_3__2__27_, connection_3__2__26_, 
        connection_3__2__25_, connection_3__2__24_, connection_3__2__23_, 
        connection_3__2__22_, connection_3__2__21_, connection_3__2__20_, 
        connection_3__2__19_, connection_3__2__18_, connection_3__2__17_, 
        connection_3__2__16_, connection_3__2__15_, connection_3__2__14_, 
        connection_3__2__13_, connection_3__2__12_, connection_3__2__11_, 
        connection_3__2__10_, connection_3__2__9_, connection_3__2__8_, 
        connection_3__2__7_, connection_3__2__6_, connection_3__2__5_, 
        connection_3__2__4_, connection_3__2__3_, connection_3__2__2_, 
        connection_3__2__1_, connection_3__2__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[61:60]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_30 first_half_stages_2__group_first_half_1__switch_first_half_0__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__6_, 
        connection_valid_2__4_}), .i_data_bus({connection_2__6__31_, 
        connection_2__6__30_, connection_2__6__29_, connection_2__6__28_, 
        connection_2__6__27_, connection_2__6__26_, connection_2__6__25_, 
        connection_2__6__24_, connection_2__6__23_, connection_2__6__22_, 
        connection_2__6__21_, connection_2__6__20_, connection_2__6__19_, 
        connection_2__6__18_, connection_2__6__17_, connection_2__6__16_, 
        connection_2__6__15_, connection_2__6__14_, connection_2__6__13_, 
        connection_2__6__12_, connection_2__6__11_, connection_2__6__10_, 
        connection_2__6__9_, connection_2__6__8_, connection_2__6__7_, 
        connection_2__6__6_, connection_2__6__5_, connection_2__6__4_, 
        connection_2__6__3_, connection_2__6__2_, connection_2__6__1_, 
        connection_2__6__0_, connection_2__4__31_, connection_2__4__30_, 
        connection_2__4__29_, connection_2__4__28_, connection_2__4__27_, 
        connection_2__4__26_, connection_2__4__25_, connection_2__4__24_, 
        connection_2__4__23_, connection_2__4__22_, connection_2__4__21_, 
        connection_2__4__20_, connection_2__4__19_, connection_2__4__18_, 
        connection_2__4__17_, connection_2__4__16_, connection_2__4__15_, 
        connection_2__4__14_, connection_2__4__13_, connection_2__4__12_, 
        connection_2__4__11_, connection_2__4__10_, connection_2__4__9_, 
        connection_2__4__8_, connection_2__4__7_, connection_2__4__6_, 
        connection_2__4__5_, connection_2__4__4_, connection_2__4__3_, 
        connection_2__4__2_, connection_2__4__1_, connection_2__4__0_}), 
        .o_valid({connection_valid_3__5_, connection_valid_3__4_}), 
        .o_data_bus({connection_3__5__31_, connection_3__5__30_, 
        connection_3__5__29_, connection_3__5__28_, connection_3__5__27_, 
        connection_3__5__26_, connection_3__5__25_, connection_3__5__24_, 
        connection_3__5__23_, connection_3__5__22_, connection_3__5__21_, 
        connection_3__5__20_, connection_3__5__19_, connection_3__5__18_, 
        connection_3__5__17_, connection_3__5__16_, connection_3__5__15_, 
        connection_3__5__14_, connection_3__5__13_, connection_3__5__12_, 
        connection_3__5__11_, connection_3__5__10_, connection_3__5__9_, 
        connection_3__5__8_, connection_3__5__7_, connection_3__5__6_, 
        connection_3__5__5_, connection_3__5__4_, connection_3__5__3_, 
        connection_3__5__2_, connection_3__5__1_, connection_3__5__0_, 
        connection_3__4__31_, connection_3__4__30_, connection_3__4__29_, 
        connection_3__4__28_, connection_3__4__27_, connection_3__4__26_, 
        connection_3__4__25_, connection_3__4__24_, connection_3__4__23_, 
        connection_3__4__22_, connection_3__4__21_, connection_3__4__20_, 
        connection_3__4__19_, connection_3__4__18_, connection_3__4__17_, 
        connection_3__4__16_, connection_3__4__15_, connection_3__4__14_, 
        connection_3__4__13_, connection_3__4__12_, connection_3__4__11_, 
        connection_3__4__10_, connection_3__4__9_, connection_3__4__8_, 
        connection_3__4__7_, connection_3__4__6_, connection_3__4__5_, 
        connection_3__4__4_, connection_3__4__3_, connection_3__4__2_, 
        connection_3__4__1_, connection_3__4__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[59:58]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_29 first_half_stages_2__group_first_half_1__switch_first_half_1__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__7_, 
        connection_valid_2__5_}), .i_data_bus({connection_2__7__31_, 
        connection_2__7__30_, connection_2__7__29_, connection_2__7__28_, 
        connection_2__7__27_, connection_2__7__26_, connection_2__7__25_, 
        connection_2__7__24_, connection_2__7__23_, connection_2__7__22_, 
        connection_2__7__21_, connection_2__7__20_, connection_2__7__19_, 
        connection_2__7__18_, connection_2__7__17_, connection_2__7__16_, 
        connection_2__7__15_, connection_2__7__14_, connection_2__7__13_, 
        connection_2__7__12_, connection_2__7__11_, connection_2__7__10_, 
        connection_2__7__9_, connection_2__7__8_, connection_2__7__7_, 
        connection_2__7__6_, connection_2__7__5_, connection_2__7__4_, 
        connection_2__7__3_, connection_2__7__2_, connection_2__7__1_, 
        connection_2__7__0_, connection_2__5__31_, connection_2__5__30_, 
        connection_2__5__29_, connection_2__5__28_, connection_2__5__27_, 
        connection_2__5__26_, connection_2__5__25_, connection_2__5__24_, 
        connection_2__5__23_, connection_2__5__22_, connection_2__5__21_, 
        connection_2__5__20_, connection_2__5__19_, connection_2__5__18_, 
        connection_2__5__17_, connection_2__5__16_, connection_2__5__15_, 
        connection_2__5__14_, connection_2__5__13_, connection_2__5__12_, 
        connection_2__5__11_, connection_2__5__10_, connection_2__5__9_, 
        connection_2__5__8_, connection_2__5__7_, connection_2__5__6_, 
        connection_2__5__5_, connection_2__5__4_, connection_2__5__3_, 
        connection_2__5__2_, connection_2__5__1_, connection_2__5__0_}), 
        .o_valid({connection_valid_3__7_, connection_valid_3__6_}), 
        .o_data_bus({connection_3__7__31_, connection_3__7__30_, 
        connection_3__7__29_, connection_3__7__28_, connection_3__7__27_, 
        connection_3__7__26_, connection_3__7__25_, connection_3__7__24_, 
        connection_3__7__23_, connection_3__7__22_, connection_3__7__21_, 
        connection_3__7__20_, connection_3__7__19_, connection_3__7__18_, 
        connection_3__7__17_, connection_3__7__16_, connection_3__7__15_, 
        connection_3__7__14_, connection_3__7__13_, connection_3__7__12_, 
        connection_3__7__11_, connection_3__7__10_, connection_3__7__9_, 
        connection_3__7__8_, connection_3__7__7_, connection_3__7__6_, 
        connection_3__7__5_, connection_3__7__4_, connection_3__7__3_, 
        connection_3__7__2_, connection_3__7__1_, connection_3__7__0_, 
        connection_3__6__31_, connection_3__6__30_, connection_3__6__29_, 
        connection_3__6__28_, connection_3__6__27_, connection_3__6__26_, 
        connection_3__6__25_, connection_3__6__24_, connection_3__6__23_, 
        connection_3__6__22_, connection_3__6__21_, connection_3__6__20_, 
        connection_3__6__19_, connection_3__6__18_, connection_3__6__17_, 
        connection_3__6__16_, connection_3__6__15_, connection_3__6__14_, 
        connection_3__6__13_, connection_3__6__12_, connection_3__6__11_, 
        connection_3__6__10_, connection_3__6__9_, connection_3__6__8_, 
        connection_3__6__7_, connection_3__6__6_, connection_3__6__5_, 
        connection_3__6__4_, connection_3__6__3_, connection_3__6__2_, 
        connection_3__6__1_, connection_3__6__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[57:56]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_28 first_half_stages_2__group_first_half_2__switch_first_half_0__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__10_, 
        connection_valid_2__8_}), .i_data_bus({connection_2__10__31_, 
        connection_2__10__30_, connection_2__10__29_, connection_2__10__28_, 
        connection_2__10__27_, connection_2__10__26_, connection_2__10__25_, 
        connection_2__10__24_, connection_2__10__23_, connection_2__10__22_, 
        connection_2__10__21_, connection_2__10__20_, connection_2__10__19_, 
        connection_2__10__18_, connection_2__10__17_, connection_2__10__16_, 
        connection_2__10__15_, connection_2__10__14_, connection_2__10__13_, 
        connection_2__10__12_, connection_2__10__11_, connection_2__10__10_, 
        connection_2__10__9_, connection_2__10__8_, connection_2__10__7_, 
        connection_2__10__6_, connection_2__10__5_, connection_2__10__4_, 
        connection_2__10__3_, connection_2__10__2_, connection_2__10__1_, 
        connection_2__10__0_, connection_2__8__31_, connection_2__8__30_, 
        connection_2__8__29_, connection_2__8__28_, connection_2__8__27_, 
        connection_2__8__26_, connection_2__8__25_, connection_2__8__24_, 
        connection_2__8__23_, connection_2__8__22_, connection_2__8__21_, 
        connection_2__8__20_, connection_2__8__19_, connection_2__8__18_, 
        connection_2__8__17_, connection_2__8__16_, connection_2__8__15_, 
        connection_2__8__14_, connection_2__8__13_, connection_2__8__12_, 
        connection_2__8__11_, connection_2__8__10_, connection_2__8__9_, 
        connection_2__8__8_, connection_2__8__7_, connection_2__8__6_, 
        connection_2__8__5_, connection_2__8__4_, connection_2__8__3_, 
        connection_2__8__2_, connection_2__8__1_, connection_2__8__0_}), 
        .o_valid({connection_valid_3__9_, connection_valid_3__8_}), 
        .o_data_bus({connection_3__9__31_, connection_3__9__30_, 
        connection_3__9__29_, connection_3__9__28_, connection_3__9__27_, 
        connection_3__9__26_, connection_3__9__25_, connection_3__9__24_, 
        connection_3__9__23_, connection_3__9__22_, connection_3__9__21_, 
        connection_3__9__20_, connection_3__9__19_, connection_3__9__18_, 
        connection_3__9__17_, connection_3__9__16_, connection_3__9__15_, 
        connection_3__9__14_, connection_3__9__13_, connection_3__9__12_, 
        connection_3__9__11_, connection_3__9__10_, connection_3__9__9_, 
        connection_3__9__8_, connection_3__9__7_, connection_3__9__6_, 
        connection_3__9__5_, connection_3__9__4_, connection_3__9__3_, 
        connection_3__9__2_, connection_3__9__1_, connection_3__9__0_, 
        connection_3__8__31_, connection_3__8__30_, connection_3__8__29_, 
        connection_3__8__28_, connection_3__8__27_, connection_3__8__26_, 
        connection_3__8__25_, connection_3__8__24_, connection_3__8__23_, 
        connection_3__8__22_, connection_3__8__21_, connection_3__8__20_, 
        connection_3__8__19_, connection_3__8__18_, connection_3__8__17_, 
        connection_3__8__16_, connection_3__8__15_, connection_3__8__14_, 
        connection_3__8__13_, connection_3__8__12_, connection_3__8__11_, 
        connection_3__8__10_, connection_3__8__9_, connection_3__8__8_, 
        connection_3__8__7_, connection_3__8__6_, connection_3__8__5_, 
        connection_3__8__4_, connection_3__8__3_, connection_3__8__2_, 
        connection_3__8__1_, connection_3__8__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[55:54]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_27 first_half_stages_2__group_first_half_2__switch_first_half_1__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__11_, 
        connection_valid_2__9_}), .i_data_bus({connection_2__11__31_, 
        connection_2__11__30_, connection_2__11__29_, connection_2__11__28_, 
        connection_2__11__27_, connection_2__11__26_, connection_2__11__25_, 
        connection_2__11__24_, connection_2__11__23_, connection_2__11__22_, 
        connection_2__11__21_, connection_2__11__20_, connection_2__11__19_, 
        connection_2__11__18_, connection_2__11__17_, connection_2__11__16_, 
        connection_2__11__15_, connection_2__11__14_, connection_2__11__13_, 
        connection_2__11__12_, connection_2__11__11_, connection_2__11__10_, 
        connection_2__11__9_, connection_2__11__8_, connection_2__11__7_, 
        connection_2__11__6_, connection_2__11__5_, connection_2__11__4_, 
        connection_2__11__3_, connection_2__11__2_, connection_2__11__1_, 
        connection_2__11__0_, connection_2__9__31_, connection_2__9__30_, 
        connection_2__9__29_, connection_2__9__28_, connection_2__9__27_, 
        connection_2__9__26_, connection_2__9__25_, connection_2__9__24_, 
        connection_2__9__23_, connection_2__9__22_, connection_2__9__21_, 
        connection_2__9__20_, connection_2__9__19_, connection_2__9__18_, 
        connection_2__9__17_, connection_2__9__16_, connection_2__9__15_, 
        connection_2__9__14_, connection_2__9__13_, connection_2__9__12_, 
        connection_2__9__11_, connection_2__9__10_, connection_2__9__9_, 
        connection_2__9__8_, connection_2__9__7_, connection_2__9__6_, 
        connection_2__9__5_, connection_2__9__4_, connection_2__9__3_, 
        connection_2__9__2_, connection_2__9__1_, connection_2__9__0_}), 
        .o_valid({connection_valid_3__11_, connection_valid_3__10_}), 
        .o_data_bus({connection_3__11__31_, connection_3__11__30_, 
        connection_3__11__29_, connection_3__11__28_, connection_3__11__27_, 
        connection_3__11__26_, connection_3__11__25_, connection_3__11__24_, 
        connection_3__11__23_, connection_3__11__22_, connection_3__11__21_, 
        connection_3__11__20_, connection_3__11__19_, connection_3__11__18_, 
        connection_3__11__17_, connection_3__11__16_, connection_3__11__15_, 
        connection_3__11__14_, connection_3__11__13_, connection_3__11__12_, 
        connection_3__11__11_, connection_3__11__10_, connection_3__11__9_, 
        connection_3__11__8_, connection_3__11__7_, connection_3__11__6_, 
        connection_3__11__5_, connection_3__11__4_, connection_3__11__3_, 
        connection_3__11__2_, connection_3__11__1_, connection_3__11__0_, 
        connection_3__10__31_, connection_3__10__30_, connection_3__10__29_, 
        connection_3__10__28_, connection_3__10__27_, connection_3__10__26_, 
        connection_3__10__25_, connection_3__10__24_, connection_3__10__23_, 
        connection_3__10__22_, connection_3__10__21_, connection_3__10__20_, 
        connection_3__10__19_, connection_3__10__18_, connection_3__10__17_, 
        connection_3__10__16_, connection_3__10__15_, connection_3__10__14_, 
        connection_3__10__13_, connection_3__10__12_, connection_3__10__11_, 
        connection_3__10__10_, connection_3__10__9_, connection_3__10__8_, 
        connection_3__10__7_, connection_3__10__6_, connection_3__10__5_, 
        connection_3__10__4_, connection_3__10__3_, connection_3__10__2_, 
        connection_3__10__1_, connection_3__10__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[53:52]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_26 first_half_stages_2__group_first_half_3__switch_first_half_0__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__14_, 
        connection_valid_2__12_}), .i_data_bus({connection_2__14__31_, 
        connection_2__14__30_, connection_2__14__29_, connection_2__14__28_, 
        connection_2__14__27_, connection_2__14__26_, connection_2__14__25_, 
        connection_2__14__24_, connection_2__14__23_, connection_2__14__22_, 
        connection_2__14__21_, connection_2__14__20_, connection_2__14__19_, 
        connection_2__14__18_, connection_2__14__17_, connection_2__14__16_, 
        connection_2__14__15_, connection_2__14__14_, connection_2__14__13_, 
        connection_2__14__12_, connection_2__14__11_, connection_2__14__10_, 
        connection_2__14__9_, connection_2__14__8_, connection_2__14__7_, 
        connection_2__14__6_, connection_2__14__5_, connection_2__14__4_, 
        connection_2__14__3_, connection_2__14__2_, connection_2__14__1_, 
        connection_2__14__0_, connection_2__12__31_, connection_2__12__30_, 
        connection_2__12__29_, connection_2__12__28_, connection_2__12__27_, 
        connection_2__12__26_, connection_2__12__25_, connection_2__12__24_, 
        connection_2__12__23_, connection_2__12__22_, connection_2__12__21_, 
        connection_2__12__20_, connection_2__12__19_, connection_2__12__18_, 
        connection_2__12__17_, connection_2__12__16_, connection_2__12__15_, 
        connection_2__12__14_, connection_2__12__13_, connection_2__12__12_, 
        connection_2__12__11_, connection_2__12__10_, connection_2__12__9_, 
        connection_2__12__8_, connection_2__12__7_, connection_2__12__6_, 
        connection_2__12__5_, connection_2__12__4_, connection_2__12__3_, 
        connection_2__12__2_, connection_2__12__1_, connection_2__12__0_}), 
        .o_valid({connection_valid_3__13_, connection_valid_3__12_}), 
        .o_data_bus({connection_3__13__31_, connection_3__13__30_, 
        connection_3__13__29_, connection_3__13__28_, connection_3__13__27_, 
        connection_3__13__26_, connection_3__13__25_, connection_3__13__24_, 
        connection_3__13__23_, connection_3__13__22_, connection_3__13__21_, 
        connection_3__13__20_, connection_3__13__19_, connection_3__13__18_, 
        connection_3__13__17_, connection_3__13__16_, connection_3__13__15_, 
        connection_3__13__14_, connection_3__13__13_, connection_3__13__12_, 
        connection_3__13__11_, connection_3__13__10_, connection_3__13__9_, 
        connection_3__13__8_, connection_3__13__7_, connection_3__13__6_, 
        connection_3__13__5_, connection_3__13__4_, connection_3__13__3_, 
        connection_3__13__2_, connection_3__13__1_, connection_3__13__0_, 
        connection_3__12__31_, connection_3__12__30_, connection_3__12__29_, 
        connection_3__12__28_, connection_3__12__27_, connection_3__12__26_, 
        connection_3__12__25_, connection_3__12__24_, connection_3__12__23_, 
        connection_3__12__22_, connection_3__12__21_, connection_3__12__20_, 
        connection_3__12__19_, connection_3__12__18_, connection_3__12__17_, 
        connection_3__12__16_, connection_3__12__15_, connection_3__12__14_, 
        connection_3__12__13_, connection_3__12__12_, connection_3__12__11_, 
        connection_3__12__10_, connection_3__12__9_, connection_3__12__8_, 
        connection_3__12__7_, connection_3__12__6_, connection_3__12__5_, 
        connection_3__12__4_, connection_3__12__3_, connection_3__12__2_, 
        connection_3__12__1_, connection_3__12__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[51:50]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_25 first_half_stages_2__group_first_half_3__switch_first_half_1__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__15_, 
        connection_valid_2__13_}), .i_data_bus({connection_2__15__31_, 
        connection_2__15__30_, connection_2__15__29_, connection_2__15__28_, 
        connection_2__15__27_, connection_2__15__26_, connection_2__15__25_, 
        connection_2__15__24_, connection_2__15__23_, connection_2__15__22_, 
        connection_2__15__21_, connection_2__15__20_, connection_2__15__19_, 
        connection_2__15__18_, connection_2__15__17_, connection_2__15__16_, 
        connection_2__15__15_, connection_2__15__14_, connection_2__15__13_, 
        connection_2__15__12_, connection_2__15__11_, connection_2__15__10_, 
        connection_2__15__9_, connection_2__15__8_, connection_2__15__7_, 
        connection_2__15__6_, connection_2__15__5_, connection_2__15__4_, 
        connection_2__15__3_, connection_2__15__2_, connection_2__15__1_, 
        connection_2__15__0_, connection_2__13__31_, connection_2__13__30_, 
        connection_2__13__29_, connection_2__13__28_, connection_2__13__27_, 
        connection_2__13__26_, connection_2__13__25_, connection_2__13__24_, 
        connection_2__13__23_, connection_2__13__22_, connection_2__13__21_, 
        connection_2__13__20_, connection_2__13__19_, connection_2__13__18_, 
        connection_2__13__17_, connection_2__13__16_, connection_2__13__15_, 
        connection_2__13__14_, connection_2__13__13_, connection_2__13__12_, 
        connection_2__13__11_, connection_2__13__10_, connection_2__13__9_, 
        connection_2__13__8_, connection_2__13__7_, connection_2__13__6_, 
        connection_2__13__5_, connection_2__13__4_, connection_2__13__3_, 
        connection_2__13__2_, connection_2__13__1_, connection_2__13__0_}), 
        .o_valid({connection_valid_3__15_, connection_valid_3__14_}), 
        .o_data_bus({connection_3__15__31_, connection_3__15__30_, 
        connection_3__15__29_, connection_3__15__28_, connection_3__15__27_, 
        connection_3__15__26_, connection_3__15__25_, connection_3__15__24_, 
        connection_3__15__23_, connection_3__15__22_, connection_3__15__21_, 
        connection_3__15__20_, connection_3__15__19_, connection_3__15__18_, 
        connection_3__15__17_, connection_3__15__16_, connection_3__15__15_, 
        connection_3__15__14_, connection_3__15__13_, connection_3__15__12_, 
        connection_3__15__11_, connection_3__15__10_, connection_3__15__9_, 
        connection_3__15__8_, connection_3__15__7_, connection_3__15__6_, 
        connection_3__15__5_, connection_3__15__4_, connection_3__15__3_, 
        connection_3__15__2_, connection_3__15__1_, connection_3__15__0_, 
        connection_3__14__31_, connection_3__14__30_, connection_3__14__29_, 
        connection_3__14__28_, connection_3__14__27_, connection_3__14__26_, 
        connection_3__14__25_, connection_3__14__24_, connection_3__14__23_, 
        connection_3__14__22_, connection_3__14__21_, connection_3__14__20_, 
        connection_3__14__19_, connection_3__14__18_, connection_3__14__17_, 
        connection_3__14__16_, connection_3__14__15_, connection_3__14__14_, 
        connection_3__14__13_, connection_3__14__12_, connection_3__14__11_, 
        connection_3__14__10_, connection_3__14__9_, connection_3__14__8_, 
        connection_3__14__7_, connection_3__14__6_, connection_3__14__5_, 
        connection_3__14__4_, connection_3__14__3_, connection_3__14__2_, 
        connection_3__14__1_, connection_3__14__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[49:48]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_24 second_half_stages_3__group_sec_half_0__switch_sec_half_0__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__2_, 
        connection_valid_3__0_}), .i_data_bus({connection_3__2__31_, 
        connection_3__2__30_, connection_3__2__29_, connection_3__2__28_, 
        connection_3__2__27_, connection_3__2__26_, connection_3__2__25_, 
        connection_3__2__24_, connection_3__2__23_, connection_3__2__22_, 
        connection_3__2__21_, connection_3__2__20_, connection_3__2__19_, 
        connection_3__2__18_, connection_3__2__17_, connection_3__2__16_, 
        connection_3__2__15_, connection_3__2__14_, connection_3__2__13_, 
        connection_3__2__12_, connection_3__2__11_, connection_3__2__10_, 
        connection_3__2__9_, connection_3__2__8_, connection_3__2__7_, 
        connection_3__2__6_, connection_3__2__5_, connection_3__2__4_, 
        connection_3__2__3_, connection_3__2__2_, connection_3__2__1_, 
        connection_3__2__0_, connection_3__0__31_, connection_3__0__30_, 
        connection_3__0__29_, connection_3__0__28_, connection_3__0__27_, 
        connection_3__0__26_, connection_3__0__25_, connection_3__0__24_, 
        connection_3__0__23_, connection_3__0__22_, connection_3__0__21_, 
        connection_3__0__20_, connection_3__0__19_, connection_3__0__18_, 
        connection_3__0__17_, connection_3__0__16_, connection_3__0__15_, 
        connection_3__0__14_, connection_3__0__13_, connection_3__0__12_, 
        connection_3__0__11_, connection_3__0__10_, connection_3__0__9_, 
        connection_3__0__8_, connection_3__0__7_, connection_3__0__6_, 
        connection_3__0__5_, connection_3__0__4_, connection_3__0__3_, 
        connection_3__0__2_, connection_3__0__1_, connection_3__0__0_}), 
        .o_valid({connection_valid_4__1_, connection_valid_4__0_}), 
        .o_data_bus({connection_4__1__31_, connection_4__1__30_, 
        connection_4__1__29_, connection_4__1__28_, connection_4__1__27_, 
        connection_4__1__26_, connection_4__1__25_, connection_4__1__24_, 
        connection_4__1__23_, connection_4__1__22_, connection_4__1__21_, 
        connection_4__1__20_, connection_4__1__19_, connection_4__1__18_, 
        connection_4__1__17_, connection_4__1__16_, connection_4__1__15_, 
        connection_4__1__14_, connection_4__1__13_, connection_4__1__12_, 
        connection_4__1__11_, connection_4__1__10_, connection_4__1__9_, 
        connection_4__1__8_, connection_4__1__7_, connection_4__1__6_, 
        connection_4__1__5_, connection_4__1__4_, connection_4__1__3_, 
        connection_4__1__2_, connection_4__1__1_, connection_4__1__0_, 
        connection_4__0__31_, connection_4__0__30_, connection_4__0__29_, 
        connection_4__0__28_, connection_4__0__27_, connection_4__0__26_, 
        connection_4__0__25_, connection_4__0__24_, connection_4__0__23_, 
        connection_4__0__22_, connection_4__0__21_, connection_4__0__20_, 
        connection_4__0__19_, connection_4__0__18_, connection_4__0__17_, 
        connection_4__0__16_, connection_4__0__15_, connection_4__0__14_, 
        connection_4__0__13_, connection_4__0__12_, connection_4__0__11_, 
        connection_4__0__10_, connection_4__0__9_, connection_4__0__8_, 
        connection_4__0__7_, connection_4__0__6_, connection_4__0__5_, 
        connection_4__0__4_, connection_4__0__3_, connection_4__0__2_, 
        connection_4__0__1_, connection_4__0__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[47:46]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_23 second_half_stages_3__group_sec_half_0__switch_sec_half_1__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__3_, 
        connection_valid_3__1_}), .i_data_bus({connection_3__3__31_, 
        connection_3__3__30_, connection_3__3__29_, connection_3__3__28_, 
        connection_3__3__27_, connection_3__3__26_, connection_3__3__25_, 
        connection_3__3__24_, connection_3__3__23_, connection_3__3__22_, 
        connection_3__3__21_, connection_3__3__20_, connection_3__3__19_, 
        connection_3__3__18_, connection_3__3__17_, connection_3__3__16_, 
        connection_3__3__15_, connection_3__3__14_, connection_3__3__13_, 
        connection_3__3__12_, connection_3__3__11_, connection_3__3__10_, 
        connection_3__3__9_, connection_3__3__8_, connection_3__3__7_, 
        connection_3__3__6_, connection_3__3__5_, connection_3__3__4_, 
        connection_3__3__3_, connection_3__3__2_, connection_3__3__1_, 
        connection_3__3__0_, connection_3__1__31_, connection_3__1__30_, 
        connection_3__1__29_, connection_3__1__28_, connection_3__1__27_, 
        connection_3__1__26_, connection_3__1__25_, connection_3__1__24_, 
        connection_3__1__23_, connection_3__1__22_, connection_3__1__21_, 
        connection_3__1__20_, connection_3__1__19_, connection_3__1__18_, 
        connection_3__1__17_, connection_3__1__16_, connection_3__1__15_, 
        connection_3__1__14_, connection_3__1__13_, connection_3__1__12_, 
        connection_3__1__11_, connection_3__1__10_, connection_3__1__9_, 
        connection_3__1__8_, connection_3__1__7_, connection_3__1__6_, 
        connection_3__1__5_, connection_3__1__4_, connection_3__1__3_, 
        connection_3__1__2_, connection_3__1__1_, connection_3__1__0_}), 
        .o_valid({connection_valid_4__3_, connection_valid_4__2_}), 
        .o_data_bus({connection_4__3__31_, connection_4__3__30_, 
        connection_4__3__29_, connection_4__3__28_, connection_4__3__27_, 
        connection_4__3__26_, connection_4__3__25_, connection_4__3__24_, 
        connection_4__3__23_, connection_4__3__22_, connection_4__3__21_, 
        connection_4__3__20_, connection_4__3__19_, connection_4__3__18_, 
        connection_4__3__17_, connection_4__3__16_, connection_4__3__15_, 
        connection_4__3__14_, connection_4__3__13_, connection_4__3__12_, 
        connection_4__3__11_, connection_4__3__10_, connection_4__3__9_, 
        connection_4__3__8_, connection_4__3__7_, connection_4__3__6_, 
        connection_4__3__5_, connection_4__3__4_, connection_4__3__3_, 
        connection_4__3__2_, connection_4__3__1_, connection_4__3__0_, 
        connection_4__2__31_, connection_4__2__30_, connection_4__2__29_, 
        connection_4__2__28_, connection_4__2__27_, connection_4__2__26_, 
        connection_4__2__25_, connection_4__2__24_, connection_4__2__23_, 
        connection_4__2__22_, connection_4__2__21_, connection_4__2__20_, 
        connection_4__2__19_, connection_4__2__18_, connection_4__2__17_, 
        connection_4__2__16_, connection_4__2__15_, connection_4__2__14_, 
        connection_4__2__13_, connection_4__2__12_, connection_4__2__11_, 
        connection_4__2__10_, connection_4__2__9_, connection_4__2__8_, 
        connection_4__2__7_, connection_4__2__6_, connection_4__2__5_, 
        connection_4__2__4_, connection_4__2__3_, connection_4__2__2_, 
        connection_4__2__1_, connection_4__2__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[45:44]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_22 second_half_stages_3__group_sec_half_1__switch_sec_half_0__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__6_, 
        connection_valid_3__4_}), .i_data_bus({connection_3__6__31_, 
        connection_3__6__30_, connection_3__6__29_, connection_3__6__28_, 
        connection_3__6__27_, connection_3__6__26_, connection_3__6__25_, 
        connection_3__6__24_, connection_3__6__23_, connection_3__6__22_, 
        connection_3__6__21_, connection_3__6__20_, connection_3__6__19_, 
        connection_3__6__18_, connection_3__6__17_, connection_3__6__16_, 
        connection_3__6__15_, connection_3__6__14_, connection_3__6__13_, 
        connection_3__6__12_, connection_3__6__11_, connection_3__6__10_, 
        connection_3__6__9_, connection_3__6__8_, connection_3__6__7_, 
        connection_3__6__6_, connection_3__6__5_, connection_3__6__4_, 
        connection_3__6__3_, connection_3__6__2_, connection_3__6__1_, 
        connection_3__6__0_, connection_3__4__31_, connection_3__4__30_, 
        connection_3__4__29_, connection_3__4__28_, connection_3__4__27_, 
        connection_3__4__26_, connection_3__4__25_, connection_3__4__24_, 
        connection_3__4__23_, connection_3__4__22_, connection_3__4__21_, 
        connection_3__4__20_, connection_3__4__19_, connection_3__4__18_, 
        connection_3__4__17_, connection_3__4__16_, connection_3__4__15_, 
        connection_3__4__14_, connection_3__4__13_, connection_3__4__12_, 
        connection_3__4__11_, connection_3__4__10_, connection_3__4__9_, 
        connection_3__4__8_, connection_3__4__7_, connection_3__4__6_, 
        connection_3__4__5_, connection_3__4__4_, connection_3__4__3_, 
        connection_3__4__2_, connection_3__4__1_, connection_3__4__0_}), 
        .o_valid({connection_valid_4__5_, connection_valid_4__4_}), 
        .o_data_bus({connection_4__5__31_, connection_4__5__30_, 
        connection_4__5__29_, connection_4__5__28_, connection_4__5__27_, 
        connection_4__5__26_, connection_4__5__25_, connection_4__5__24_, 
        connection_4__5__23_, connection_4__5__22_, connection_4__5__21_, 
        connection_4__5__20_, connection_4__5__19_, connection_4__5__18_, 
        connection_4__5__17_, connection_4__5__16_, connection_4__5__15_, 
        connection_4__5__14_, connection_4__5__13_, connection_4__5__12_, 
        connection_4__5__11_, connection_4__5__10_, connection_4__5__9_, 
        connection_4__5__8_, connection_4__5__7_, connection_4__5__6_, 
        connection_4__5__5_, connection_4__5__4_, connection_4__5__3_, 
        connection_4__5__2_, connection_4__5__1_, connection_4__5__0_, 
        connection_4__4__31_, connection_4__4__30_, connection_4__4__29_, 
        connection_4__4__28_, connection_4__4__27_, connection_4__4__26_, 
        connection_4__4__25_, connection_4__4__24_, connection_4__4__23_, 
        connection_4__4__22_, connection_4__4__21_, connection_4__4__20_, 
        connection_4__4__19_, connection_4__4__18_, connection_4__4__17_, 
        connection_4__4__16_, connection_4__4__15_, connection_4__4__14_, 
        connection_4__4__13_, connection_4__4__12_, connection_4__4__11_, 
        connection_4__4__10_, connection_4__4__9_, connection_4__4__8_, 
        connection_4__4__7_, connection_4__4__6_, connection_4__4__5_, 
        connection_4__4__4_, connection_4__4__3_, connection_4__4__2_, 
        connection_4__4__1_, connection_4__4__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[43:42]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_21 second_half_stages_3__group_sec_half_1__switch_sec_half_1__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__7_, 
        connection_valid_3__5_}), .i_data_bus({connection_3__7__31_, 
        connection_3__7__30_, connection_3__7__29_, connection_3__7__28_, 
        connection_3__7__27_, connection_3__7__26_, connection_3__7__25_, 
        connection_3__7__24_, connection_3__7__23_, connection_3__7__22_, 
        connection_3__7__21_, connection_3__7__20_, connection_3__7__19_, 
        connection_3__7__18_, connection_3__7__17_, connection_3__7__16_, 
        connection_3__7__15_, connection_3__7__14_, connection_3__7__13_, 
        connection_3__7__12_, connection_3__7__11_, connection_3__7__10_, 
        connection_3__7__9_, connection_3__7__8_, connection_3__7__7_, 
        connection_3__7__6_, connection_3__7__5_, connection_3__7__4_, 
        connection_3__7__3_, connection_3__7__2_, connection_3__7__1_, 
        connection_3__7__0_, connection_3__5__31_, connection_3__5__30_, 
        connection_3__5__29_, connection_3__5__28_, connection_3__5__27_, 
        connection_3__5__26_, connection_3__5__25_, connection_3__5__24_, 
        connection_3__5__23_, connection_3__5__22_, connection_3__5__21_, 
        connection_3__5__20_, connection_3__5__19_, connection_3__5__18_, 
        connection_3__5__17_, connection_3__5__16_, connection_3__5__15_, 
        connection_3__5__14_, connection_3__5__13_, connection_3__5__12_, 
        connection_3__5__11_, connection_3__5__10_, connection_3__5__9_, 
        connection_3__5__8_, connection_3__5__7_, connection_3__5__6_, 
        connection_3__5__5_, connection_3__5__4_, connection_3__5__3_, 
        connection_3__5__2_, connection_3__5__1_, connection_3__5__0_}), 
        .o_valid({connection_valid_4__7_, connection_valid_4__6_}), 
        .o_data_bus({connection_4__7__31_, connection_4__7__30_, 
        connection_4__7__29_, connection_4__7__28_, connection_4__7__27_, 
        connection_4__7__26_, connection_4__7__25_, connection_4__7__24_, 
        connection_4__7__23_, connection_4__7__22_, connection_4__7__21_, 
        connection_4__7__20_, connection_4__7__19_, connection_4__7__18_, 
        connection_4__7__17_, connection_4__7__16_, connection_4__7__15_, 
        connection_4__7__14_, connection_4__7__13_, connection_4__7__12_, 
        connection_4__7__11_, connection_4__7__10_, connection_4__7__9_, 
        connection_4__7__8_, connection_4__7__7_, connection_4__7__6_, 
        connection_4__7__5_, connection_4__7__4_, connection_4__7__3_, 
        connection_4__7__2_, connection_4__7__1_, connection_4__7__0_, 
        connection_4__6__31_, connection_4__6__30_, connection_4__6__29_, 
        connection_4__6__28_, connection_4__6__27_, connection_4__6__26_, 
        connection_4__6__25_, connection_4__6__24_, connection_4__6__23_, 
        connection_4__6__22_, connection_4__6__21_, connection_4__6__20_, 
        connection_4__6__19_, connection_4__6__18_, connection_4__6__17_, 
        connection_4__6__16_, connection_4__6__15_, connection_4__6__14_, 
        connection_4__6__13_, connection_4__6__12_, connection_4__6__11_, 
        connection_4__6__10_, connection_4__6__9_, connection_4__6__8_, 
        connection_4__6__7_, connection_4__6__6_, connection_4__6__5_, 
        connection_4__6__4_, connection_4__6__3_, connection_4__6__2_, 
        connection_4__6__1_, connection_4__6__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[41:40]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_20 second_half_stages_3__group_sec_half_2__switch_sec_half_0__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__10_, 
        connection_valid_3__8_}), .i_data_bus({connection_3__10__31_, 
        connection_3__10__30_, connection_3__10__29_, connection_3__10__28_, 
        connection_3__10__27_, connection_3__10__26_, connection_3__10__25_, 
        connection_3__10__24_, connection_3__10__23_, connection_3__10__22_, 
        connection_3__10__21_, connection_3__10__20_, connection_3__10__19_, 
        connection_3__10__18_, connection_3__10__17_, connection_3__10__16_, 
        connection_3__10__15_, connection_3__10__14_, connection_3__10__13_, 
        connection_3__10__12_, connection_3__10__11_, connection_3__10__10_, 
        connection_3__10__9_, connection_3__10__8_, connection_3__10__7_, 
        connection_3__10__6_, connection_3__10__5_, connection_3__10__4_, 
        connection_3__10__3_, connection_3__10__2_, connection_3__10__1_, 
        connection_3__10__0_, connection_3__8__31_, connection_3__8__30_, 
        connection_3__8__29_, connection_3__8__28_, connection_3__8__27_, 
        connection_3__8__26_, connection_3__8__25_, connection_3__8__24_, 
        connection_3__8__23_, connection_3__8__22_, connection_3__8__21_, 
        connection_3__8__20_, connection_3__8__19_, connection_3__8__18_, 
        connection_3__8__17_, connection_3__8__16_, connection_3__8__15_, 
        connection_3__8__14_, connection_3__8__13_, connection_3__8__12_, 
        connection_3__8__11_, connection_3__8__10_, connection_3__8__9_, 
        connection_3__8__8_, connection_3__8__7_, connection_3__8__6_, 
        connection_3__8__5_, connection_3__8__4_, connection_3__8__3_, 
        connection_3__8__2_, connection_3__8__1_, connection_3__8__0_}), 
        .o_valid({connection_valid_4__9_, connection_valid_4__8_}), 
        .o_data_bus({connection_4__9__31_, connection_4__9__30_, 
        connection_4__9__29_, connection_4__9__28_, connection_4__9__27_, 
        connection_4__9__26_, connection_4__9__25_, connection_4__9__24_, 
        connection_4__9__23_, connection_4__9__22_, connection_4__9__21_, 
        connection_4__9__20_, connection_4__9__19_, connection_4__9__18_, 
        connection_4__9__17_, connection_4__9__16_, connection_4__9__15_, 
        connection_4__9__14_, connection_4__9__13_, connection_4__9__12_, 
        connection_4__9__11_, connection_4__9__10_, connection_4__9__9_, 
        connection_4__9__8_, connection_4__9__7_, connection_4__9__6_, 
        connection_4__9__5_, connection_4__9__4_, connection_4__9__3_, 
        connection_4__9__2_, connection_4__9__1_, connection_4__9__0_, 
        connection_4__8__31_, connection_4__8__30_, connection_4__8__29_, 
        connection_4__8__28_, connection_4__8__27_, connection_4__8__26_, 
        connection_4__8__25_, connection_4__8__24_, connection_4__8__23_, 
        connection_4__8__22_, connection_4__8__21_, connection_4__8__20_, 
        connection_4__8__19_, connection_4__8__18_, connection_4__8__17_, 
        connection_4__8__16_, connection_4__8__15_, connection_4__8__14_, 
        connection_4__8__13_, connection_4__8__12_, connection_4__8__11_, 
        connection_4__8__10_, connection_4__8__9_, connection_4__8__8_, 
        connection_4__8__7_, connection_4__8__6_, connection_4__8__5_, 
        connection_4__8__4_, connection_4__8__3_, connection_4__8__2_, 
        connection_4__8__1_, connection_4__8__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[39:38]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_19 second_half_stages_3__group_sec_half_2__switch_sec_half_1__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__11_, 
        connection_valid_3__9_}), .i_data_bus({connection_3__11__31_, 
        connection_3__11__30_, connection_3__11__29_, connection_3__11__28_, 
        connection_3__11__27_, connection_3__11__26_, connection_3__11__25_, 
        connection_3__11__24_, connection_3__11__23_, connection_3__11__22_, 
        connection_3__11__21_, connection_3__11__20_, connection_3__11__19_, 
        connection_3__11__18_, connection_3__11__17_, connection_3__11__16_, 
        connection_3__11__15_, connection_3__11__14_, connection_3__11__13_, 
        connection_3__11__12_, connection_3__11__11_, connection_3__11__10_, 
        connection_3__11__9_, connection_3__11__8_, connection_3__11__7_, 
        connection_3__11__6_, connection_3__11__5_, connection_3__11__4_, 
        connection_3__11__3_, connection_3__11__2_, connection_3__11__1_, 
        connection_3__11__0_, connection_3__9__31_, connection_3__9__30_, 
        connection_3__9__29_, connection_3__9__28_, connection_3__9__27_, 
        connection_3__9__26_, connection_3__9__25_, connection_3__9__24_, 
        connection_3__9__23_, connection_3__9__22_, connection_3__9__21_, 
        connection_3__9__20_, connection_3__9__19_, connection_3__9__18_, 
        connection_3__9__17_, connection_3__9__16_, connection_3__9__15_, 
        connection_3__9__14_, connection_3__9__13_, connection_3__9__12_, 
        connection_3__9__11_, connection_3__9__10_, connection_3__9__9_, 
        connection_3__9__8_, connection_3__9__7_, connection_3__9__6_, 
        connection_3__9__5_, connection_3__9__4_, connection_3__9__3_, 
        connection_3__9__2_, connection_3__9__1_, connection_3__9__0_}), 
        .o_valid({connection_valid_4__11_, connection_valid_4__10_}), 
        .o_data_bus({connection_4__11__31_, connection_4__11__30_, 
        connection_4__11__29_, connection_4__11__28_, connection_4__11__27_, 
        connection_4__11__26_, connection_4__11__25_, connection_4__11__24_, 
        connection_4__11__23_, connection_4__11__22_, connection_4__11__21_, 
        connection_4__11__20_, connection_4__11__19_, connection_4__11__18_, 
        connection_4__11__17_, connection_4__11__16_, connection_4__11__15_, 
        connection_4__11__14_, connection_4__11__13_, connection_4__11__12_, 
        connection_4__11__11_, connection_4__11__10_, connection_4__11__9_, 
        connection_4__11__8_, connection_4__11__7_, connection_4__11__6_, 
        connection_4__11__5_, connection_4__11__4_, connection_4__11__3_, 
        connection_4__11__2_, connection_4__11__1_, connection_4__11__0_, 
        connection_4__10__31_, connection_4__10__30_, connection_4__10__29_, 
        connection_4__10__28_, connection_4__10__27_, connection_4__10__26_, 
        connection_4__10__25_, connection_4__10__24_, connection_4__10__23_, 
        connection_4__10__22_, connection_4__10__21_, connection_4__10__20_, 
        connection_4__10__19_, connection_4__10__18_, connection_4__10__17_, 
        connection_4__10__16_, connection_4__10__15_, connection_4__10__14_, 
        connection_4__10__13_, connection_4__10__12_, connection_4__10__11_, 
        connection_4__10__10_, connection_4__10__9_, connection_4__10__8_, 
        connection_4__10__7_, connection_4__10__6_, connection_4__10__5_, 
        connection_4__10__4_, connection_4__10__3_, connection_4__10__2_, 
        connection_4__10__1_, connection_4__10__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[37:36]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_18 second_half_stages_3__group_sec_half_3__switch_sec_half_0__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__14_, 
        connection_valid_3__12_}), .i_data_bus({connection_3__14__31_, 
        connection_3__14__30_, connection_3__14__29_, connection_3__14__28_, 
        connection_3__14__27_, connection_3__14__26_, connection_3__14__25_, 
        connection_3__14__24_, connection_3__14__23_, connection_3__14__22_, 
        connection_3__14__21_, connection_3__14__20_, connection_3__14__19_, 
        connection_3__14__18_, connection_3__14__17_, connection_3__14__16_, 
        connection_3__14__15_, connection_3__14__14_, connection_3__14__13_, 
        connection_3__14__12_, connection_3__14__11_, connection_3__14__10_, 
        connection_3__14__9_, connection_3__14__8_, connection_3__14__7_, 
        connection_3__14__6_, connection_3__14__5_, connection_3__14__4_, 
        connection_3__14__3_, connection_3__14__2_, connection_3__14__1_, 
        connection_3__14__0_, connection_3__12__31_, connection_3__12__30_, 
        connection_3__12__29_, connection_3__12__28_, connection_3__12__27_, 
        connection_3__12__26_, connection_3__12__25_, connection_3__12__24_, 
        connection_3__12__23_, connection_3__12__22_, connection_3__12__21_, 
        connection_3__12__20_, connection_3__12__19_, connection_3__12__18_, 
        connection_3__12__17_, connection_3__12__16_, connection_3__12__15_, 
        connection_3__12__14_, connection_3__12__13_, connection_3__12__12_, 
        connection_3__12__11_, connection_3__12__10_, connection_3__12__9_, 
        connection_3__12__8_, connection_3__12__7_, connection_3__12__6_, 
        connection_3__12__5_, connection_3__12__4_, connection_3__12__3_, 
        connection_3__12__2_, connection_3__12__1_, connection_3__12__0_}), 
        .o_valid({connection_valid_4__13_, connection_valid_4__12_}), 
        .o_data_bus({connection_4__13__31_, connection_4__13__30_, 
        connection_4__13__29_, connection_4__13__28_, connection_4__13__27_, 
        connection_4__13__26_, connection_4__13__25_, connection_4__13__24_, 
        connection_4__13__23_, connection_4__13__22_, connection_4__13__21_, 
        connection_4__13__20_, connection_4__13__19_, connection_4__13__18_, 
        connection_4__13__17_, connection_4__13__16_, connection_4__13__15_, 
        connection_4__13__14_, connection_4__13__13_, connection_4__13__12_, 
        connection_4__13__11_, connection_4__13__10_, connection_4__13__9_, 
        connection_4__13__8_, connection_4__13__7_, connection_4__13__6_, 
        connection_4__13__5_, connection_4__13__4_, connection_4__13__3_, 
        connection_4__13__2_, connection_4__13__1_, connection_4__13__0_, 
        connection_4__12__31_, connection_4__12__30_, connection_4__12__29_, 
        connection_4__12__28_, connection_4__12__27_, connection_4__12__26_, 
        connection_4__12__25_, connection_4__12__24_, connection_4__12__23_, 
        connection_4__12__22_, connection_4__12__21_, connection_4__12__20_, 
        connection_4__12__19_, connection_4__12__18_, connection_4__12__17_, 
        connection_4__12__16_, connection_4__12__15_, connection_4__12__14_, 
        connection_4__12__13_, connection_4__12__12_, connection_4__12__11_, 
        connection_4__12__10_, connection_4__12__9_, connection_4__12__8_, 
        connection_4__12__7_, connection_4__12__6_, connection_4__12__5_, 
        connection_4__12__4_, connection_4__12__3_, connection_4__12__2_, 
        connection_4__12__1_, connection_4__12__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[35:34]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_17 second_half_stages_3__group_sec_half_3__switch_sec_half_1__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__15_, 
        connection_valid_3__13_}), .i_data_bus({connection_3__15__31_, 
        connection_3__15__30_, connection_3__15__29_, connection_3__15__28_, 
        connection_3__15__27_, connection_3__15__26_, connection_3__15__25_, 
        connection_3__15__24_, connection_3__15__23_, connection_3__15__22_, 
        connection_3__15__21_, connection_3__15__20_, connection_3__15__19_, 
        connection_3__15__18_, connection_3__15__17_, connection_3__15__16_, 
        connection_3__15__15_, connection_3__15__14_, connection_3__15__13_, 
        connection_3__15__12_, connection_3__15__11_, connection_3__15__10_, 
        connection_3__15__9_, connection_3__15__8_, connection_3__15__7_, 
        connection_3__15__6_, connection_3__15__5_, connection_3__15__4_, 
        connection_3__15__3_, connection_3__15__2_, connection_3__15__1_, 
        connection_3__15__0_, connection_3__13__31_, connection_3__13__30_, 
        connection_3__13__29_, connection_3__13__28_, connection_3__13__27_, 
        connection_3__13__26_, connection_3__13__25_, connection_3__13__24_, 
        connection_3__13__23_, connection_3__13__22_, connection_3__13__21_, 
        connection_3__13__20_, connection_3__13__19_, connection_3__13__18_, 
        connection_3__13__17_, connection_3__13__16_, connection_3__13__15_, 
        connection_3__13__14_, connection_3__13__13_, connection_3__13__12_, 
        connection_3__13__11_, connection_3__13__10_, connection_3__13__9_, 
        connection_3__13__8_, connection_3__13__7_, connection_3__13__6_, 
        connection_3__13__5_, connection_3__13__4_, connection_3__13__3_, 
        connection_3__13__2_, connection_3__13__1_, connection_3__13__0_}), 
        .o_valid({connection_valid_4__15_, connection_valid_4__14_}), 
        .o_data_bus({connection_4__15__31_, connection_4__15__30_, 
        connection_4__15__29_, connection_4__15__28_, connection_4__15__27_, 
        connection_4__15__26_, connection_4__15__25_, connection_4__15__24_, 
        connection_4__15__23_, connection_4__15__22_, connection_4__15__21_, 
        connection_4__15__20_, connection_4__15__19_, connection_4__15__18_, 
        connection_4__15__17_, connection_4__15__16_, connection_4__15__15_, 
        connection_4__15__14_, connection_4__15__13_, connection_4__15__12_, 
        connection_4__15__11_, connection_4__15__10_, connection_4__15__9_, 
        connection_4__15__8_, connection_4__15__7_, connection_4__15__6_, 
        connection_4__15__5_, connection_4__15__4_, connection_4__15__3_, 
        connection_4__15__2_, connection_4__15__1_, connection_4__15__0_, 
        connection_4__14__31_, connection_4__14__30_, connection_4__14__29_, 
        connection_4__14__28_, connection_4__14__27_, connection_4__14__26_, 
        connection_4__14__25_, connection_4__14__24_, connection_4__14__23_, 
        connection_4__14__22_, connection_4__14__21_, connection_4__14__20_, 
        connection_4__14__19_, connection_4__14__18_, connection_4__14__17_, 
        connection_4__14__16_, connection_4__14__15_, connection_4__14__14_, 
        connection_4__14__13_, connection_4__14__12_, connection_4__14__11_, 
        connection_4__14__10_, connection_4__14__9_, connection_4__14__8_, 
        connection_4__14__7_, connection_4__14__6_, connection_4__14__5_, 
        connection_4__14__4_, connection_4__14__3_, connection_4__14__2_, 
        connection_4__14__1_, connection_4__14__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[33:32]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_16 second_half_stages_4__group_sec_half_0__switch_sec_half_0__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__4_, 
        connection_valid_4__0_}), .i_data_bus({connection_4__4__31_, 
        connection_4__4__30_, connection_4__4__29_, connection_4__4__28_, 
        connection_4__4__27_, connection_4__4__26_, connection_4__4__25_, 
        connection_4__4__24_, connection_4__4__23_, connection_4__4__22_, 
        connection_4__4__21_, connection_4__4__20_, connection_4__4__19_, 
        connection_4__4__18_, connection_4__4__17_, connection_4__4__16_, 
        connection_4__4__15_, connection_4__4__14_, connection_4__4__13_, 
        connection_4__4__12_, connection_4__4__11_, connection_4__4__10_, 
        connection_4__4__9_, connection_4__4__8_, connection_4__4__7_, 
        connection_4__4__6_, connection_4__4__5_, connection_4__4__4_, 
        connection_4__4__3_, connection_4__4__2_, connection_4__4__1_, 
        connection_4__4__0_, connection_4__0__31_, connection_4__0__30_, 
        connection_4__0__29_, connection_4__0__28_, connection_4__0__27_, 
        connection_4__0__26_, connection_4__0__25_, connection_4__0__24_, 
        connection_4__0__23_, connection_4__0__22_, connection_4__0__21_, 
        connection_4__0__20_, connection_4__0__19_, connection_4__0__18_, 
        connection_4__0__17_, connection_4__0__16_, connection_4__0__15_, 
        connection_4__0__14_, connection_4__0__13_, connection_4__0__12_, 
        connection_4__0__11_, connection_4__0__10_, connection_4__0__9_, 
        connection_4__0__8_, connection_4__0__7_, connection_4__0__6_, 
        connection_4__0__5_, connection_4__0__4_, connection_4__0__3_, 
        connection_4__0__2_, connection_4__0__1_, connection_4__0__0_}), 
        .o_valid({connection_valid_5__1_, connection_valid_5__0_}), 
        .o_data_bus({connection_5__1__31_, connection_5__1__30_, 
        connection_5__1__29_, connection_5__1__28_, connection_5__1__27_, 
        connection_5__1__26_, connection_5__1__25_, connection_5__1__24_, 
        connection_5__1__23_, connection_5__1__22_, connection_5__1__21_, 
        connection_5__1__20_, connection_5__1__19_, connection_5__1__18_, 
        connection_5__1__17_, connection_5__1__16_, connection_5__1__15_, 
        connection_5__1__14_, connection_5__1__13_, connection_5__1__12_, 
        connection_5__1__11_, connection_5__1__10_, connection_5__1__9_, 
        connection_5__1__8_, connection_5__1__7_, connection_5__1__6_, 
        connection_5__1__5_, connection_5__1__4_, connection_5__1__3_, 
        connection_5__1__2_, connection_5__1__1_, connection_5__1__0_, 
        connection_5__0__31_, connection_5__0__30_, connection_5__0__29_, 
        connection_5__0__28_, connection_5__0__27_, connection_5__0__26_, 
        connection_5__0__25_, connection_5__0__24_, connection_5__0__23_, 
        connection_5__0__22_, connection_5__0__21_, connection_5__0__20_, 
        connection_5__0__19_, connection_5__0__18_, connection_5__0__17_, 
        connection_5__0__16_, connection_5__0__15_, connection_5__0__14_, 
        connection_5__0__13_, connection_5__0__12_, connection_5__0__11_, 
        connection_5__0__10_, connection_5__0__9_, connection_5__0__8_, 
        connection_5__0__7_, connection_5__0__6_, connection_5__0__5_, 
        connection_5__0__4_, connection_5__0__3_, connection_5__0__2_, 
        connection_5__0__1_, connection_5__0__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[31:30]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_15 second_half_stages_4__group_sec_half_0__switch_sec_half_1__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__5_, 
        connection_valid_4__1_}), .i_data_bus({connection_4__5__31_, 
        connection_4__5__30_, connection_4__5__29_, connection_4__5__28_, 
        connection_4__5__27_, connection_4__5__26_, connection_4__5__25_, 
        connection_4__5__24_, connection_4__5__23_, connection_4__5__22_, 
        connection_4__5__21_, connection_4__5__20_, connection_4__5__19_, 
        connection_4__5__18_, connection_4__5__17_, connection_4__5__16_, 
        connection_4__5__15_, connection_4__5__14_, connection_4__5__13_, 
        connection_4__5__12_, connection_4__5__11_, connection_4__5__10_, 
        connection_4__5__9_, connection_4__5__8_, connection_4__5__7_, 
        connection_4__5__6_, connection_4__5__5_, connection_4__5__4_, 
        connection_4__5__3_, connection_4__5__2_, connection_4__5__1_, 
        connection_4__5__0_, connection_4__1__31_, connection_4__1__30_, 
        connection_4__1__29_, connection_4__1__28_, connection_4__1__27_, 
        connection_4__1__26_, connection_4__1__25_, connection_4__1__24_, 
        connection_4__1__23_, connection_4__1__22_, connection_4__1__21_, 
        connection_4__1__20_, connection_4__1__19_, connection_4__1__18_, 
        connection_4__1__17_, connection_4__1__16_, connection_4__1__15_, 
        connection_4__1__14_, connection_4__1__13_, connection_4__1__12_, 
        connection_4__1__11_, connection_4__1__10_, connection_4__1__9_, 
        connection_4__1__8_, connection_4__1__7_, connection_4__1__6_, 
        connection_4__1__5_, connection_4__1__4_, connection_4__1__3_, 
        connection_4__1__2_, connection_4__1__1_, connection_4__1__0_}), 
        .o_valid({connection_valid_5__3_, connection_valid_5__2_}), 
        .o_data_bus({connection_5__3__31_, connection_5__3__30_, 
        connection_5__3__29_, connection_5__3__28_, connection_5__3__27_, 
        connection_5__3__26_, connection_5__3__25_, connection_5__3__24_, 
        connection_5__3__23_, connection_5__3__22_, connection_5__3__21_, 
        connection_5__3__20_, connection_5__3__19_, connection_5__3__18_, 
        connection_5__3__17_, connection_5__3__16_, connection_5__3__15_, 
        connection_5__3__14_, connection_5__3__13_, connection_5__3__12_, 
        connection_5__3__11_, connection_5__3__10_, connection_5__3__9_, 
        connection_5__3__8_, connection_5__3__7_, connection_5__3__6_, 
        connection_5__3__5_, connection_5__3__4_, connection_5__3__3_, 
        connection_5__3__2_, connection_5__3__1_, connection_5__3__0_, 
        connection_5__2__31_, connection_5__2__30_, connection_5__2__29_, 
        connection_5__2__28_, connection_5__2__27_, connection_5__2__26_, 
        connection_5__2__25_, connection_5__2__24_, connection_5__2__23_, 
        connection_5__2__22_, connection_5__2__21_, connection_5__2__20_, 
        connection_5__2__19_, connection_5__2__18_, connection_5__2__17_, 
        connection_5__2__16_, connection_5__2__15_, connection_5__2__14_, 
        connection_5__2__13_, connection_5__2__12_, connection_5__2__11_, 
        connection_5__2__10_, connection_5__2__9_, connection_5__2__8_, 
        connection_5__2__7_, connection_5__2__6_, connection_5__2__5_, 
        connection_5__2__4_, connection_5__2__3_, connection_5__2__2_, 
        connection_5__2__1_, connection_5__2__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[29:28]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_14 second_half_stages_4__group_sec_half_0__switch_sec_half_2__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__6_, 
        connection_valid_4__2_}), .i_data_bus({connection_4__6__31_, 
        connection_4__6__30_, connection_4__6__29_, connection_4__6__28_, 
        connection_4__6__27_, connection_4__6__26_, connection_4__6__25_, 
        connection_4__6__24_, connection_4__6__23_, connection_4__6__22_, 
        connection_4__6__21_, connection_4__6__20_, connection_4__6__19_, 
        connection_4__6__18_, connection_4__6__17_, connection_4__6__16_, 
        connection_4__6__15_, connection_4__6__14_, connection_4__6__13_, 
        connection_4__6__12_, connection_4__6__11_, connection_4__6__10_, 
        connection_4__6__9_, connection_4__6__8_, connection_4__6__7_, 
        connection_4__6__6_, connection_4__6__5_, connection_4__6__4_, 
        connection_4__6__3_, connection_4__6__2_, connection_4__6__1_, 
        connection_4__6__0_, connection_4__2__31_, connection_4__2__30_, 
        connection_4__2__29_, connection_4__2__28_, connection_4__2__27_, 
        connection_4__2__26_, connection_4__2__25_, connection_4__2__24_, 
        connection_4__2__23_, connection_4__2__22_, connection_4__2__21_, 
        connection_4__2__20_, connection_4__2__19_, connection_4__2__18_, 
        connection_4__2__17_, connection_4__2__16_, connection_4__2__15_, 
        connection_4__2__14_, connection_4__2__13_, connection_4__2__12_, 
        connection_4__2__11_, connection_4__2__10_, connection_4__2__9_, 
        connection_4__2__8_, connection_4__2__7_, connection_4__2__6_, 
        connection_4__2__5_, connection_4__2__4_, connection_4__2__3_, 
        connection_4__2__2_, connection_4__2__1_, connection_4__2__0_}), 
        .o_valid({connection_valid_5__5_, connection_valid_5__4_}), 
        .o_data_bus({connection_5__5__31_, connection_5__5__30_, 
        connection_5__5__29_, connection_5__5__28_, connection_5__5__27_, 
        connection_5__5__26_, connection_5__5__25_, connection_5__5__24_, 
        connection_5__5__23_, connection_5__5__22_, connection_5__5__21_, 
        connection_5__5__20_, connection_5__5__19_, connection_5__5__18_, 
        connection_5__5__17_, connection_5__5__16_, connection_5__5__15_, 
        connection_5__5__14_, connection_5__5__13_, connection_5__5__12_, 
        connection_5__5__11_, connection_5__5__10_, connection_5__5__9_, 
        connection_5__5__8_, connection_5__5__7_, connection_5__5__6_, 
        connection_5__5__5_, connection_5__5__4_, connection_5__5__3_, 
        connection_5__5__2_, connection_5__5__1_, connection_5__5__0_, 
        connection_5__4__31_, connection_5__4__30_, connection_5__4__29_, 
        connection_5__4__28_, connection_5__4__27_, connection_5__4__26_, 
        connection_5__4__25_, connection_5__4__24_, connection_5__4__23_, 
        connection_5__4__22_, connection_5__4__21_, connection_5__4__20_, 
        connection_5__4__19_, connection_5__4__18_, connection_5__4__17_, 
        connection_5__4__16_, connection_5__4__15_, connection_5__4__14_, 
        connection_5__4__13_, connection_5__4__12_, connection_5__4__11_, 
        connection_5__4__10_, connection_5__4__9_, connection_5__4__8_, 
        connection_5__4__7_, connection_5__4__6_, connection_5__4__5_, 
        connection_5__4__4_, connection_5__4__3_, connection_5__4__2_, 
        connection_5__4__1_, connection_5__4__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[27:26]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_13 second_half_stages_4__group_sec_half_0__switch_sec_half_3__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__7_, 
        connection_valid_4__3_}), .i_data_bus({connection_4__7__31_, 
        connection_4__7__30_, connection_4__7__29_, connection_4__7__28_, 
        connection_4__7__27_, connection_4__7__26_, connection_4__7__25_, 
        connection_4__7__24_, connection_4__7__23_, connection_4__7__22_, 
        connection_4__7__21_, connection_4__7__20_, connection_4__7__19_, 
        connection_4__7__18_, connection_4__7__17_, connection_4__7__16_, 
        connection_4__7__15_, connection_4__7__14_, connection_4__7__13_, 
        connection_4__7__12_, connection_4__7__11_, connection_4__7__10_, 
        connection_4__7__9_, connection_4__7__8_, connection_4__7__7_, 
        connection_4__7__6_, connection_4__7__5_, connection_4__7__4_, 
        connection_4__7__3_, connection_4__7__2_, connection_4__7__1_, 
        connection_4__7__0_, connection_4__3__31_, connection_4__3__30_, 
        connection_4__3__29_, connection_4__3__28_, connection_4__3__27_, 
        connection_4__3__26_, connection_4__3__25_, connection_4__3__24_, 
        connection_4__3__23_, connection_4__3__22_, connection_4__3__21_, 
        connection_4__3__20_, connection_4__3__19_, connection_4__3__18_, 
        connection_4__3__17_, connection_4__3__16_, connection_4__3__15_, 
        connection_4__3__14_, connection_4__3__13_, connection_4__3__12_, 
        connection_4__3__11_, connection_4__3__10_, connection_4__3__9_, 
        connection_4__3__8_, connection_4__3__7_, connection_4__3__6_, 
        connection_4__3__5_, connection_4__3__4_, connection_4__3__3_, 
        connection_4__3__2_, connection_4__3__1_, connection_4__3__0_}), 
        .o_valid({connection_valid_5__7_, connection_valid_5__6_}), 
        .o_data_bus({connection_5__7__31_, connection_5__7__30_, 
        connection_5__7__29_, connection_5__7__28_, connection_5__7__27_, 
        connection_5__7__26_, connection_5__7__25_, connection_5__7__24_, 
        connection_5__7__23_, connection_5__7__22_, connection_5__7__21_, 
        connection_5__7__20_, connection_5__7__19_, connection_5__7__18_, 
        connection_5__7__17_, connection_5__7__16_, connection_5__7__15_, 
        connection_5__7__14_, connection_5__7__13_, connection_5__7__12_, 
        connection_5__7__11_, connection_5__7__10_, connection_5__7__9_, 
        connection_5__7__8_, connection_5__7__7_, connection_5__7__6_, 
        connection_5__7__5_, connection_5__7__4_, connection_5__7__3_, 
        connection_5__7__2_, connection_5__7__1_, connection_5__7__0_, 
        connection_5__6__31_, connection_5__6__30_, connection_5__6__29_, 
        connection_5__6__28_, connection_5__6__27_, connection_5__6__26_, 
        connection_5__6__25_, connection_5__6__24_, connection_5__6__23_, 
        connection_5__6__22_, connection_5__6__21_, connection_5__6__20_, 
        connection_5__6__19_, connection_5__6__18_, connection_5__6__17_, 
        connection_5__6__16_, connection_5__6__15_, connection_5__6__14_, 
        connection_5__6__13_, connection_5__6__12_, connection_5__6__11_, 
        connection_5__6__10_, connection_5__6__9_, connection_5__6__8_, 
        connection_5__6__7_, connection_5__6__6_, connection_5__6__5_, 
        connection_5__6__4_, connection_5__6__3_, connection_5__6__2_, 
        connection_5__6__1_, connection_5__6__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[25:24]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_12 second_half_stages_4__group_sec_half_1__switch_sec_half_0__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__12_, 
        connection_valid_4__8_}), .i_data_bus({connection_4__12__31_, 
        connection_4__12__30_, connection_4__12__29_, connection_4__12__28_, 
        connection_4__12__27_, connection_4__12__26_, connection_4__12__25_, 
        connection_4__12__24_, connection_4__12__23_, connection_4__12__22_, 
        connection_4__12__21_, connection_4__12__20_, connection_4__12__19_, 
        connection_4__12__18_, connection_4__12__17_, connection_4__12__16_, 
        connection_4__12__15_, connection_4__12__14_, connection_4__12__13_, 
        connection_4__12__12_, connection_4__12__11_, connection_4__12__10_, 
        connection_4__12__9_, connection_4__12__8_, connection_4__12__7_, 
        connection_4__12__6_, connection_4__12__5_, connection_4__12__4_, 
        connection_4__12__3_, connection_4__12__2_, connection_4__12__1_, 
        connection_4__12__0_, connection_4__8__31_, connection_4__8__30_, 
        connection_4__8__29_, connection_4__8__28_, connection_4__8__27_, 
        connection_4__8__26_, connection_4__8__25_, connection_4__8__24_, 
        connection_4__8__23_, connection_4__8__22_, connection_4__8__21_, 
        connection_4__8__20_, connection_4__8__19_, connection_4__8__18_, 
        connection_4__8__17_, connection_4__8__16_, connection_4__8__15_, 
        connection_4__8__14_, connection_4__8__13_, connection_4__8__12_, 
        connection_4__8__11_, connection_4__8__10_, connection_4__8__9_, 
        connection_4__8__8_, connection_4__8__7_, connection_4__8__6_, 
        connection_4__8__5_, connection_4__8__4_, connection_4__8__3_, 
        connection_4__8__2_, connection_4__8__1_, connection_4__8__0_}), 
        .o_valid({connection_valid_5__9_, connection_valid_5__8_}), 
        .o_data_bus({connection_5__9__31_, connection_5__9__30_, 
        connection_5__9__29_, connection_5__9__28_, connection_5__9__27_, 
        connection_5__9__26_, connection_5__9__25_, connection_5__9__24_, 
        connection_5__9__23_, connection_5__9__22_, connection_5__9__21_, 
        connection_5__9__20_, connection_5__9__19_, connection_5__9__18_, 
        connection_5__9__17_, connection_5__9__16_, connection_5__9__15_, 
        connection_5__9__14_, connection_5__9__13_, connection_5__9__12_, 
        connection_5__9__11_, connection_5__9__10_, connection_5__9__9_, 
        connection_5__9__8_, connection_5__9__7_, connection_5__9__6_, 
        connection_5__9__5_, connection_5__9__4_, connection_5__9__3_, 
        connection_5__9__2_, connection_5__9__1_, connection_5__9__0_, 
        connection_5__8__31_, connection_5__8__30_, connection_5__8__29_, 
        connection_5__8__28_, connection_5__8__27_, connection_5__8__26_, 
        connection_5__8__25_, connection_5__8__24_, connection_5__8__23_, 
        connection_5__8__22_, connection_5__8__21_, connection_5__8__20_, 
        connection_5__8__19_, connection_5__8__18_, connection_5__8__17_, 
        connection_5__8__16_, connection_5__8__15_, connection_5__8__14_, 
        connection_5__8__13_, connection_5__8__12_, connection_5__8__11_, 
        connection_5__8__10_, connection_5__8__9_, connection_5__8__8_, 
        connection_5__8__7_, connection_5__8__6_, connection_5__8__5_, 
        connection_5__8__4_, connection_5__8__3_, connection_5__8__2_, 
        connection_5__8__1_, connection_5__8__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[23:22]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_11 second_half_stages_4__group_sec_half_1__switch_sec_half_1__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__13_, 
        connection_valid_4__9_}), .i_data_bus({connection_4__13__31_, 
        connection_4__13__30_, connection_4__13__29_, connection_4__13__28_, 
        connection_4__13__27_, connection_4__13__26_, connection_4__13__25_, 
        connection_4__13__24_, connection_4__13__23_, connection_4__13__22_, 
        connection_4__13__21_, connection_4__13__20_, connection_4__13__19_, 
        connection_4__13__18_, connection_4__13__17_, connection_4__13__16_, 
        connection_4__13__15_, connection_4__13__14_, connection_4__13__13_, 
        connection_4__13__12_, connection_4__13__11_, connection_4__13__10_, 
        connection_4__13__9_, connection_4__13__8_, connection_4__13__7_, 
        connection_4__13__6_, connection_4__13__5_, connection_4__13__4_, 
        connection_4__13__3_, connection_4__13__2_, connection_4__13__1_, 
        connection_4__13__0_, connection_4__9__31_, connection_4__9__30_, 
        connection_4__9__29_, connection_4__9__28_, connection_4__9__27_, 
        connection_4__9__26_, connection_4__9__25_, connection_4__9__24_, 
        connection_4__9__23_, connection_4__9__22_, connection_4__9__21_, 
        connection_4__9__20_, connection_4__9__19_, connection_4__9__18_, 
        connection_4__9__17_, connection_4__9__16_, connection_4__9__15_, 
        connection_4__9__14_, connection_4__9__13_, connection_4__9__12_, 
        connection_4__9__11_, connection_4__9__10_, connection_4__9__9_, 
        connection_4__9__8_, connection_4__9__7_, connection_4__9__6_, 
        connection_4__9__5_, connection_4__9__4_, connection_4__9__3_, 
        connection_4__9__2_, connection_4__9__1_, connection_4__9__0_}), 
        .o_valid({connection_valid_5__11_, connection_valid_5__10_}), 
        .o_data_bus({connection_5__11__31_, connection_5__11__30_, 
        connection_5__11__29_, connection_5__11__28_, connection_5__11__27_, 
        connection_5__11__26_, connection_5__11__25_, connection_5__11__24_, 
        connection_5__11__23_, connection_5__11__22_, connection_5__11__21_, 
        connection_5__11__20_, connection_5__11__19_, connection_5__11__18_, 
        connection_5__11__17_, connection_5__11__16_, connection_5__11__15_, 
        connection_5__11__14_, connection_5__11__13_, connection_5__11__12_, 
        connection_5__11__11_, connection_5__11__10_, connection_5__11__9_, 
        connection_5__11__8_, connection_5__11__7_, connection_5__11__6_, 
        connection_5__11__5_, connection_5__11__4_, connection_5__11__3_, 
        connection_5__11__2_, connection_5__11__1_, connection_5__11__0_, 
        connection_5__10__31_, connection_5__10__30_, connection_5__10__29_, 
        connection_5__10__28_, connection_5__10__27_, connection_5__10__26_, 
        connection_5__10__25_, connection_5__10__24_, connection_5__10__23_, 
        connection_5__10__22_, connection_5__10__21_, connection_5__10__20_, 
        connection_5__10__19_, connection_5__10__18_, connection_5__10__17_, 
        connection_5__10__16_, connection_5__10__15_, connection_5__10__14_, 
        connection_5__10__13_, connection_5__10__12_, connection_5__10__11_, 
        connection_5__10__10_, connection_5__10__9_, connection_5__10__8_, 
        connection_5__10__7_, connection_5__10__6_, connection_5__10__5_, 
        connection_5__10__4_, connection_5__10__3_, connection_5__10__2_, 
        connection_5__10__1_, connection_5__10__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[21:20]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_10 second_half_stages_4__group_sec_half_1__switch_sec_half_2__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__14_, 
        connection_valid_4__10_}), .i_data_bus({connection_4__14__31_, 
        connection_4__14__30_, connection_4__14__29_, connection_4__14__28_, 
        connection_4__14__27_, connection_4__14__26_, connection_4__14__25_, 
        connection_4__14__24_, connection_4__14__23_, connection_4__14__22_, 
        connection_4__14__21_, connection_4__14__20_, connection_4__14__19_, 
        connection_4__14__18_, connection_4__14__17_, connection_4__14__16_, 
        connection_4__14__15_, connection_4__14__14_, connection_4__14__13_, 
        connection_4__14__12_, connection_4__14__11_, connection_4__14__10_, 
        connection_4__14__9_, connection_4__14__8_, connection_4__14__7_, 
        connection_4__14__6_, connection_4__14__5_, connection_4__14__4_, 
        connection_4__14__3_, connection_4__14__2_, connection_4__14__1_, 
        connection_4__14__0_, connection_4__10__31_, connection_4__10__30_, 
        connection_4__10__29_, connection_4__10__28_, connection_4__10__27_, 
        connection_4__10__26_, connection_4__10__25_, connection_4__10__24_, 
        connection_4__10__23_, connection_4__10__22_, connection_4__10__21_, 
        connection_4__10__20_, connection_4__10__19_, connection_4__10__18_, 
        connection_4__10__17_, connection_4__10__16_, connection_4__10__15_, 
        connection_4__10__14_, connection_4__10__13_, connection_4__10__12_, 
        connection_4__10__11_, connection_4__10__10_, connection_4__10__9_, 
        connection_4__10__8_, connection_4__10__7_, connection_4__10__6_, 
        connection_4__10__5_, connection_4__10__4_, connection_4__10__3_, 
        connection_4__10__2_, connection_4__10__1_, connection_4__10__0_}), 
        .o_valid({connection_valid_5__13_, connection_valid_5__12_}), 
        .o_data_bus({connection_5__13__31_, connection_5__13__30_, 
        connection_5__13__29_, connection_5__13__28_, connection_5__13__27_, 
        connection_5__13__26_, connection_5__13__25_, connection_5__13__24_, 
        connection_5__13__23_, connection_5__13__22_, connection_5__13__21_, 
        connection_5__13__20_, connection_5__13__19_, connection_5__13__18_, 
        connection_5__13__17_, connection_5__13__16_, connection_5__13__15_, 
        connection_5__13__14_, connection_5__13__13_, connection_5__13__12_, 
        connection_5__13__11_, connection_5__13__10_, connection_5__13__9_, 
        connection_5__13__8_, connection_5__13__7_, connection_5__13__6_, 
        connection_5__13__5_, connection_5__13__4_, connection_5__13__3_, 
        connection_5__13__2_, connection_5__13__1_, connection_5__13__0_, 
        connection_5__12__31_, connection_5__12__30_, connection_5__12__29_, 
        connection_5__12__28_, connection_5__12__27_, connection_5__12__26_, 
        connection_5__12__25_, connection_5__12__24_, connection_5__12__23_, 
        connection_5__12__22_, connection_5__12__21_, connection_5__12__20_, 
        connection_5__12__19_, connection_5__12__18_, connection_5__12__17_, 
        connection_5__12__16_, connection_5__12__15_, connection_5__12__14_, 
        connection_5__12__13_, connection_5__12__12_, connection_5__12__11_, 
        connection_5__12__10_, connection_5__12__9_, connection_5__12__8_, 
        connection_5__12__7_, connection_5__12__6_, connection_5__12__5_, 
        connection_5__12__4_, connection_5__12__3_, connection_5__12__2_, 
        connection_5__12__1_, connection_5__12__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[19:18]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_9 second_half_stages_4__group_sec_half_1__switch_sec_half_3__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__15_, 
        connection_valid_4__11_}), .i_data_bus({connection_4__15__31_, 
        connection_4__15__30_, connection_4__15__29_, connection_4__15__28_, 
        connection_4__15__27_, connection_4__15__26_, connection_4__15__25_, 
        connection_4__15__24_, connection_4__15__23_, connection_4__15__22_, 
        connection_4__15__21_, connection_4__15__20_, connection_4__15__19_, 
        connection_4__15__18_, connection_4__15__17_, connection_4__15__16_, 
        connection_4__15__15_, connection_4__15__14_, connection_4__15__13_, 
        connection_4__15__12_, connection_4__15__11_, connection_4__15__10_, 
        connection_4__15__9_, connection_4__15__8_, connection_4__15__7_, 
        connection_4__15__6_, connection_4__15__5_, connection_4__15__4_, 
        connection_4__15__3_, connection_4__15__2_, connection_4__15__1_, 
        connection_4__15__0_, connection_4__11__31_, connection_4__11__30_, 
        connection_4__11__29_, connection_4__11__28_, connection_4__11__27_, 
        connection_4__11__26_, connection_4__11__25_, connection_4__11__24_, 
        connection_4__11__23_, connection_4__11__22_, connection_4__11__21_, 
        connection_4__11__20_, connection_4__11__19_, connection_4__11__18_, 
        connection_4__11__17_, connection_4__11__16_, connection_4__11__15_, 
        connection_4__11__14_, connection_4__11__13_, connection_4__11__12_, 
        connection_4__11__11_, connection_4__11__10_, connection_4__11__9_, 
        connection_4__11__8_, connection_4__11__7_, connection_4__11__6_, 
        connection_4__11__5_, connection_4__11__4_, connection_4__11__3_, 
        connection_4__11__2_, connection_4__11__1_, connection_4__11__0_}), 
        .o_valid({connection_valid_5__15_, connection_valid_5__14_}), 
        .o_data_bus({connection_5__15__31_, connection_5__15__30_, 
        connection_5__15__29_, connection_5__15__28_, connection_5__15__27_, 
        connection_5__15__26_, connection_5__15__25_, connection_5__15__24_, 
        connection_5__15__23_, connection_5__15__22_, connection_5__15__21_, 
        connection_5__15__20_, connection_5__15__19_, connection_5__15__18_, 
        connection_5__15__17_, connection_5__15__16_, connection_5__15__15_, 
        connection_5__15__14_, connection_5__15__13_, connection_5__15__12_, 
        connection_5__15__11_, connection_5__15__10_, connection_5__15__9_, 
        connection_5__15__8_, connection_5__15__7_, connection_5__15__6_, 
        connection_5__15__5_, connection_5__15__4_, connection_5__15__3_, 
        connection_5__15__2_, connection_5__15__1_, connection_5__15__0_, 
        connection_5__14__31_, connection_5__14__30_, connection_5__14__29_, 
        connection_5__14__28_, connection_5__14__27_, connection_5__14__26_, 
        connection_5__14__25_, connection_5__14__24_, connection_5__14__23_, 
        connection_5__14__22_, connection_5__14__21_, connection_5__14__20_, 
        connection_5__14__19_, connection_5__14__18_, connection_5__14__17_, 
        connection_5__14__16_, connection_5__14__15_, connection_5__14__14_, 
        connection_5__14__13_, connection_5__14__12_, connection_5__14__11_, 
        connection_5__14__10_, connection_5__14__9_, connection_5__14__8_, 
        connection_5__14__7_, connection_5__14__6_, connection_5__14__5_, 
        connection_5__14__4_, connection_5__14__3_, connection_5__14__2_, 
        connection_5__14__1_, connection_5__14__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[17:16]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_8 second_half_stages_5__group_sec_half_0__switch_sec_half_0__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__8_, 
        connection_valid_5__0_}), .i_data_bus({connection_5__8__31_, 
        connection_5__8__30_, connection_5__8__29_, connection_5__8__28_, 
        connection_5__8__27_, connection_5__8__26_, connection_5__8__25_, 
        connection_5__8__24_, connection_5__8__23_, connection_5__8__22_, 
        connection_5__8__21_, connection_5__8__20_, connection_5__8__19_, 
        connection_5__8__18_, connection_5__8__17_, connection_5__8__16_, 
        connection_5__8__15_, connection_5__8__14_, connection_5__8__13_, 
        connection_5__8__12_, connection_5__8__11_, connection_5__8__10_, 
        connection_5__8__9_, connection_5__8__8_, connection_5__8__7_, 
        connection_5__8__6_, connection_5__8__5_, connection_5__8__4_, 
        connection_5__8__3_, connection_5__8__2_, connection_5__8__1_, 
        connection_5__8__0_, connection_5__0__31_, connection_5__0__30_, 
        connection_5__0__29_, connection_5__0__28_, connection_5__0__27_, 
        connection_5__0__26_, connection_5__0__25_, connection_5__0__24_, 
        connection_5__0__23_, connection_5__0__22_, connection_5__0__21_, 
        connection_5__0__20_, connection_5__0__19_, connection_5__0__18_, 
        connection_5__0__17_, connection_5__0__16_, connection_5__0__15_, 
        connection_5__0__14_, connection_5__0__13_, connection_5__0__12_, 
        connection_5__0__11_, connection_5__0__10_, connection_5__0__9_, 
        connection_5__0__8_, connection_5__0__7_, connection_5__0__6_, 
        connection_5__0__5_, connection_5__0__4_, connection_5__0__3_, 
        connection_5__0__2_, connection_5__0__1_, connection_5__0__0_}), 
        .o_valid({n565, n566}), .o_data_bus({n1015, n1016, n1017, n1018, n1019, 
        n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, 
        n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, 
        n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, 
        n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, 
        n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, 
        n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078}), 
        .i_en(i_en), .i_cmd(cmd_pipeline_stage_5__pipeline_i_cmd_reg[15:14])
         );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_7 second_half_stages_5__group_sec_half_0__switch_sec_half_1__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__9_, 
        connection_valid_5__1_}), .i_data_bus({connection_5__9__31_, 
        connection_5__9__30_, connection_5__9__29_, connection_5__9__28_, 
        connection_5__9__27_, connection_5__9__26_, connection_5__9__25_, 
        connection_5__9__24_, connection_5__9__23_, connection_5__9__22_, 
        connection_5__9__21_, connection_5__9__20_, connection_5__9__19_, 
        connection_5__9__18_, connection_5__9__17_, connection_5__9__16_, 
        connection_5__9__15_, connection_5__9__14_, connection_5__9__13_, 
        connection_5__9__12_, connection_5__9__11_, connection_5__9__10_, 
        connection_5__9__9_, connection_5__9__8_, connection_5__9__7_, 
        connection_5__9__6_, connection_5__9__5_, connection_5__9__4_, 
        connection_5__9__3_, connection_5__9__2_, connection_5__9__1_, 
        connection_5__9__0_, connection_5__1__31_, connection_5__1__30_, 
        connection_5__1__29_, connection_5__1__28_, connection_5__1__27_, 
        connection_5__1__26_, connection_5__1__25_, connection_5__1__24_, 
        connection_5__1__23_, connection_5__1__22_, connection_5__1__21_, 
        connection_5__1__20_, connection_5__1__19_, connection_5__1__18_, 
        connection_5__1__17_, connection_5__1__16_, connection_5__1__15_, 
        connection_5__1__14_, connection_5__1__13_, connection_5__1__12_, 
        connection_5__1__11_, connection_5__1__10_, connection_5__1__9_, 
        connection_5__1__8_, connection_5__1__7_, connection_5__1__6_, 
        connection_5__1__5_, connection_5__1__4_, connection_5__1__3_, 
        connection_5__1__2_, connection_5__1__1_, connection_5__1__0_}), 
        .o_valid({n563, n564}), .o_data_bus({n951, n952, n953, n954, n955, 
        n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, 
        n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, 
        n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, 
        n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, 
        n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
        n1013, n1014}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[13:12]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_6 second_half_stages_5__group_sec_half_0__switch_sec_half_2__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__10_, 
        connection_valid_5__2_}), .i_data_bus({connection_5__10__31_, 
        connection_5__10__30_, connection_5__10__29_, connection_5__10__28_, 
        connection_5__10__27_, connection_5__10__26_, connection_5__10__25_, 
        connection_5__10__24_, connection_5__10__23_, connection_5__10__22_, 
        connection_5__10__21_, connection_5__10__20_, connection_5__10__19_, 
        connection_5__10__18_, connection_5__10__17_, connection_5__10__16_, 
        connection_5__10__15_, connection_5__10__14_, connection_5__10__13_, 
        connection_5__10__12_, connection_5__10__11_, connection_5__10__10_, 
        connection_5__10__9_, connection_5__10__8_, connection_5__10__7_, 
        connection_5__10__6_, connection_5__10__5_, connection_5__10__4_, 
        connection_5__10__3_, connection_5__10__2_, connection_5__10__1_, 
        connection_5__10__0_, connection_5__2__31_, connection_5__2__30_, 
        connection_5__2__29_, connection_5__2__28_, connection_5__2__27_, 
        connection_5__2__26_, connection_5__2__25_, connection_5__2__24_, 
        connection_5__2__23_, connection_5__2__22_, connection_5__2__21_, 
        connection_5__2__20_, connection_5__2__19_, connection_5__2__18_, 
        connection_5__2__17_, connection_5__2__16_, connection_5__2__15_, 
        connection_5__2__14_, connection_5__2__13_, connection_5__2__12_, 
        connection_5__2__11_, connection_5__2__10_, connection_5__2__9_, 
        connection_5__2__8_, connection_5__2__7_, connection_5__2__6_, 
        connection_5__2__5_, connection_5__2__4_, connection_5__2__3_, 
        connection_5__2__2_, connection_5__2__1_, connection_5__2__0_}), 
        .o_valid({n561, n562}), .o_data_bus({n887, n888, n889, n890, n891, 
        n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, 
        n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, 
        n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, 
        n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, 
        n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950}), 
        .i_en(i_en), .i_cmd(cmd_pipeline_stage_5__pipeline_i_cmd_reg[11:10])
         );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_5 second_half_stages_5__group_sec_half_0__switch_sec_half_3__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__11_, 
        connection_valid_5__3_}), .i_data_bus({connection_5__11__31_, 
        connection_5__11__30_, connection_5__11__29_, connection_5__11__28_, 
        connection_5__11__27_, connection_5__11__26_, connection_5__11__25_, 
        connection_5__11__24_, connection_5__11__23_, connection_5__11__22_, 
        connection_5__11__21_, connection_5__11__20_, connection_5__11__19_, 
        connection_5__11__18_, connection_5__11__17_, connection_5__11__16_, 
        connection_5__11__15_, connection_5__11__14_, connection_5__11__13_, 
        connection_5__11__12_, connection_5__11__11_, connection_5__11__10_, 
        connection_5__11__9_, connection_5__11__8_, connection_5__11__7_, 
        connection_5__11__6_, connection_5__11__5_, connection_5__11__4_, 
        connection_5__11__3_, connection_5__11__2_, connection_5__11__1_, 
        connection_5__11__0_, connection_5__3__31_, connection_5__3__30_, 
        connection_5__3__29_, connection_5__3__28_, connection_5__3__27_, 
        connection_5__3__26_, connection_5__3__25_, connection_5__3__24_, 
        connection_5__3__23_, connection_5__3__22_, connection_5__3__21_, 
        connection_5__3__20_, connection_5__3__19_, connection_5__3__18_, 
        connection_5__3__17_, connection_5__3__16_, connection_5__3__15_, 
        connection_5__3__14_, connection_5__3__13_, connection_5__3__12_, 
        connection_5__3__11_, connection_5__3__10_, connection_5__3__9_, 
        connection_5__3__8_, connection_5__3__7_, connection_5__3__6_, 
        connection_5__3__5_, connection_5__3__4_, connection_5__3__3_, 
        connection_5__3__2_, connection_5__3__1_, connection_5__3__0_}), 
        .o_valid({n559, n560}), .o_data_bus({n823, n824, n825, n826, n827, 
        n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, 
        n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, 
        n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, 
        n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, 
        n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886}), 
        .i_en(i_en), .i_cmd(cmd_pipeline_stage_5__pipeline_i_cmd_reg[9:8]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_4 second_half_stages_5__group_sec_half_0__switch_sec_half_4__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__12_, 
        connection_valid_5__4_}), .i_data_bus({connection_5__12__31_, 
        connection_5__12__30_, connection_5__12__29_, connection_5__12__28_, 
        connection_5__12__27_, connection_5__12__26_, connection_5__12__25_, 
        connection_5__12__24_, connection_5__12__23_, connection_5__12__22_, 
        connection_5__12__21_, connection_5__12__20_, connection_5__12__19_, 
        connection_5__12__18_, connection_5__12__17_, connection_5__12__16_, 
        connection_5__12__15_, connection_5__12__14_, connection_5__12__13_, 
        connection_5__12__12_, connection_5__12__11_, connection_5__12__10_, 
        connection_5__12__9_, connection_5__12__8_, connection_5__12__7_, 
        connection_5__12__6_, connection_5__12__5_, connection_5__12__4_, 
        connection_5__12__3_, connection_5__12__2_, connection_5__12__1_, 
        connection_5__12__0_, connection_5__4__31_, connection_5__4__30_, 
        connection_5__4__29_, connection_5__4__28_, connection_5__4__27_, 
        connection_5__4__26_, connection_5__4__25_, connection_5__4__24_, 
        connection_5__4__23_, connection_5__4__22_, connection_5__4__21_, 
        connection_5__4__20_, connection_5__4__19_, connection_5__4__18_, 
        connection_5__4__17_, connection_5__4__16_, connection_5__4__15_, 
        connection_5__4__14_, connection_5__4__13_, connection_5__4__12_, 
        connection_5__4__11_, connection_5__4__10_, connection_5__4__9_, 
        connection_5__4__8_, connection_5__4__7_, connection_5__4__6_, 
        connection_5__4__5_, connection_5__4__4_, connection_5__4__3_, 
        connection_5__4__2_, connection_5__4__1_, connection_5__4__0_}), 
        .o_valid({n557, n558}), .o_data_bus({n759, n760, n761, n762, n763, 
        n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, 
        n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, 
        n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, 
        n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, 
        n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822}), 
        .i_en(i_en), .i_cmd(cmd_pipeline_stage_5__pipeline_i_cmd_reg[7:6]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_3 second_half_stages_5__group_sec_half_0__switch_sec_half_5__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__13_, 
        connection_valid_5__5_}), .i_data_bus({connection_5__13__31_, 
        connection_5__13__30_, connection_5__13__29_, connection_5__13__28_, 
        connection_5__13__27_, connection_5__13__26_, connection_5__13__25_, 
        connection_5__13__24_, connection_5__13__23_, connection_5__13__22_, 
        connection_5__13__21_, connection_5__13__20_, connection_5__13__19_, 
        connection_5__13__18_, connection_5__13__17_, connection_5__13__16_, 
        connection_5__13__15_, connection_5__13__14_, connection_5__13__13_, 
        connection_5__13__12_, connection_5__13__11_, connection_5__13__10_, 
        connection_5__13__9_, connection_5__13__8_, connection_5__13__7_, 
        connection_5__13__6_, connection_5__13__5_, connection_5__13__4_, 
        connection_5__13__3_, connection_5__13__2_, connection_5__13__1_, 
        connection_5__13__0_, connection_5__5__31_, connection_5__5__30_, 
        connection_5__5__29_, connection_5__5__28_, connection_5__5__27_, 
        connection_5__5__26_, connection_5__5__25_, connection_5__5__24_, 
        connection_5__5__23_, connection_5__5__22_, connection_5__5__21_, 
        connection_5__5__20_, connection_5__5__19_, connection_5__5__18_, 
        connection_5__5__17_, connection_5__5__16_, connection_5__5__15_, 
        connection_5__5__14_, connection_5__5__13_, connection_5__5__12_, 
        connection_5__5__11_, connection_5__5__10_, connection_5__5__9_, 
        connection_5__5__8_, connection_5__5__7_, connection_5__5__6_, 
        connection_5__5__5_, connection_5__5__4_, connection_5__5__3_, 
        connection_5__5__2_, connection_5__5__1_, connection_5__5__0_}), 
        .o_valid({n555, n556}), .o_data_bus({n695, n696, n697, n698, n699, 
        n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, 
        n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, 
        n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, 
        n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, 
        n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758}), 
        .i_en(i_en), .i_cmd(cmd_pipeline_stage_5__pipeline_i_cmd_reg[5:4]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_2 second_half_stages_5__group_sec_half_0__switch_sec_half_6__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__14_, 
        connection_valid_5__6_}), .i_data_bus({connection_5__14__31_, 
        connection_5__14__30_, connection_5__14__29_, connection_5__14__28_, 
        connection_5__14__27_, connection_5__14__26_, connection_5__14__25_, 
        connection_5__14__24_, connection_5__14__23_, connection_5__14__22_, 
        connection_5__14__21_, connection_5__14__20_, connection_5__14__19_, 
        connection_5__14__18_, connection_5__14__17_, connection_5__14__16_, 
        connection_5__14__15_, connection_5__14__14_, connection_5__14__13_, 
        connection_5__14__12_, connection_5__14__11_, connection_5__14__10_, 
        connection_5__14__9_, connection_5__14__8_, connection_5__14__7_, 
        connection_5__14__6_, connection_5__14__5_, connection_5__14__4_, 
        connection_5__14__3_, connection_5__14__2_, connection_5__14__1_, 
        connection_5__14__0_, connection_5__6__31_, connection_5__6__30_, 
        connection_5__6__29_, connection_5__6__28_, connection_5__6__27_, 
        connection_5__6__26_, connection_5__6__25_, connection_5__6__24_, 
        connection_5__6__23_, connection_5__6__22_, connection_5__6__21_, 
        connection_5__6__20_, connection_5__6__19_, connection_5__6__18_, 
        connection_5__6__17_, connection_5__6__16_, connection_5__6__15_, 
        connection_5__6__14_, connection_5__6__13_, connection_5__6__12_, 
        connection_5__6__11_, connection_5__6__10_, connection_5__6__9_, 
        connection_5__6__8_, connection_5__6__7_, connection_5__6__6_, 
        connection_5__6__5_, connection_5__6__4_, connection_5__6__3_, 
        connection_5__6__2_, connection_5__6__1_, connection_5__6__0_}), 
        .o_valid({n553, n554}), .o_data_bus({n631, n632, n633, n634, n635, 
        n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, 
        n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, 
        n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, 
        n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, 
        n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694}), 
        .i_en(i_en), .i_cmd(cmd_pipeline_stage_5__pipeline_i_cmd_reg[3:2]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_1 second_half_stages_5__group_sec_half_0__switch_sec_half_7__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__15_, 
        connection_valid_5__7_}), .i_data_bus({connection_5__15__31_, 
        connection_5__15__30_, connection_5__15__29_, connection_5__15__28_, 
        connection_5__15__27_, connection_5__15__26_, connection_5__15__25_, 
        connection_5__15__24_, connection_5__15__23_, connection_5__15__22_, 
        connection_5__15__21_, connection_5__15__20_, connection_5__15__19_, 
        connection_5__15__18_, connection_5__15__17_, connection_5__15__16_, 
        connection_5__15__15_, connection_5__15__14_, connection_5__15__13_, 
        connection_5__15__12_, connection_5__15__11_, connection_5__15__10_, 
        connection_5__15__9_, connection_5__15__8_, connection_5__15__7_, 
        connection_5__15__6_, connection_5__15__5_, connection_5__15__4_, 
        connection_5__15__3_, connection_5__15__2_, connection_5__15__1_, 
        connection_5__15__0_, connection_5__7__31_, connection_5__7__30_, 
        connection_5__7__29_, connection_5__7__28_, connection_5__7__27_, 
        connection_5__7__26_, connection_5__7__25_, connection_5__7__24_, 
        connection_5__7__23_, connection_5__7__22_, connection_5__7__21_, 
        connection_5__7__20_, connection_5__7__19_, connection_5__7__18_, 
        connection_5__7__17_, connection_5__7__16_, connection_5__7__15_, 
        connection_5__7__14_, connection_5__7__13_, connection_5__7__12_, 
        connection_5__7__11_, connection_5__7__10_, connection_5__7__9_, 
        connection_5__7__8_, connection_5__7__7_, connection_5__7__6_, 
        connection_5__7__5_, connection_5__7__4_, connection_5__7__3_, 
        connection_5__7__2_, connection_5__7__1_, connection_5__7__0_}), 
        .o_valid({n551, n552}), .o_data_bus({n567, n568, n569, n570, n571, 
        n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, 
        n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, 
        n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, 
        n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, 
        n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630}), 
        .i_en(i_en), .i_cmd(cmd_pipeline_stage_5__pipeline_i_cmd_reg[1:0]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__0__1_ ( .D(
        i_cmd[33]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[79])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__0__0_ ( .D(
        i_cmd[32]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[78])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__1__1_ ( .D(
        i_cmd[35]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[77])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__1__0_ ( .D(
        i_cmd[34]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[76])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__2__1_ ( .D(
        i_cmd[37]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[75])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__2__0_ ( .D(
        i_cmd[36]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[74])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__3__1_ ( .D(
        i_cmd[39]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[73])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__3__0_ ( .D(
        i_cmd[38]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[72])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__4__1_ ( .D(
        i_cmd[41]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[71])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__4__0_ ( .D(
        i_cmd[40]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[70])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__5__1_ ( .D(
        i_cmd[43]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[69])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__5__0_ ( .D(
        i_cmd[42]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[68])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__6__1_ ( .D(
        i_cmd[45]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[67])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__6__0_ ( .D(
        i_cmd[44]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[66])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__7__1_ ( .D(
        i_cmd[47]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[65])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__7__0_ ( .D(
        i_cmd[46]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[64])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__0__1_ ( .D(
        i_cmd[49]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[63])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__0__0_ ( .D(
        i_cmd[48]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[62])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__1__1_ ( .D(
        i_cmd[51]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[61])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__1__0_ ( .D(
        i_cmd[50]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[60])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__2__1_ ( .D(
        i_cmd[53]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[59])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__2__0_ ( .D(
        i_cmd[52]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[58])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__3__1_ ( .D(
        i_cmd[55]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[57])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__3__0_ ( .D(
        i_cmd[54]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[56])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__4__1_ ( .D(
        i_cmd[57]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[55])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__4__0_ ( .D(
        i_cmd[56]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[54])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__5__1_ ( .D(
        i_cmd[59]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[53])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__5__0_ ( .D(
        i_cmd[58]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[52])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__6__1_ ( .D(
        i_cmd[61]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[51])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__6__0_ ( .D(
        i_cmd[60]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[50])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__7__1_ ( .D(
        i_cmd[63]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[49])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__7__0_ ( .D(
        i_cmd[62]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[48])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__0__1_ ( .D(
        i_cmd[65]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[47])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__0__0_ ( .D(
        i_cmd[64]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[46])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__1__1_ ( .D(
        i_cmd[67]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[45])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__1__0_ ( .D(
        i_cmd[66]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[44])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__2__1_ ( .D(
        i_cmd[69]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[43])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__2__0_ ( .D(
        i_cmd[68]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[42])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__3__1_ ( .D(
        i_cmd[71]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[41])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__3__0_ ( .D(
        i_cmd[70]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[40])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__4__1_ ( .D(
        i_cmd[73]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[39])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__4__0_ ( .D(
        i_cmd[72]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[38])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__5__1_ ( .D(
        i_cmd[75]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[37])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__5__0_ ( .D(
        i_cmd[74]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[36])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__6__1_ ( .D(
        i_cmd[77]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[35])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__6__0_ ( .D(
        i_cmd[76]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[34])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__7__1_ ( .D(
        i_cmd[79]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[33])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__7__0_ ( .D(
        i_cmd[78]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[32])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__0__1_ ( .D(
        i_cmd[81]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[31])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__0__0_ ( .D(
        i_cmd[80]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[30])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__1__1_ ( .D(
        i_cmd[83]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[29])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__1__0_ ( .D(
        i_cmd[82]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[28])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__2__1_ ( .D(
        i_cmd[85]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[27])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__2__0_ ( .D(
        i_cmd[84]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[26])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__3__1_ ( .D(
        i_cmd[87]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[25])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__3__0_ ( .D(
        i_cmd[86]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[24])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__4__1_ ( .D(
        i_cmd[89]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[23])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__4__0_ ( .D(
        i_cmd[88]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[22])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__5__1_ ( .D(
        i_cmd[91]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[21])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__5__0_ ( .D(
        i_cmd[90]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[20])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__6__1_ ( .D(
        i_cmd[93]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[19])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__6__0_ ( .D(
        i_cmd[92]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[18])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__7__1_ ( .D(
        i_cmd[95]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[17])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__7__0_ ( .D(
        i_cmd[94]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[16])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__0__1_ ( .D(
        i_cmd[97]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[15])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__0__0_ ( .D(
        i_cmd[96]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[14])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__1__1_ ( .D(
        i_cmd[99]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[13])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__1__0_ ( .D(
        i_cmd[98]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[12])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__2__1_ ( .D(
        i_cmd[101]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[11]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__2__0_ ( .D(
        i_cmd[100]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[10]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__3__1_ ( .D(
        i_cmd[103]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[9])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__3__0_ ( .D(
        i_cmd[102]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[8])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__4__1_ ( .D(
        i_cmd[105]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[7])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__4__0_ ( .D(
        i_cmd[104]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[6])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__5__1_ ( .D(
        i_cmd[107]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[5])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__5__0_ ( .D(
        i_cmd[106]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[4])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__6__1_ ( .D(
        i_cmd[109]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[3])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__6__0_ ( .D(
        i_cmd[108]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[2])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__7__1_ ( .D(
        i_cmd[111]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[1])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__7__0_ ( .D(
        i_cmd[110]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[0])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__0__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[63]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[63]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__0__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[62]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[62]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__1__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[61]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[61]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__1__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[60]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[60]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__2__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[59]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[59]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__2__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[58]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[58]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__3__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[57]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[57]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__3__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[56]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[56]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__4__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[55]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[55]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__4__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[54]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[54]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__5__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[53]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[53]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__5__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[52]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[52]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__6__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[51]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[51]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__6__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[50]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[50]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__7__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[49]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[49]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__7__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[48]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[48]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__0__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[47]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[47]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__0__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[46]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[46]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__1__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[45]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[45]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__1__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[44]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[44]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__2__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[43]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[43]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__2__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[42]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[42]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__3__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[41]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[41]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__3__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[40]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[40]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__4__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[39]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[39]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__4__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[38]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[38]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__5__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[37]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[37]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__5__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[36]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[36]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__6__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[35]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[35]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__6__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[34]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[34]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__7__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[33]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[33]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__7__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[32]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[32]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__0__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[31]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[31]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__0__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[30]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[30]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__1__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[29]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[29]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__1__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[28]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[28]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__2__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[27]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[27]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__2__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[26]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[26]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__3__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[25]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[25]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__3__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[24]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[24]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__4__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[23]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[23]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__4__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[22]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[22]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__5__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[21]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[21]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__5__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[20]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[20]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__6__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[19]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[19]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__6__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[18]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[18]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__7__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[17]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[17]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__7__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[16]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[16]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__0__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[15]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[15]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__0__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[14]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[14]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__1__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[13]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[13]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__1__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[12]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[12]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__2__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[11]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[11]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__2__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[10]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[10]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__3__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[9]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[9]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__3__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[8]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[8]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__4__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[7]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[7]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__4__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[6]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[6]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__5__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[5]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[5]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__5__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[4]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[4]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__6__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[3]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[3]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__6__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[2]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[2]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__7__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[1]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[1]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__7__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[0]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[0]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__0__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[47]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[47]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__0__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[46]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[46]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__1__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[45]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[45]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__1__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[44]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[44]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__2__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[43]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[43]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__2__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[42]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[42]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__3__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[41]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[41]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__3__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[40]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[40]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__4__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[39]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[39]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__4__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[38]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[38]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__5__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[37]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[37]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__5__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[36]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[36]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__6__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[35]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[35]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__6__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[34]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[34]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__7__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[33]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[33]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__7__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[32]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[32]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__0__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[31]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[31]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__0__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[30]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[30]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__1__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[29]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[29]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__1__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[28]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[28]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__2__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[27]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[27]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__2__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[26]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[26]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__3__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[25]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[25]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__3__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[24]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[24]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__4__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[23]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[23]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__4__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[22]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[22]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__5__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[21]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[21]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__5__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[20]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[20]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__6__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[19]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[19]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__6__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[18]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[18]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__7__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[17]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[17]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__7__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[16]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[16]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__0__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[15]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[15]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__0__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[14]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[14]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__1__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[13]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[13]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__1__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[12]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[12]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__2__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[11]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[11]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__2__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[10]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[10]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__3__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[9]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[9]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__3__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[8]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[8]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__4__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[7]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[7]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__4__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[6]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[6]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__5__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[5]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[5]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__5__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[4]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[4]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__6__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[3]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[3]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__6__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[2]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[2]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__7__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[1]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[1]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__7__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[0]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[0]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__0__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[31]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[31]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__0__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[30]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[30]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__1__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[29]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[29]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__1__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[28]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[28]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__2__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[27]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[27]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__2__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[26]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[26]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__3__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[25]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[25]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__3__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[24]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[24]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__4__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[23]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[23]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__4__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[22]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[22]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__5__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[21]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[21]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__5__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[20]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[20]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__6__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[19]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[19]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__6__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[18]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[18]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__7__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[17]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[17]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__7__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[16]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[16]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__0__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[15]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[15]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__0__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[14]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[14]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__1__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[13]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[13]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__1__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[12]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[12]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__2__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[11]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[11]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__2__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[10]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[10]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__3__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[9]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[9]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__3__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[8]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[8]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__4__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[7]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[7]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__4__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[6]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[6]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__5__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[5]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[5]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__5__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[4]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[4]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__6__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[3]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[3]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__6__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[2]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[2]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__7__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[1]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[1]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__7__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[0]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[0]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__0__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[15]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[15]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__0__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[14]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[14]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__1__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[13]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[13]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__1__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[12]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[12]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__2__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[11]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[11]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__2__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[10]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[10]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__3__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[9]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[9]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__3__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[8]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[8]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__4__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[7]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[7]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__4__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[6]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[6]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__5__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[5]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[5]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__5__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[4]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[4]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__6__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[3]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[3]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__6__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[2]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[2]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__7__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[1]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[1]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__7__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[0]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[0]) );
  DFQD4BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__4__1_ ( .D(
        i_cmd[25]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[87])
         );
  DFQD4BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__5__1_ ( .D(
        i_cmd[27]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[85])
         );
  DFQD4BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__6__1_ ( .D(
        i_cmd[29]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[83])
         );
  DFQD4BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__7__1_ ( .D(
        i_cmd[31]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[81])
         );
  DFQD4BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__0__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[14]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[14]) );
  DFQD4BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__0__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[15]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[15]) );
  DFQD4BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__7__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[1]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[1]) );
  DFQD2BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__6__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[34]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[34]) );
  DFQD2BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__7__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[32]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[32]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__0__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[30]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[30]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__1__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[28]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[28]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__2__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[26]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[26]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__3__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[24]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[24]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__4__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[22]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[22]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__5__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[20]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[20]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__6__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[18]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[18]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__7__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[16]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[16]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__6__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[2]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[2]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__5__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[4]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[4]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__4__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[6]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[6]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__3__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[8]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[8]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__2__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[10]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[10]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__1__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[12]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[12]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__5__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[36]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[36]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__4__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[38]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[38]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__3__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[40]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[40]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__2__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[42]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[42]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__1__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[44]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[44]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__0__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[46]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[46]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__7__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[48]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[48]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__6__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[50]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[50]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__5__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[52]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[52]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__4__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[54]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[54]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__3__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[56]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[56]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__2__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[58]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[58]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__1__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[60]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[60]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__0__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[62]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[62]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__7__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[64]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[64]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__6__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[66]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[66]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__5__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[68]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[68]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__4__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[70]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[70]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__3__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[72]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[72]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__2__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[74]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[74]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__1__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[76]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[76]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__0__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[78]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[78]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__7__0_ ( .D(
        i_cmd[30]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[80])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__6__0_ ( .D(
        i_cmd[28]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[82])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__5__0_ ( .D(
        i_cmd[26]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[84])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__4__0_ ( .D(
        i_cmd[24]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[86])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__3__0_ ( .D(
        i_cmd[22]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[88])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__2__0_ ( .D(
        i_cmd[20]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[90])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__1__0_ ( .D(
        i_cmd[18]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[92])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__0__0_ ( .D(
        i_cmd[16]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[94])
         );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__7__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[0]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[0]) );
  DFQD2BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__1__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[77]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[77]) );
  DFQD2BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__1__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[61]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[61]) );
  DFQD2BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__2__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[59]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[59]) );
  DFQD2BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__3__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[57]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[57]) );
  DFQD2BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__5__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[53]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[53]) );
  DFQD2BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__0__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[47]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[47]) );
  DFQD2BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__1__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[45]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[45]) );
  DFQD2BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__2__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[43]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[43]) );
  DFQD2BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__3__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[41]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[41]) );
  DFQD2BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__4__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[39]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[39]) );
  DFQD2BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__5__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[37]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[37]) );
  DFQD2BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__0__1_ ( .D(
        i_cmd[17]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[95])
         );
  DFQD2BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__1__1_ ( .D(
        i_cmd[19]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[93])
         );
  DFQD2BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__2__1_ ( .D(
        i_cmd[21]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[91])
         );
  DFQD2BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__3__1_ ( .D(
        i_cmd[23]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[89])
         );
  DFQD2BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__0__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[79]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[79]) );
  DFQD2BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__2__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[75]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[75]) );
  DFQD2BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__3__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[73]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[73]) );
  DFQD2BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__4__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[71]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[71]) );
  DFQD2BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__5__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[69]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[69]) );
  DFQD2BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__6__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[67]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[67]) );
  DFQD2BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__7__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[65]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[65]) );
  DFQD2BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__0__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[63]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[63]) );
  DFQD2BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__4__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[55]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[55]) );
  DFQD2BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__6__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[51]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[51]) );
  DFQD2BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__7__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[49]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[49]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__6__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[3]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[3]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__5__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[5]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[5]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__4__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[7]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[7]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__3__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[9]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[9]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__2__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[11]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[11]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__1__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[13]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[13]) );
  DFQD2BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__7__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[33]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[33]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__4__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[23]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[23]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__6__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[19]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[19]) );
  DFQD2BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__6__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[35]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[35]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__0__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[31]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[31]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__1__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[29]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[29]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__2__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[27]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[27]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__3__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[25]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[25]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__5__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[21]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[21]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__7__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[17]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[17]) );
  INVD12BWP30P140 U5 ( .I(n11), .ZN(o_data_bus[19]) );
  INVD3BWP30P140 U6 ( .I(n1059), .ZN(n11) );
  INVD12BWP30P140 U7 ( .I(n12), .ZN(o_data_bus[20]) );
  INVD3BWP30P140 U8 ( .I(n1058), .ZN(n12) );
  INVD12BWP30P140 U9 ( .I(n13), .ZN(o_data_bus[21]) );
  INVD3BWP30P140 U10 ( .I(n1057), .ZN(n13) );
  INVD12BWP30P140 U11 ( .I(n14), .ZN(o_data_bus[22]) );
  INVD3BWP30P140 U12 ( .I(n1056), .ZN(n14) );
  INVD12BWP30P140 U13 ( .I(n15), .ZN(o_data_bus[23]) );
  INVD3BWP30P140 U14 ( .I(n1055), .ZN(n15) );
  INVD12BWP30P140 U15 ( .I(n16), .ZN(o_data_bus[24]) );
  INVD3BWP30P140 U16 ( .I(n1054), .ZN(n16) );
  INVD12BWP30P140 U17 ( .I(n17), .ZN(o_data_bus[25]) );
  INVD3BWP30P140 U18 ( .I(n1053), .ZN(n17) );
  INVD12BWP30P140 U19 ( .I(n18), .ZN(o_data_bus[26]) );
  INVD3BWP30P140 U20 ( .I(n1052), .ZN(n18) );
  INVD12BWP30P140 U21 ( .I(n19), .ZN(o_data_bus[27]) );
  INVD3BWP30P140 U22 ( .I(n1051), .ZN(n19) );
  INVD12BWP30P140 U23 ( .I(n20), .ZN(o_data_bus[28]) );
  INVD3BWP30P140 U24 ( .I(n1050), .ZN(n20) );
  INVD12BWP30P140 U25 ( .I(n21), .ZN(o_data_bus[29]) );
  INVD3BWP30P140 U26 ( .I(n1049), .ZN(n21) );
  INVD12BWP30P140 U27 ( .I(n22), .ZN(o_data_bus[30]) );
  INVD3BWP30P140 U28 ( .I(n1048), .ZN(n22) );
  INVD12BWP30P140 U29 ( .I(n23), .ZN(o_data_bus[31]) );
  INVD3BWP30P140 U30 ( .I(n1047), .ZN(n23) );
  INVD12BWP30P140 U31 ( .I(n24), .ZN(o_data_bus[453]) );
  INVD3BWP30P140 U32 ( .I(n625), .ZN(n24) );
  INVD12BWP30P140 U33 ( .I(n25), .ZN(o_data_bus[455]) );
  INVD3BWP30P140 U34 ( .I(n623), .ZN(n25) );
  INVD12BWP30P140 U35 ( .I(n26), .ZN(o_data_bus[470]) );
  INVD3BWP30P140 U36 ( .I(n608), .ZN(n26) );
  INVD12BWP30P140 U37 ( .I(n27), .ZN(o_data_bus[472]) );
  INVD3BWP30P140 U38 ( .I(n606), .ZN(n27) );
  INVD12BWP30P140 U39 ( .I(n28), .ZN(o_data_bus[474]) );
  INVD3BWP30P140 U40 ( .I(n604), .ZN(n28) );
  INVD12BWP30P140 U41 ( .I(n29), .ZN(o_data_bus[476]) );
  INVD3BWP30P140 U42 ( .I(n602), .ZN(n29) );
  INVD12BWP30P140 U43 ( .I(n30), .ZN(o_data_bus[478]) );
  INVD3BWP30P140 U44 ( .I(n600), .ZN(n30) );
  BUFFD12BWP30P140 U45 ( .I(n565), .Z(o_valid[1]) );
  BUFFD12BWP30P140 U46 ( .I(n563), .Z(o_valid[3]) );
  BUFFD12BWP30P140 U47 ( .I(n561), .Z(o_valid[5]) );
  BUFFD12BWP30P140 U48 ( .I(n559), .Z(o_valid[7]) );
  BUFFD12BWP30P140 U49 ( .I(n557), .Z(o_valid[9]) );
  BUFFD12BWP30P140 U50 ( .I(n555), .Z(o_valid[11]) );
  BUFFD12BWP30P140 U51 ( .I(n553), .Z(o_valid[13]) );
  BUFFD12BWP30P140 U52 ( .I(n551), .Z(o_valid[15]) );
  BUFFD12BWP30P140 U53 ( .I(n1074), .Z(o_data_bus[4]) );
  BUFFD12BWP30P140 U54 ( .I(n1075), .Z(o_data_bus[3]) );
  BUFFD12BWP30P140 U55 ( .I(n1076), .Z(o_data_bus[2]) );
  BUFFD12BWP30P140 U56 ( .I(n1077), .Z(o_data_bus[1]) );
  BUFFD12BWP30P140 U57 ( .I(n1078), .Z(o_data_bus[0]) );
  BUFFD12BWP30P140 U58 ( .I(n1071), .Z(o_data_bus[7]) );
  BUFFD12BWP30P140 U59 ( .I(n1072), .Z(o_data_bus[6]) );
  BUFFD12BWP30P140 U60 ( .I(n1073), .Z(o_data_bus[5]) );
  BUFFD12BWP30P140 U61 ( .I(n1060), .Z(o_data_bus[18]) );
  BUFFD12BWP30P140 U62 ( .I(n1061), .Z(o_data_bus[17]) );
  BUFFD12BWP30P140 U63 ( .I(n1062), .Z(o_data_bus[16]) );
  BUFFD12BWP30P140 U64 ( .I(n1063), .Z(o_data_bus[15]) );
  BUFFD12BWP30P140 U65 ( .I(n1064), .Z(o_data_bus[14]) );
  BUFFD12BWP30P140 U66 ( .I(n1065), .Z(o_data_bus[13]) );
  BUFFD12BWP30P140 U67 ( .I(n1066), .Z(o_data_bus[12]) );
  BUFFD12BWP30P140 U68 ( .I(n1067), .Z(o_data_bus[11]) );
  BUFFD12BWP30P140 U69 ( .I(n1068), .Z(o_data_bus[10]) );
  BUFFD12BWP30P140 U70 ( .I(n1069), .Z(o_data_bus[9]) );
  BUFFD12BWP30P140 U71 ( .I(n1070), .Z(o_data_bus[8]) );
  BUFFD12BWP30P140 U72 ( .I(n1046), .Z(o_data_bus[32]) );
  BUFFD12BWP30P140 U73 ( .I(n1045), .Z(o_data_bus[33]) );
  BUFFD12BWP30P140 U74 ( .I(n1044), .Z(o_data_bus[34]) );
  BUFFD12BWP30P140 U75 ( .I(n1043), .Z(o_data_bus[35]) );
  BUFFD12BWP30P140 U76 ( .I(n1042), .Z(o_data_bus[36]) );
  BUFFD12BWP30P140 U77 ( .I(n1041), .Z(o_data_bus[37]) );
  BUFFD12BWP30P140 U78 ( .I(n1040), .Z(o_data_bus[38]) );
  BUFFD12BWP30P140 U79 ( .I(n1039), .Z(o_data_bus[39]) );
  BUFFD12BWP30P140 U80 ( .I(n1038), .Z(o_data_bus[40]) );
  BUFFD12BWP30P140 U81 ( .I(n1037), .Z(o_data_bus[41]) );
  BUFFD12BWP30P140 U82 ( .I(n1036), .Z(o_data_bus[42]) );
  BUFFD12BWP30P140 U83 ( .I(n1035), .Z(o_data_bus[43]) );
  BUFFD12BWP30P140 U84 ( .I(n1034), .Z(o_data_bus[44]) );
  BUFFD12BWP30P140 U85 ( .I(n1033), .Z(o_data_bus[45]) );
  BUFFD12BWP30P140 U86 ( .I(n1032), .Z(o_data_bus[46]) );
  BUFFD12BWP30P140 U87 ( .I(n1031), .Z(o_data_bus[47]) );
  BUFFD12BWP30P140 U88 ( .I(n1030), .Z(o_data_bus[48]) );
  BUFFD12BWP30P140 U89 ( .I(n1029), .Z(o_data_bus[49]) );
  BUFFD12BWP30P140 U90 ( .I(n1028), .Z(o_data_bus[50]) );
  BUFFD12BWP30P140 U91 ( .I(n1027), .Z(o_data_bus[51]) );
  BUFFD12BWP30P140 U92 ( .I(n1026), .Z(o_data_bus[52]) );
  BUFFD12BWP30P140 U93 ( .I(n1025), .Z(o_data_bus[53]) );
  BUFFD12BWP30P140 U94 ( .I(n1024), .Z(o_data_bus[54]) );
  BUFFD12BWP30P140 U95 ( .I(n1023), .Z(o_data_bus[55]) );
  BUFFD12BWP30P140 U96 ( .I(n1022), .Z(o_data_bus[56]) );
  BUFFD12BWP30P140 U97 ( .I(n1021), .Z(o_data_bus[57]) );
  BUFFD12BWP30P140 U98 ( .I(n1020), .Z(o_data_bus[58]) );
  BUFFD12BWP30P140 U99 ( .I(n1019), .Z(o_data_bus[59]) );
  BUFFD12BWP30P140 U100 ( .I(n1018), .Z(o_data_bus[60]) );
  BUFFD12BWP30P140 U101 ( .I(n1017), .Z(o_data_bus[61]) );
  BUFFD12BWP30P140 U102 ( .I(n1016), .Z(o_data_bus[62]) );
  BUFFD12BWP30P140 U103 ( .I(n1015), .Z(o_data_bus[63]) );
  BUFFD12BWP30P140 U104 ( .I(n1014), .Z(o_data_bus[64]) );
  BUFFD12BWP30P140 U105 ( .I(n1013), .Z(o_data_bus[65]) );
  BUFFD12BWP30P140 U106 ( .I(n1012), .Z(o_data_bus[66]) );
  BUFFD12BWP30P140 U107 ( .I(n1011), .Z(o_data_bus[67]) );
  BUFFD12BWP30P140 U108 ( .I(n1010), .Z(o_data_bus[68]) );
  BUFFD12BWP30P140 U109 ( .I(n1009), .Z(o_data_bus[69]) );
  BUFFD12BWP30P140 U110 ( .I(n1008), .Z(o_data_bus[70]) );
  BUFFD12BWP30P140 U111 ( .I(n1007), .Z(o_data_bus[71]) );
  BUFFD12BWP30P140 U112 ( .I(n1006), .Z(o_data_bus[72]) );
  BUFFD12BWP30P140 U113 ( .I(n1005), .Z(o_data_bus[73]) );
  BUFFD12BWP30P140 U114 ( .I(n1004), .Z(o_data_bus[74]) );
  BUFFD12BWP30P140 U115 ( .I(n1003), .Z(o_data_bus[75]) );
  BUFFD12BWP30P140 U116 ( .I(n1002), .Z(o_data_bus[76]) );
  BUFFD12BWP30P140 U117 ( .I(n1001), .Z(o_data_bus[77]) );
  BUFFD12BWP30P140 U118 ( .I(n1000), .Z(o_data_bus[78]) );
  BUFFD12BWP30P140 U119 ( .I(n999), .Z(o_data_bus[79]) );
  BUFFD12BWP30P140 U120 ( .I(n998), .Z(o_data_bus[80]) );
  BUFFD12BWP30P140 U121 ( .I(n997), .Z(o_data_bus[81]) );
  BUFFD12BWP30P140 U122 ( .I(n996), .Z(o_data_bus[82]) );
  BUFFD12BWP30P140 U123 ( .I(n995), .Z(o_data_bus[83]) );
  BUFFD12BWP30P140 U124 ( .I(n994), .Z(o_data_bus[84]) );
  BUFFD12BWP30P140 U125 ( .I(n993), .Z(o_data_bus[85]) );
  BUFFD12BWP30P140 U126 ( .I(n992), .Z(o_data_bus[86]) );
  BUFFD12BWP30P140 U127 ( .I(n991), .Z(o_data_bus[87]) );
  BUFFD12BWP30P140 U128 ( .I(n990), .Z(o_data_bus[88]) );
  BUFFD12BWP30P140 U129 ( .I(n989), .Z(o_data_bus[89]) );
  BUFFD12BWP30P140 U130 ( .I(n988), .Z(o_data_bus[90]) );
  BUFFD12BWP30P140 U131 ( .I(n987), .Z(o_data_bus[91]) );
  BUFFD12BWP30P140 U132 ( .I(n986), .Z(o_data_bus[92]) );
  BUFFD12BWP30P140 U133 ( .I(n985), .Z(o_data_bus[93]) );
  BUFFD12BWP30P140 U134 ( .I(n984), .Z(o_data_bus[94]) );
  BUFFD12BWP30P140 U135 ( .I(n983), .Z(o_data_bus[95]) );
  BUFFD12BWP30P140 U136 ( .I(n982), .Z(o_data_bus[96]) );
  BUFFD12BWP30P140 U137 ( .I(n981), .Z(o_data_bus[97]) );
  BUFFD12BWP30P140 U138 ( .I(n980), .Z(o_data_bus[98]) );
  BUFFD12BWP30P140 U139 ( .I(n979), .Z(o_data_bus[99]) );
  BUFFD12BWP30P140 U140 ( .I(n978), .Z(o_data_bus[100]) );
  BUFFD12BWP30P140 U141 ( .I(n977), .Z(o_data_bus[101]) );
  BUFFD12BWP30P140 U142 ( .I(n976), .Z(o_data_bus[102]) );
  BUFFD12BWP30P140 U143 ( .I(n975), .Z(o_data_bus[103]) );
  BUFFD12BWP30P140 U144 ( .I(n974), .Z(o_data_bus[104]) );
  BUFFD12BWP30P140 U145 ( .I(n973), .Z(o_data_bus[105]) );
  BUFFD12BWP30P140 U146 ( .I(n972), .Z(o_data_bus[106]) );
  BUFFD12BWP30P140 U147 ( .I(n971), .Z(o_data_bus[107]) );
  BUFFD12BWP30P140 U148 ( .I(n970), .Z(o_data_bus[108]) );
  BUFFD12BWP30P140 U149 ( .I(n969), .Z(o_data_bus[109]) );
  BUFFD12BWP30P140 U150 ( .I(n968), .Z(o_data_bus[110]) );
  BUFFD12BWP30P140 U151 ( .I(n967), .Z(o_data_bus[111]) );
  BUFFD12BWP30P140 U152 ( .I(n966), .Z(o_data_bus[112]) );
  BUFFD12BWP30P140 U153 ( .I(n965), .Z(o_data_bus[113]) );
  BUFFD12BWP30P140 U154 ( .I(n964), .Z(o_data_bus[114]) );
  BUFFD12BWP30P140 U155 ( .I(n963), .Z(o_data_bus[115]) );
  BUFFD12BWP30P140 U156 ( .I(n962), .Z(o_data_bus[116]) );
  BUFFD12BWP30P140 U157 ( .I(n961), .Z(o_data_bus[117]) );
  BUFFD12BWP30P140 U158 ( .I(n960), .Z(o_data_bus[118]) );
  BUFFD12BWP30P140 U159 ( .I(n959), .Z(o_data_bus[119]) );
  BUFFD12BWP30P140 U160 ( .I(n958), .Z(o_data_bus[120]) );
  BUFFD12BWP30P140 U161 ( .I(n957), .Z(o_data_bus[121]) );
  BUFFD12BWP30P140 U162 ( .I(n956), .Z(o_data_bus[122]) );
  BUFFD12BWP30P140 U163 ( .I(n955), .Z(o_data_bus[123]) );
  BUFFD12BWP30P140 U164 ( .I(n954), .Z(o_data_bus[124]) );
  BUFFD12BWP30P140 U165 ( .I(n953), .Z(o_data_bus[125]) );
  BUFFD12BWP30P140 U166 ( .I(n952), .Z(o_data_bus[126]) );
  BUFFD12BWP30P140 U167 ( .I(n951), .Z(o_data_bus[127]) );
  BUFFD12BWP30P140 U168 ( .I(n950), .Z(o_data_bus[128]) );
  BUFFD12BWP30P140 U169 ( .I(n949), .Z(o_data_bus[129]) );
  BUFFD12BWP30P140 U170 ( .I(n948), .Z(o_data_bus[130]) );
  BUFFD12BWP30P140 U171 ( .I(n947), .Z(o_data_bus[131]) );
  BUFFD12BWP30P140 U172 ( .I(n946), .Z(o_data_bus[132]) );
  BUFFD12BWP30P140 U173 ( .I(n945), .Z(o_data_bus[133]) );
  BUFFD12BWP30P140 U174 ( .I(n944), .Z(o_data_bus[134]) );
  BUFFD12BWP30P140 U175 ( .I(n943), .Z(o_data_bus[135]) );
  BUFFD12BWP30P140 U176 ( .I(n942), .Z(o_data_bus[136]) );
  BUFFD12BWP30P140 U177 ( .I(n941), .Z(o_data_bus[137]) );
  BUFFD12BWP30P140 U178 ( .I(n940), .Z(o_data_bus[138]) );
  BUFFD12BWP30P140 U179 ( .I(n939), .Z(o_data_bus[139]) );
  BUFFD12BWP30P140 U180 ( .I(n938), .Z(o_data_bus[140]) );
  BUFFD12BWP30P140 U181 ( .I(n937), .Z(o_data_bus[141]) );
  BUFFD12BWP30P140 U182 ( .I(n936), .Z(o_data_bus[142]) );
  BUFFD12BWP30P140 U183 ( .I(n935), .Z(o_data_bus[143]) );
  BUFFD12BWP30P140 U184 ( .I(n934), .Z(o_data_bus[144]) );
  BUFFD12BWP30P140 U185 ( .I(n933), .Z(o_data_bus[145]) );
  BUFFD12BWP30P140 U186 ( .I(n932), .Z(o_data_bus[146]) );
  BUFFD12BWP30P140 U187 ( .I(n931), .Z(o_data_bus[147]) );
  BUFFD12BWP30P140 U188 ( .I(n930), .Z(o_data_bus[148]) );
  BUFFD12BWP30P140 U189 ( .I(n929), .Z(o_data_bus[149]) );
  BUFFD12BWP30P140 U190 ( .I(n928), .Z(o_data_bus[150]) );
  BUFFD12BWP30P140 U191 ( .I(n927), .Z(o_data_bus[151]) );
  BUFFD12BWP30P140 U192 ( .I(n926), .Z(o_data_bus[152]) );
  BUFFD12BWP30P140 U193 ( .I(n925), .Z(o_data_bus[153]) );
  BUFFD12BWP30P140 U194 ( .I(n924), .Z(o_data_bus[154]) );
  BUFFD12BWP30P140 U195 ( .I(n923), .Z(o_data_bus[155]) );
  BUFFD12BWP30P140 U196 ( .I(n922), .Z(o_data_bus[156]) );
  BUFFD12BWP30P140 U197 ( .I(n921), .Z(o_data_bus[157]) );
  BUFFD12BWP30P140 U198 ( .I(n920), .Z(o_data_bus[158]) );
  BUFFD12BWP30P140 U199 ( .I(n919), .Z(o_data_bus[159]) );
  BUFFD12BWP30P140 U200 ( .I(n918), .Z(o_data_bus[160]) );
  BUFFD12BWP30P140 U201 ( .I(n917), .Z(o_data_bus[161]) );
  BUFFD12BWP30P140 U202 ( .I(n916), .Z(o_data_bus[162]) );
  BUFFD12BWP30P140 U203 ( .I(n915), .Z(o_data_bus[163]) );
  BUFFD12BWP30P140 U204 ( .I(n914), .Z(o_data_bus[164]) );
  BUFFD12BWP30P140 U205 ( .I(n913), .Z(o_data_bus[165]) );
  BUFFD12BWP30P140 U206 ( .I(n912), .Z(o_data_bus[166]) );
  BUFFD12BWP30P140 U207 ( .I(n911), .Z(o_data_bus[167]) );
  BUFFD12BWP30P140 U208 ( .I(n910), .Z(o_data_bus[168]) );
  BUFFD12BWP30P140 U209 ( .I(n909), .Z(o_data_bus[169]) );
  BUFFD12BWP30P140 U210 ( .I(n908), .Z(o_data_bus[170]) );
  BUFFD12BWP30P140 U211 ( .I(n907), .Z(o_data_bus[171]) );
  BUFFD12BWP30P140 U212 ( .I(n906), .Z(o_data_bus[172]) );
  BUFFD12BWP30P140 U213 ( .I(n905), .Z(o_data_bus[173]) );
  BUFFD12BWP30P140 U214 ( .I(n904), .Z(o_data_bus[174]) );
  BUFFD12BWP30P140 U215 ( .I(n903), .Z(o_data_bus[175]) );
  BUFFD12BWP30P140 U216 ( .I(n902), .Z(o_data_bus[176]) );
  BUFFD12BWP30P140 U217 ( .I(n901), .Z(o_data_bus[177]) );
  BUFFD12BWP30P140 U218 ( .I(n900), .Z(o_data_bus[178]) );
  BUFFD12BWP30P140 U219 ( .I(n899), .Z(o_data_bus[179]) );
  BUFFD12BWP30P140 U220 ( .I(n898), .Z(o_data_bus[180]) );
  BUFFD12BWP30P140 U221 ( .I(n897), .Z(o_data_bus[181]) );
  BUFFD12BWP30P140 U222 ( .I(n896), .Z(o_data_bus[182]) );
  BUFFD12BWP30P140 U223 ( .I(n895), .Z(o_data_bus[183]) );
  BUFFD12BWP30P140 U224 ( .I(n894), .Z(o_data_bus[184]) );
  BUFFD12BWP30P140 U225 ( .I(n893), .Z(o_data_bus[185]) );
  BUFFD12BWP30P140 U226 ( .I(n892), .Z(o_data_bus[186]) );
  BUFFD12BWP30P140 U227 ( .I(n891), .Z(o_data_bus[187]) );
  BUFFD12BWP30P140 U228 ( .I(n890), .Z(o_data_bus[188]) );
  BUFFD12BWP30P140 U229 ( .I(n889), .Z(o_data_bus[189]) );
  BUFFD12BWP30P140 U230 ( .I(n888), .Z(o_data_bus[190]) );
  BUFFD12BWP30P140 U231 ( .I(n887), .Z(o_data_bus[191]) );
  BUFFD12BWP30P140 U232 ( .I(n886), .Z(o_data_bus[192]) );
  BUFFD12BWP30P140 U233 ( .I(n885), .Z(o_data_bus[193]) );
  BUFFD12BWP30P140 U234 ( .I(n884), .Z(o_data_bus[194]) );
  BUFFD12BWP30P140 U235 ( .I(n883), .Z(o_data_bus[195]) );
  BUFFD12BWP30P140 U236 ( .I(n882), .Z(o_data_bus[196]) );
  BUFFD12BWP30P140 U237 ( .I(n881), .Z(o_data_bus[197]) );
  BUFFD12BWP30P140 U238 ( .I(n880), .Z(o_data_bus[198]) );
  BUFFD12BWP30P140 U239 ( .I(n879), .Z(o_data_bus[199]) );
  BUFFD12BWP30P140 U240 ( .I(n878), .Z(o_data_bus[200]) );
  BUFFD12BWP30P140 U241 ( .I(n877), .Z(o_data_bus[201]) );
  BUFFD12BWP30P140 U242 ( .I(n876), .Z(o_data_bus[202]) );
  BUFFD12BWP30P140 U243 ( .I(n875), .Z(o_data_bus[203]) );
  BUFFD12BWP30P140 U244 ( .I(n874), .Z(o_data_bus[204]) );
  BUFFD12BWP30P140 U245 ( .I(n873), .Z(o_data_bus[205]) );
  BUFFD12BWP30P140 U246 ( .I(n872), .Z(o_data_bus[206]) );
  BUFFD12BWP30P140 U247 ( .I(n871), .Z(o_data_bus[207]) );
  BUFFD12BWP30P140 U248 ( .I(n870), .Z(o_data_bus[208]) );
  BUFFD12BWP30P140 U249 ( .I(n869), .Z(o_data_bus[209]) );
  BUFFD12BWP30P140 U250 ( .I(n868), .Z(o_data_bus[210]) );
  BUFFD12BWP30P140 U251 ( .I(n867), .Z(o_data_bus[211]) );
  BUFFD12BWP30P140 U252 ( .I(n866), .Z(o_data_bus[212]) );
  BUFFD12BWP30P140 U253 ( .I(n865), .Z(o_data_bus[213]) );
  BUFFD12BWP30P140 U254 ( .I(n864), .Z(o_data_bus[214]) );
  BUFFD12BWP30P140 U255 ( .I(n863), .Z(o_data_bus[215]) );
  BUFFD12BWP30P140 U256 ( .I(n862), .Z(o_data_bus[216]) );
  BUFFD12BWP30P140 U257 ( .I(n861), .Z(o_data_bus[217]) );
  BUFFD12BWP30P140 U258 ( .I(n860), .Z(o_data_bus[218]) );
  BUFFD12BWP30P140 U259 ( .I(n859), .Z(o_data_bus[219]) );
  BUFFD12BWP30P140 U260 ( .I(n858), .Z(o_data_bus[220]) );
  BUFFD12BWP30P140 U261 ( .I(n857), .Z(o_data_bus[221]) );
  BUFFD12BWP30P140 U262 ( .I(n856), .Z(o_data_bus[222]) );
  BUFFD12BWP30P140 U263 ( .I(n855), .Z(o_data_bus[223]) );
  BUFFD12BWP30P140 U264 ( .I(n854), .Z(o_data_bus[224]) );
  BUFFD12BWP30P140 U265 ( .I(n853), .Z(o_data_bus[225]) );
  BUFFD12BWP30P140 U266 ( .I(n852), .Z(o_data_bus[226]) );
  BUFFD12BWP30P140 U267 ( .I(n851), .Z(o_data_bus[227]) );
  BUFFD12BWP30P140 U268 ( .I(n850), .Z(o_data_bus[228]) );
  BUFFD12BWP30P140 U269 ( .I(n849), .Z(o_data_bus[229]) );
  BUFFD12BWP30P140 U270 ( .I(n848), .Z(o_data_bus[230]) );
  BUFFD12BWP30P140 U271 ( .I(n847), .Z(o_data_bus[231]) );
  BUFFD12BWP30P140 U272 ( .I(n846), .Z(o_data_bus[232]) );
  BUFFD12BWP30P140 U273 ( .I(n845), .Z(o_data_bus[233]) );
  BUFFD12BWP30P140 U274 ( .I(n844), .Z(o_data_bus[234]) );
  BUFFD12BWP30P140 U275 ( .I(n843), .Z(o_data_bus[235]) );
  BUFFD12BWP30P140 U276 ( .I(n842), .Z(o_data_bus[236]) );
  BUFFD12BWP30P140 U277 ( .I(n841), .Z(o_data_bus[237]) );
  BUFFD12BWP30P140 U278 ( .I(n840), .Z(o_data_bus[238]) );
  BUFFD12BWP30P140 U279 ( .I(n839), .Z(o_data_bus[239]) );
  BUFFD12BWP30P140 U280 ( .I(n838), .Z(o_data_bus[240]) );
  BUFFD12BWP30P140 U281 ( .I(n837), .Z(o_data_bus[241]) );
  BUFFD12BWP30P140 U282 ( .I(n836), .Z(o_data_bus[242]) );
  BUFFD12BWP30P140 U283 ( .I(n835), .Z(o_data_bus[243]) );
  BUFFD12BWP30P140 U284 ( .I(n834), .Z(o_data_bus[244]) );
  BUFFD12BWP30P140 U285 ( .I(n833), .Z(o_data_bus[245]) );
  BUFFD12BWP30P140 U286 ( .I(n832), .Z(o_data_bus[246]) );
  BUFFD12BWP30P140 U287 ( .I(n831), .Z(o_data_bus[247]) );
  BUFFD12BWP30P140 U288 ( .I(n830), .Z(o_data_bus[248]) );
  BUFFD12BWP30P140 U289 ( .I(n829), .Z(o_data_bus[249]) );
  BUFFD12BWP30P140 U290 ( .I(n828), .Z(o_data_bus[250]) );
  BUFFD12BWP30P140 U291 ( .I(n827), .Z(o_data_bus[251]) );
  BUFFD12BWP30P140 U292 ( .I(n826), .Z(o_data_bus[252]) );
  BUFFD12BWP30P140 U293 ( .I(n825), .Z(o_data_bus[253]) );
  BUFFD12BWP30P140 U294 ( .I(n824), .Z(o_data_bus[254]) );
  BUFFD12BWP30P140 U295 ( .I(n823), .Z(o_data_bus[255]) );
  BUFFD12BWP30P140 U296 ( .I(n822), .Z(o_data_bus[256]) );
  BUFFD12BWP30P140 U297 ( .I(n821), .Z(o_data_bus[257]) );
  BUFFD12BWP30P140 U298 ( .I(n820), .Z(o_data_bus[258]) );
  BUFFD12BWP30P140 U299 ( .I(n819), .Z(o_data_bus[259]) );
  BUFFD12BWP30P140 U300 ( .I(n818), .Z(o_data_bus[260]) );
  BUFFD12BWP30P140 U301 ( .I(n817), .Z(o_data_bus[261]) );
  BUFFD12BWP30P140 U302 ( .I(n816), .Z(o_data_bus[262]) );
  BUFFD12BWP30P140 U303 ( .I(n815), .Z(o_data_bus[263]) );
  BUFFD12BWP30P140 U304 ( .I(n814), .Z(o_data_bus[264]) );
  BUFFD12BWP30P140 U305 ( .I(n813), .Z(o_data_bus[265]) );
  BUFFD12BWP30P140 U306 ( .I(n812), .Z(o_data_bus[266]) );
  BUFFD12BWP30P140 U307 ( .I(n811), .Z(o_data_bus[267]) );
  BUFFD12BWP30P140 U308 ( .I(n810), .Z(o_data_bus[268]) );
  BUFFD12BWP30P140 U309 ( .I(n809), .Z(o_data_bus[269]) );
  BUFFD12BWP30P140 U310 ( .I(n808), .Z(o_data_bus[270]) );
  BUFFD12BWP30P140 U311 ( .I(n807), .Z(o_data_bus[271]) );
  BUFFD12BWP30P140 U312 ( .I(n806), .Z(o_data_bus[272]) );
  BUFFD12BWP30P140 U313 ( .I(n805), .Z(o_data_bus[273]) );
  BUFFD12BWP30P140 U314 ( .I(n804), .Z(o_data_bus[274]) );
  BUFFD12BWP30P140 U315 ( .I(n803), .Z(o_data_bus[275]) );
  BUFFD12BWP30P140 U316 ( .I(n802), .Z(o_data_bus[276]) );
  BUFFD12BWP30P140 U317 ( .I(n801), .Z(o_data_bus[277]) );
  BUFFD12BWP30P140 U318 ( .I(n800), .Z(o_data_bus[278]) );
  BUFFD12BWP30P140 U319 ( .I(n799), .Z(o_data_bus[279]) );
  BUFFD12BWP30P140 U320 ( .I(n798), .Z(o_data_bus[280]) );
  BUFFD12BWP30P140 U321 ( .I(n797), .Z(o_data_bus[281]) );
  BUFFD12BWP30P140 U322 ( .I(n796), .Z(o_data_bus[282]) );
  BUFFD12BWP30P140 U323 ( .I(n795), .Z(o_data_bus[283]) );
  BUFFD12BWP30P140 U324 ( .I(n794), .Z(o_data_bus[284]) );
  BUFFD12BWP30P140 U325 ( .I(n793), .Z(o_data_bus[285]) );
  BUFFD12BWP30P140 U326 ( .I(n792), .Z(o_data_bus[286]) );
  BUFFD12BWP30P140 U327 ( .I(n791), .Z(o_data_bus[287]) );
  BUFFD12BWP30P140 U328 ( .I(n790), .Z(o_data_bus[288]) );
  BUFFD12BWP30P140 U329 ( .I(n789), .Z(o_data_bus[289]) );
  BUFFD12BWP30P140 U330 ( .I(n788), .Z(o_data_bus[290]) );
  BUFFD12BWP30P140 U331 ( .I(n787), .Z(o_data_bus[291]) );
  BUFFD12BWP30P140 U332 ( .I(n786), .Z(o_data_bus[292]) );
  BUFFD12BWP30P140 U333 ( .I(n785), .Z(o_data_bus[293]) );
  BUFFD12BWP30P140 U334 ( .I(n784), .Z(o_data_bus[294]) );
  BUFFD12BWP30P140 U335 ( .I(n783), .Z(o_data_bus[295]) );
  BUFFD12BWP30P140 U336 ( .I(n782), .Z(o_data_bus[296]) );
  BUFFD12BWP30P140 U337 ( .I(n781), .Z(o_data_bus[297]) );
  BUFFD12BWP30P140 U338 ( .I(n780), .Z(o_data_bus[298]) );
  BUFFD12BWP30P140 U339 ( .I(n779), .Z(o_data_bus[299]) );
  BUFFD12BWP30P140 U340 ( .I(n778), .Z(o_data_bus[300]) );
  BUFFD12BWP30P140 U341 ( .I(n777), .Z(o_data_bus[301]) );
  BUFFD12BWP30P140 U342 ( .I(n776), .Z(o_data_bus[302]) );
  BUFFD12BWP30P140 U343 ( .I(n775), .Z(o_data_bus[303]) );
  BUFFD12BWP30P140 U344 ( .I(n774), .Z(o_data_bus[304]) );
  BUFFD12BWP30P140 U345 ( .I(n773), .Z(o_data_bus[305]) );
  BUFFD12BWP30P140 U346 ( .I(n772), .Z(o_data_bus[306]) );
  BUFFD12BWP30P140 U347 ( .I(n771), .Z(o_data_bus[307]) );
  BUFFD12BWP30P140 U348 ( .I(n770), .Z(o_data_bus[308]) );
  BUFFD12BWP30P140 U349 ( .I(n769), .Z(o_data_bus[309]) );
  BUFFD12BWP30P140 U350 ( .I(n768), .Z(o_data_bus[310]) );
  BUFFD12BWP30P140 U351 ( .I(n767), .Z(o_data_bus[311]) );
  BUFFD12BWP30P140 U352 ( .I(n766), .Z(o_data_bus[312]) );
  BUFFD12BWP30P140 U353 ( .I(n765), .Z(o_data_bus[313]) );
  BUFFD12BWP30P140 U354 ( .I(n764), .Z(o_data_bus[314]) );
  BUFFD12BWP30P140 U355 ( .I(n763), .Z(o_data_bus[315]) );
  BUFFD12BWP30P140 U356 ( .I(n762), .Z(o_data_bus[316]) );
  BUFFD12BWP30P140 U357 ( .I(n761), .Z(o_data_bus[317]) );
  BUFFD12BWP30P140 U358 ( .I(n760), .Z(o_data_bus[318]) );
  BUFFD12BWP30P140 U359 ( .I(n759), .Z(o_data_bus[319]) );
  BUFFD12BWP30P140 U360 ( .I(n758), .Z(o_data_bus[320]) );
  BUFFD12BWP30P140 U361 ( .I(n757), .Z(o_data_bus[321]) );
  BUFFD12BWP30P140 U362 ( .I(n756), .Z(o_data_bus[322]) );
  BUFFD12BWP30P140 U363 ( .I(n755), .Z(o_data_bus[323]) );
  BUFFD12BWP30P140 U364 ( .I(n754), .Z(o_data_bus[324]) );
  BUFFD12BWP30P140 U365 ( .I(n753), .Z(o_data_bus[325]) );
  BUFFD12BWP30P140 U366 ( .I(n752), .Z(o_data_bus[326]) );
  BUFFD12BWP30P140 U367 ( .I(n751), .Z(o_data_bus[327]) );
  BUFFD12BWP30P140 U368 ( .I(n750), .Z(o_data_bus[328]) );
  BUFFD12BWP30P140 U369 ( .I(n749), .Z(o_data_bus[329]) );
  BUFFD12BWP30P140 U370 ( .I(n748), .Z(o_data_bus[330]) );
  BUFFD12BWP30P140 U371 ( .I(n747), .Z(o_data_bus[331]) );
  BUFFD12BWP30P140 U372 ( .I(n746), .Z(o_data_bus[332]) );
  BUFFD12BWP30P140 U373 ( .I(n745), .Z(o_data_bus[333]) );
  BUFFD12BWP30P140 U374 ( .I(n744), .Z(o_data_bus[334]) );
  BUFFD12BWP30P140 U375 ( .I(n743), .Z(o_data_bus[335]) );
  BUFFD12BWP30P140 U376 ( .I(n742), .Z(o_data_bus[336]) );
  BUFFD12BWP30P140 U377 ( .I(n741), .Z(o_data_bus[337]) );
  BUFFD12BWP30P140 U378 ( .I(n740), .Z(o_data_bus[338]) );
  BUFFD12BWP30P140 U379 ( .I(n739), .Z(o_data_bus[339]) );
  BUFFD12BWP30P140 U380 ( .I(n738), .Z(o_data_bus[340]) );
  BUFFD12BWP30P140 U381 ( .I(n737), .Z(o_data_bus[341]) );
  BUFFD12BWP30P140 U382 ( .I(n736), .Z(o_data_bus[342]) );
  BUFFD12BWP30P140 U383 ( .I(n735), .Z(o_data_bus[343]) );
  BUFFD12BWP30P140 U384 ( .I(n734), .Z(o_data_bus[344]) );
  BUFFD12BWP30P140 U385 ( .I(n733), .Z(o_data_bus[345]) );
  BUFFD12BWP30P140 U386 ( .I(n732), .Z(o_data_bus[346]) );
  BUFFD12BWP30P140 U387 ( .I(n731), .Z(o_data_bus[347]) );
  BUFFD12BWP30P140 U388 ( .I(n730), .Z(o_data_bus[348]) );
  BUFFD12BWP30P140 U389 ( .I(n729), .Z(o_data_bus[349]) );
  BUFFD12BWP30P140 U390 ( .I(n728), .Z(o_data_bus[350]) );
  BUFFD12BWP30P140 U391 ( .I(n727), .Z(o_data_bus[351]) );
  BUFFD12BWP30P140 U392 ( .I(n726), .Z(o_data_bus[352]) );
  BUFFD12BWP30P140 U393 ( .I(n725), .Z(o_data_bus[353]) );
  BUFFD12BWP30P140 U394 ( .I(n724), .Z(o_data_bus[354]) );
  BUFFD12BWP30P140 U395 ( .I(n723), .Z(o_data_bus[355]) );
  BUFFD12BWP30P140 U396 ( .I(n722), .Z(o_data_bus[356]) );
  BUFFD12BWP30P140 U397 ( .I(n721), .Z(o_data_bus[357]) );
  BUFFD12BWP30P140 U398 ( .I(n720), .Z(o_data_bus[358]) );
  BUFFD12BWP30P140 U399 ( .I(n719), .Z(o_data_bus[359]) );
  BUFFD12BWP30P140 U400 ( .I(n718), .Z(o_data_bus[360]) );
  BUFFD12BWP30P140 U401 ( .I(n717), .Z(o_data_bus[361]) );
  BUFFD12BWP30P140 U402 ( .I(n716), .Z(o_data_bus[362]) );
  BUFFD12BWP30P140 U403 ( .I(n715), .Z(o_data_bus[363]) );
  BUFFD12BWP30P140 U404 ( .I(n714), .Z(o_data_bus[364]) );
  BUFFD12BWP30P140 U405 ( .I(n713), .Z(o_data_bus[365]) );
  BUFFD12BWP30P140 U406 ( .I(n712), .Z(o_data_bus[366]) );
  BUFFD12BWP30P140 U407 ( .I(n711), .Z(o_data_bus[367]) );
  BUFFD12BWP30P140 U408 ( .I(n710), .Z(o_data_bus[368]) );
  BUFFD12BWP30P140 U409 ( .I(n709), .Z(o_data_bus[369]) );
  BUFFD12BWP30P140 U410 ( .I(n708), .Z(o_data_bus[370]) );
  BUFFD12BWP30P140 U411 ( .I(n707), .Z(o_data_bus[371]) );
  BUFFD12BWP30P140 U412 ( .I(n706), .Z(o_data_bus[372]) );
  BUFFD12BWP30P140 U413 ( .I(n705), .Z(o_data_bus[373]) );
  BUFFD12BWP30P140 U414 ( .I(n704), .Z(o_data_bus[374]) );
  BUFFD12BWP30P140 U415 ( .I(n703), .Z(o_data_bus[375]) );
  BUFFD12BWP30P140 U416 ( .I(n702), .Z(o_data_bus[376]) );
  BUFFD12BWP30P140 U417 ( .I(n701), .Z(o_data_bus[377]) );
  BUFFD12BWP30P140 U418 ( .I(n700), .Z(o_data_bus[378]) );
  BUFFD12BWP30P140 U419 ( .I(n699), .Z(o_data_bus[379]) );
  BUFFD12BWP30P140 U420 ( .I(n698), .Z(o_data_bus[380]) );
  BUFFD12BWP30P140 U421 ( .I(n697), .Z(o_data_bus[381]) );
  BUFFD12BWP30P140 U422 ( .I(n696), .Z(o_data_bus[382]) );
  BUFFD12BWP30P140 U423 ( .I(n695), .Z(o_data_bus[383]) );
  BUFFD12BWP30P140 U424 ( .I(n694), .Z(o_data_bus[384]) );
  BUFFD12BWP30P140 U425 ( .I(n693), .Z(o_data_bus[385]) );
  BUFFD12BWP30P140 U426 ( .I(n692), .Z(o_data_bus[386]) );
  BUFFD12BWP30P140 U427 ( .I(n691), .Z(o_data_bus[387]) );
  BUFFD12BWP30P140 U428 ( .I(n690), .Z(o_data_bus[388]) );
  BUFFD12BWP30P140 U429 ( .I(n689), .Z(o_data_bus[389]) );
  BUFFD12BWP30P140 U430 ( .I(n688), .Z(o_data_bus[390]) );
  BUFFD12BWP30P140 U431 ( .I(n687), .Z(o_data_bus[391]) );
  BUFFD12BWP30P140 U432 ( .I(n686), .Z(o_data_bus[392]) );
  BUFFD12BWP30P140 U433 ( .I(n685), .Z(o_data_bus[393]) );
  BUFFD12BWP30P140 U434 ( .I(n684), .Z(o_data_bus[394]) );
  BUFFD12BWP30P140 U435 ( .I(n683), .Z(o_data_bus[395]) );
  BUFFD12BWP30P140 U436 ( .I(n682), .Z(o_data_bus[396]) );
  BUFFD12BWP30P140 U437 ( .I(n681), .Z(o_data_bus[397]) );
  BUFFD12BWP30P140 U438 ( .I(n680), .Z(o_data_bus[398]) );
  BUFFD12BWP30P140 U439 ( .I(n679), .Z(o_data_bus[399]) );
  BUFFD12BWP30P140 U440 ( .I(n678), .Z(o_data_bus[400]) );
  BUFFD12BWP30P140 U441 ( .I(n677), .Z(o_data_bus[401]) );
  BUFFD12BWP30P140 U442 ( .I(n676), .Z(o_data_bus[402]) );
  BUFFD12BWP30P140 U443 ( .I(n675), .Z(o_data_bus[403]) );
  BUFFD12BWP30P140 U444 ( .I(n674), .Z(o_data_bus[404]) );
  BUFFD12BWP30P140 U445 ( .I(n673), .Z(o_data_bus[405]) );
  BUFFD12BWP30P140 U446 ( .I(n672), .Z(o_data_bus[406]) );
  BUFFD12BWP30P140 U447 ( .I(n671), .Z(o_data_bus[407]) );
  BUFFD12BWP30P140 U448 ( .I(n670), .Z(o_data_bus[408]) );
  BUFFD12BWP30P140 U449 ( .I(n669), .Z(o_data_bus[409]) );
  BUFFD12BWP30P140 U450 ( .I(n668), .Z(o_data_bus[410]) );
  BUFFD12BWP30P140 U451 ( .I(n667), .Z(o_data_bus[411]) );
  BUFFD12BWP30P140 U452 ( .I(n666), .Z(o_data_bus[412]) );
  BUFFD12BWP30P140 U453 ( .I(n665), .Z(o_data_bus[413]) );
  BUFFD12BWP30P140 U454 ( .I(n664), .Z(o_data_bus[414]) );
  BUFFD12BWP30P140 U455 ( .I(n663), .Z(o_data_bus[415]) );
  BUFFD12BWP30P140 U456 ( .I(n662), .Z(o_data_bus[416]) );
  BUFFD12BWP30P140 U457 ( .I(n661), .Z(o_data_bus[417]) );
  BUFFD12BWP30P140 U458 ( .I(n660), .Z(o_data_bus[418]) );
  BUFFD12BWP30P140 U459 ( .I(n659), .Z(o_data_bus[419]) );
  BUFFD12BWP30P140 U460 ( .I(n658), .Z(o_data_bus[420]) );
  BUFFD12BWP30P140 U461 ( .I(n657), .Z(o_data_bus[421]) );
  BUFFD12BWP30P140 U462 ( .I(n656), .Z(o_data_bus[422]) );
  BUFFD12BWP30P140 U463 ( .I(n655), .Z(o_data_bus[423]) );
  BUFFD12BWP30P140 U464 ( .I(n654), .Z(o_data_bus[424]) );
  BUFFD12BWP30P140 U465 ( .I(n653), .Z(o_data_bus[425]) );
  BUFFD12BWP30P140 U466 ( .I(n652), .Z(o_data_bus[426]) );
  BUFFD12BWP30P140 U467 ( .I(n651), .Z(o_data_bus[427]) );
  BUFFD12BWP30P140 U468 ( .I(n650), .Z(o_data_bus[428]) );
  BUFFD12BWP30P140 U469 ( .I(n649), .Z(o_data_bus[429]) );
  BUFFD12BWP30P140 U470 ( .I(n648), .Z(o_data_bus[430]) );
  BUFFD12BWP30P140 U471 ( .I(n647), .Z(o_data_bus[431]) );
  BUFFD12BWP30P140 U472 ( .I(n646), .Z(o_data_bus[432]) );
  BUFFD12BWP30P140 U473 ( .I(n645), .Z(o_data_bus[433]) );
  BUFFD12BWP30P140 U474 ( .I(n644), .Z(o_data_bus[434]) );
  BUFFD12BWP30P140 U475 ( .I(n643), .Z(o_data_bus[435]) );
  BUFFD12BWP30P140 U476 ( .I(n642), .Z(o_data_bus[436]) );
  BUFFD12BWP30P140 U477 ( .I(n641), .Z(o_data_bus[437]) );
  BUFFD12BWP30P140 U478 ( .I(n640), .Z(o_data_bus[438]) );
  BUFFD12BWP30P140 U479 ( .I(n639), .Z(o_data_bus[439]) );
  BUFFD12BWP30P140 U480 ( .I(n638), .Z(o_data_bus[440]) );
  BUFFD12BWP30P140 U481 ( .I(n637), .Z(o_data_bus[441]) );
  BUFFD12BWP30P140 U482 ( .I(n636), .Z(o_data_bus[442]) );
  BUFFD12BWP30P140 U483 ( .I(n635), .Z(o_data_bus[443]) );
  BUFFD12BWP30P140 U484 ( .I(n634), .Z(o_data_bus[444]) );
  BUFFD12BWP30P140 U485 ( .I(n633), .Z(o_data_bus[445]) );
  BUFFD12BWP30P140 U486 ( .I(n632), .Z(o_data_bus[446]) );
  BUFFD12BWP30P140 U487 ( .I(n631), .Z(o_data_bus[447]) );
  BUFFD12BWP30P140 U488 ( .I(n630), .Z(o_data_bus[448]) );
  BUFFD12BWP30P140 U489 ( .I(n629), .Z(o_data_bus[449]) );
  BUFFD12BWP30P140 U490 ( .I(n628), .Z(o_data_bus[450]) );
  BUFFD12BWP30P140 U491 ( .I(n627), .Z(o_data_bus[451]) );
  BUFFD12BWP30P140 U492 ( .I(n626), .Z(o_data_bus[452]) );
  BUFFD12BWP30P140 U493 ( .I(n624), .Z(o_data_bus[454]) );
  BUFFD12BWP30P140 U494 ( .I(n622), .Z(o_data_bus[456]) );
  BUFFD12BWP30P140 U495 ( .I(n621), .Z(o_data_bus[457]) );
  BUFFD12BWP30P140 U496 ( .I(n620), .Z(o_data_bus[458]) );
  BUFFD12BWP30P140 U497 ( .I(n619), .Z(o_data_bus[459]) );
  BUFFD12BWP30P140 U498 ( .I(n618), .Z(o_data_bus[460]) );
  BUFFD12BWP30P140 U499 ( .I(n617), .Z(o_data_bus[461]) );
  BUFFD12BWP30P140 U500 ( .I(n616), .Z(o_data_bus[462]) );
  BUFFD12BWP30P140 U501 ( .I(n615), .Z(o_data_bus[463]) );
  BUFFD12BWP30P140 U502 ( .I(n614), .Z(o_data_bus[464]) );
  BUFFD12BWP30P140 U503 ( .I(n613), .Z(o_data_bus[465]) );
  BUFFD12BWP30P140 U504 ( .I(n612), .Z(o_data_bus[466]) );
  BUFFD12BWP30P140 U505 ( .I(n611), .Z(o_data_bus[467]) );
  BUFFD12BWP30P140 U506 ( .I(n610), .Z(o_data_bus[468]) );
  BUFFD12BWP30P140 U507 ( .I(n609), .Z(o_data_bus[469]) );
  BUFFD12BWP30P140 U508 ( .I(n607), .Z(o_data_bus[471]) );
  BUFFD12BWP30P140 U509 ( .I(n605), .Z(o_data_bus[473]) );
  BUFFD12BWP30P140 U510 ( .I(n603), .Z(o_data_bus[475]) );
  BUFFD12BWP30P140 U511 ( .I(n601), .Z(o_data_bus[477]) );
  BUFFD12BWP30P140 U512 ( .I(n599), .Z(o_data_bus[479]) );
  BUFFD12BWP30P140 U513 ( .I(n598), .Z(o_data_bus[480]) );
  BUFFD12BWP30P140 U514 ( .I(n597), .Z(o_data_bus[481]) );
  BUFFD12BWP30P140 U515 ( .I(n596), .Z(o_data_bus[482]) );
  BUFFD12BWP30P140 U516 ( .I(n595), .Z(o_data_bus[483]) );
  BUFFD12BWP30P140 U517 ( .I(n594), .Z(o_data_bus[484]) );
  BUFFD12BWP30P140 U518 ( .I(n593), .Z(o_data_bus[485]) );
  BUFFD12BWP30P140 U519 ( .I(n592), .Z(o_data_bus[486]) );
  BUFFD12BWP30P140 U520 ( .I(n591), .Z(o_data_bus[487]) );
  BUFFD12BWP30P140 U521 ( .I(n590), .Z(o_data_bus[488]) );
  BUFFD12BWP30P140 U522 ( .I(n589), .Z(o_data_bus[489]) );
  BUFFD12BWP30P140 U523 ( .I(n588), .Z(o_data_bus[490]) );
  BUFFD12BWP30P140 U524 ( .I(n587), .Z(o_data_bus[491]) );
  BUFFD12BWP30P140 U525 ( .I(n586), .Z(o_data_bus[492]) );
  BUFFD12BWP30P140 U526 ( .I(n585), .Z(o_data_bus[493]) );
  BUFFD12BWP30P140 U527 ( .I(n584), .Z(o_data_bus[494]) );
  BUFFD12BWP30P140 U528 ( .I(n583), .Z(o_data_bus[495]) );
  BUFFD12BWP30P140 U529 ( .I(n582), .Z(o_data_bus[496]) );
  BUFFD12BWP30P140 U530 ( .I(n581), .Z(o_data_bus[497]) );
  BUFFD12BWP30P140 U531 ( .I(n580), .Z(o_data_bus[498]) );
  BUFFD12BWP30P140 U532 ( .I(n579), .Z(o_data_bus[499]) );
  BUFFD12BWP30P140 U533 ( .I(n578), .Z(o_data_bus[500]) );
  BUFFD12BWP30P140 U534 ( .I(n577), .Z(o_data_bus[501]) );
  BUFFD12BWP30P140 U535 ( .I(n576), .Z(o_data_bus[502]) );
  BUFFD12BWP30P140 U536 ( .I(n575), .Z(o_data_bus[503]) );
  BUFFD12BWP30P140 U537 ( .I(n574), .Z(o_data_bus[504]) );
  BUFFD12BWP30P140 U538 ( .I(n573), .Z(o_data_bus[505]) );
  BUFFD12BWP30P140 U539 ( .I(n572), .Z(o_data_bus[506]) );
  BUFFD12BWP30P140 U540 ( .I(n571), .Z(o_data_bus[507]) );
  BUFFD12BWP30P140 U541 ( .I(n570), .Z(o_data_bus[508]) );
  BUFFD12BWP30P140 U542 ( .I(n569), .Z(o_data_bus[509]) );
  BUFFD12BWP30P140 U543 ( .I(n568), .Z(o_data_bus[510]) );
  BUFFD12BWP30P140 U544 ( .I(n567), .Z(o_data_bus[511]) );
  BUFFD12BWP30P140 U545 ( .I(n566), .Z(o_valid[0]) );
  BUFFD12BWP30P140 U546 ( .I(n564), .Z(o_valid[2]) );
  BUFFD12BWP30P140 U547 ( .I(n562), .Z(o_valid[4]) );
  BUFFD12BWP30P140 U548 ( .I(n560), .Z(o_valid[6]) );
  BUFFD12BWP30P140 U549 ( .I(n558), .Z(o_valid[8]) );
  BUFFD12BWP30P140 U550 ( .I(n556), .Z(o_valid[10]) );
  BUFFD12BWP30P140 U551 ( .I(n554), .Z(o_valid[12]) );
  BUFFD12BWP30P140 U552 ( .I(n552), .Z(o_valid[14]) );
endmodule

