`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////////////////////
// Company: Gatech	
// Engineer: Mandovi Mukherjee
// 
// Create Date: 03/31/2021 
// System Name: accelerator
// Module Name: global controller
// Project Name: ARION DRBE
// Description: global controller top module 
// Dependencies:
// Additional Comments: 
/////////////////////////////////////////////////////////////////////////////////////////////////////

module global_controller(CLK, reset, boot_up, table_parse, input_valid, glob_scen_noc_input_valid, delay_matrix_element, obj_id_element,from_glob_prefetch_start,  from_glob_prefetch_dest,  scenario_update, local_controller_id, tapping_loc_packet);

    // parameter
    	parameter N_sample = 256;
	parameter datawidth = 16;
	parameter address_vector_width = 8; //can be 200 or 8: 8 for small tapeout
	parameter id_width = 4; // 16 local controllers in subscaled system
	parameter sample_address_width = 8; /// assuming 256 words: needs to change if arrangement is different
	parameter packet_width = 2*datawidth + address_vector_width;
	parameter delay_length = 12; // log(id_width*N_sample)
	parameter obj_id_width = 3; // log(N_obj)
	parameter tapping_loc_packet_width = sample_address_width + obj_id_width;
//=== IO Ports ===//


    // input
    	input CLK; // system clock, generated by VCO
	input reset;
	input boot_up;
	input table_parse;
	input input_valid;
	input glob_scen_noc_input_valid;
	input [delay_length - 1:0] delay_matrix_element;
	input [obj_id_width - 1:0] obj_id_element;
	input scenario_update;



    // output
	output [address_vector_width - 1:0] from_glob_prefetch_dest;
	output [sample_address_width - 1:0] from_glob_prefetch_start;
	output [id_width - 1:0] local_controller_id;
	output [tapping_loc_packet_width - 1:0] tapping_loc_packet;

//////////// internal status regs/signals //////////////////////////////////
	wire [address_vector_width - 1:0] calc_glob_prefetch_dest;

	wire [sample_address_width - 1:0] calc_glob_controller_delay;
        //wire [sample_address_width - 1:0] calc_glob_prefetch_stop;

///////////////////////////////////////////////////////////////////////////////    

////////// logic part ///////////////////////////////////////////////////////  

	assign from_glob_prefetch_start = calc_glob_controller_delay;
	assign from_glob_prefetch_dest = calc_glob_prefetch_dest;


////////////sequential logic
//
//

	 
	 
 table_parse_engine dut_parse_engine (.CLK(CLK), .reset(reset), .boot_up(boot_up), .table_parse(table_parse), .input_valid(input_valid), .glob_scen_noc_input_valid(glob_scen_noc_input_valid), .delay_matrix_element(delay_matrix_element), .obj_id_element(obj_id_element), .local_controller_id(local_controller_id), .calc_glob_controller_delay(calc_glob_controller_delay), .calc_glob_dest_addr(calc_glob_prefetch_dest),  .tapping_loc_packet(tapping_loc_packet), .scenario_update(scenario_update));

   
endmodule
    
