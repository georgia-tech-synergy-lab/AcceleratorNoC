module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_0 (
	CLK_clone24, 
	rst, 
	i_valid, 
	i_data_bus, 
	o_valid, 
	o_data_bus, 
	i_en, 
	CLK_clone28, 
	CLK_clone11, 
	CLK_clone30, 
	CLK_clone39, 
	CLK_clone22, 
	CLK_clone21, 
	CLK_clone33, 
	CLK_clone20, 
	CLK_clone18, 
	CLK_clone17, 
	CLK_clone16, 
	CLK_clone15, 
	CLK_clone13, 
	CLK_clone10, 
	CLK_clone12, 
	CLK_clone23, 
	CLK_clone9, 
	CLK_clone8, 
	CLK_clone7, 
	CLK_clone6, 
	CLK_clone5, 
	CLK_clone19, 
	CLK_clone4, 
	CLK_clone3, 
	CLK_clone14, 
	CLK_clone2, 
	CLK_clone1, 
	CLK, 
	CLK_clone44, 
	CLK_clone43, 
	CLK_clone41, 
	CLK_clone40, 
	CLK_clone42, 
	CLK_clone38, 
	CLK_clone37, 
	CLK_clone36, 
	CLK_clone35, 
	CLK_clone34, 
	CLK_clone29, 
	CLK_clone32, 
	CLK_clone31, 
	CLK_clone27, 
	CLK_clone26, 
	CLK_clone25);
   input CLK_clone24;
   input rst;
   input [0:0] i_valid;
   input [31:0] i_data_bus;
   output [7:0] o_valid;
   output [255:0] o_data_bus;
   input i_en;
   input CLK_clone28;
   input CLK_clone11;
   input CLK_clone30;
   input CLK_clone39;
   input CLK_clone22;
   input CLK_clone21;
   input CLK_clone33;
   input CLK_clone20;
   input CLK_clone18;
   input CLK_clone17;
   input CLK_clone16;
   input CLK_clone15;
   input CLK_clone13;
   input CLK_clone10;
   input CLK_clone12;
   input CLK_clone23;
   input CLK_clone9;
   input CLK_clone8;
   input CLK_clone7;
   input CLK_clone6;
   input CLK_clone5;
   input CLK_clone19;
   input CLK_clone4;
   input CLK_clone3;
   input CLK_clone14;
   input CLK_clone2;
   input CLK_clone1;
   input CLK;
   input CLK_clone44;
   input CLK_clone43;
   input CLK_clone41;
   input CLK_clone40;
   input CLK_clone42;
   input CLK_clone38;
   input CLK_clone37;
   input CLK_clone36;
   input CLK_clone35;
   input CLK_clone34;
   input CLK_clone29;
   input CLK_clone32;
   input CLK_clone31;
   input CLK_clone27;
   input CLK_clone26;
   input CLK_clone25;

   // Internal wires
   wire FE_RN_144_0;
   wire FE_RN_143_0;
   wire FE_RN_142_0;
   wire FE_RN_125_0;
   wire FE_RN_124_0;
   wire FE_RN_123_0;
   wire FE_RN_122_0;
   wire FE_RN_120_0;
   wire FE_RN_116_0;
   wire FE_OCPN1470_n1;
   wire FE_OCPN1469_n1;
   wire FE_OCPN1468_n1;
   wire FE_OCPN1467_n1;
   wire FE_OCPN1466_n1;
   wire FE_OCPN1465_n1;
   wire FE_OCPN1464_n1;
   wire FE_OCPN1376_FE_OFN344_n1;
   wire FE_OCPN1375_FE_OFN344_n1;
   wire FE_OCPN1374_FE_OFN752_n1;
   wire FE_OFN344_n1;
   wire FE_OFN343_n1;
   wire FE_OFN342_n1;
   wire FE_OFN341_n1;
   wire wire_tree_level_0__i_valid_latch_0_;
   wire N3;
   wire N4;
   wire N5;
   wire N6;
   wire N7;
   wire N8;
   wire N9;
   wire N10;
   wire N11;
   wire N12;
   wire N13;
   wire N14;
   wire N15;
   wire N16;
   wire N17;
   wire N18;
   wire N19;
   wire N20;
   wire N21;
   wire N22;
   wire N23;
   wire N24;
   wire N25;
   wire N26;
   wire N27;
   wire N28;
   wire N29;
   wire N30;
   wire N31;
   wire N32;
   wire N33;
   wire N34;
   wire N35;
   wire N68;
   wire N69;
   wire N70;
   wire N71;
   wire N72;
   wire N73;
   wire N74;
   wire N75;
   wire N76;
   wire N77;
   wire N78;
   wire N79;
   wire N80;
   wire N81;
   wire N82;
   wire N83;
   wire N84;
   wire N85;
   wire N86;
   wire N87;
   wire N88;
   wire N89;
   wire N90;
   wire N91;
   wire N92;
   wire N93;
   wire N94;
   wire N95;
   wire N96;
   wire N97;
   wire N98;
   wire N99;
   wire N101;
   wire N134;
   wire N135;
   wire N136;
   wire N137;
   wire N138;
   wire N139;
   wire N140;
   wire N141;
   wire N142;
   wire N143;
   wire N144;
   wire N145;
   wire N146;
   wire N147;
   wire N148;
   wire N149;
   wire N150;
   wire N151;
   wire N152;
   wire N153;
   wire N154;
   wire N155;
   wire N156;
   wire N157;
   wire N158;
   wire N159;
   wire N160;
   wire N161;
   wire N162;
   wire N163;
   wire N164;
   wire N165;
   wire N167;
   wire N200;
   wire N201;
   wire N202;
   wire N203;
   wire N204;
   wire N205;
   wire N206;
   wire N207;
   wire N208;
   wire N209;
   wire N210;
   wire N211;
   wire N212;
   wire N213;
   wire N214;
   wire N215;
   wire N216;
   wire N217;
   wire N218;
   wire N219;
   wire N220;
   wire N221;
   wire N222;
   wire N223;
   wire N224;
   wire N225;
   wire N226;
   wire N227;
   wire N228;
   wire N229;
   wire N230;
   wire N231;
   wire N233;
   wire N266;
   wire N267;
   wire N268;
   wire N269;
   wire N270;
   wire N271;
   wire N272;
   wire N273;
   wire N274;
   wire N275;
   wire N276;
   wire N277;
   wire N278;
   wire N279;
   wire N280;
   wire N281;
   wire N282;
   wire N283;
   wire N284;
   wire N285;
   wire N286;
   wire N287;
   wire N288;
   wire N289;
   wire N290;
   wire N291;
   wire N292;
   wire N293;
   wire N294;
   wire N295;
   wire N296;
   wire N297;
   wire N299;
   wire N332;
   wire N333;
   wire N334;
   wire N335;
   wire N336;
   wire N337;
   wire N338;
   wire N339;
   wire N340;
   wire N341;
   wire N342;
   wire N343;
   wire N344;
   wire N345;
   wire N346;
   wire N347;
   wire N348;
   wire N349;
   wire N350;
   wire N351;
   wire N352;
   wire N353;
   wire N354;
   wire N355;
   wire N356;
   wire N357;
   wire N358;
   wire N359;
   wire N360;
   wire N361;
   wire N362;
   wire N363;
   wire N365;
   wire N398;
   wire N399;
   wire N400;
   wire N401;
   wire N402;
   wire N403;
   wire N404;
   wire N405;
   wire N406;
   wire N407;
   wire N408;
   wire N409;
   wire N410;
   wire N411;
   wire N412;
   wire N413;
   wire N414;
   wire N415;
   wire N416;
   wire N417;
   wire N418;
   wire N419;
   wire N420;
   wire N421;
   wire N422;
   wire N423;
   wire N424;
   wire N425;
   wire N426;
   wire N427;
   wire N428;
   wire N429;
   wire N431;
   wire N464;
   wire N465;
   wire N466;
   wire N467;
   wire N468;
   wire N469;
   wire N470;
   wire N471;
   wire N472;
   wire N473;
   wire N474;
   wire N475;
   wire N476;
   wire N477;
   wire N478;
   wire N479;
   wire N480;
   wire N481;
   wire N482;
   wire N483;
   wire N484;
   wire N485;
   wire N486;
   wire N487;
   wire N488;
   wire N489;
   wire N490;
   wire N491;
   wire N492;
   wire N493;
   wire N494;
   wire N495;
   wire N497;
   wire n1;
   wire [31:0] wire_tree_level_0__i_data_latch;
   wire [63:0] wire_tree_level_1__i_data_latch;
   wire [1:0] wire_tree_level_1__i_valid_latch;
   wire [127:0] wire_tree_level_2__i_data_latch;
   wire [3:0] wire_tree_level_2__i_valid_latch;

   INVD6BWP30P140LVT postctshold_FE_RC_336_0 (.I(i_data_bus[13]),
	.ZN(FE_RN_144_0));
   NR2OPTPAD8BWP30P140LVT postctshold_FE_RC_335_0 (.A1(FE_RN_144_0),
	.A2(FE_RN_143_0),
	.ZN(N16));
   INVD1BWP30P140LVT postctshold_FE_RC_334_0 (.I(FE_OCPN1376_FE_OFN344_n1),
	.ZN(FE_RN_143_0));
   INVD4BWP30P140LVT postctshold_FE_RC_332_0 (.I(i_data_bus[27]),
	.ZN(FE_RN_142_0));
   NR2OPTPAD8BWP30P140LVT postctshold_FE_RC_331_0 (.A1(FE_RN_142_0),
	.A2(FE_RN_125_0),
	.ZN(N30));
   INVD1BWP30P140LVT ccpot_FE_RC_285_0 (.I(FE_OCPN1376_FE_OFN344_n1),
	.ZN(FE_RN_125_0));
   INVD1BWP30P140LVT ccpot_FE_RC_283_0 (.I(FE_OCPN1376_FE_OFN344_n1),
	.ZN(FE_RN_124_0));
   INR2D16BWP30P140LVT ccpot_FE_RC_282_0 (.A1(i_data_bus[30]),
	.B1(FE_RN_124_0),
	.ZN(N33));
   INVD1BWP30P140LVT ccpot_FE_RC_281_0 (.I(FE_OCPN1376_FE_OFN344_n1),
	.ZN(FE_RN_123_0));
   INR2D16BWP30P140LVT ccpot_FE_RC_280_0 (.A1(i_valid[0]),
	.B1(FE_RN_123_0),
	.ZN(N35));
   INVD4BWP30P140LVT ccpot_FE_RC_279_0 (.I(i_data_bus[14]),
	.ZN(FE_RN_122_0));
   INR2D4BWP30P140LVT ccpot_FE_RC_278_0 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.B1(FE_RN_122_0),
	.ZN(N17));
   INVD4BWP30P140LVT ccpot_FE_RC_275_0 (.I(i_data_bus[22]),
	.ZN(FE_RN_120_0));
   INR2D4BWP30P140LVT ccpot_FE_RC_274_0 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.B1(FE_RN_120_0),
	.ZN(N25));
   INVD4BWP30P140LVT ccpot_FE_RC_264_0 (.I(i_data_bus[15]),
	.ZN(FE_RN_116_0));
   INR2D4BWP30P140LVT ccpot_FE_RC_263_0 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.B1(FE_RN_116_0),
	.ZN(N18));
   CKBD2BWP30P140LVT placeopt_FE_OCPC1874_n1 (.I(FE_OCPN1464_n1),
	.Z(FE_OCPN1470_n1));
   INVD2BWP30P140LVT placeopt_FE_OCPC1873_n1 (.I(FE_OFN342_n1),
	.ZN(FE_OCPN1469_n1));
   INVD1BWP30P140LVT placeopt_FE_OCPC1872_n1 (.I(FE_OFN342_n1),
	.ZN(FE_OCPN1468_n1));
   INVD2BWP30P140LVT placeopt_FE_OCPC1871_n1 (.I(FE_OFN342_n1),
	.ZN(FE_OCPN1467_n1));
   INVD2BWP30P140LVT placeopt_FE_OCPC1870_n1 (.I(FE_OFN342_n1),
	.ZN(FE_OCPN1466_n1));
   INVD1BWP30P140LVT placeopt_FE_OCPC1869_n1 (.I(FE_OFN342_n1),
	.ZN(FE_OCPN1465_n1));
   INVD3BWP30P140LVT placeopt_FE_OCPC1868_n1 (.I(FE_OFN342_n1),
	.ZN(FE_OCPN1464_n1));
   INVD2BWP30P140LVT placeopt_FE_OCPC1867_n1 (.I(FE_OFN342_n1),
	.ZN(FE_OFN341_n1));
   INVD2BWP30P140LVT placeopt_FE_OCPC1866_n1 (.I(FE_OFN342_n1),
	.ZN(FE_OFN343_n1));
   INVD2BWP30P140LVT placeopt_FE_OCPC1865_n1 (.I(FE_OFN342_n1),
	.ZN(FE_OFN344_n1));
   INVD9BWP30P140LVT placeopt_FE_OCPC1863_n1 (.I(n1),
	.ZN(FE_OFN342_n1));
   CKBD2BWP30P140LVT placeopt_FE_OCPC1757_FE_OFN344_n1 (.I(FE_OCPN1375_FE_OFN344_n1),
	.Z(FE_OCPN1376_FE_OFN344_n1));
   CKBD2BWP30P140LVT placeopt_FE_OCPC1756_FE_OFN344_n1 (.I(n1),
	.Z(FE_OCPN1375_FE_OFN344_n1));
   CKBD2BWP30P140LVT placeopt_FE_OCPC1755_FE_OFN752_n1 (.I(FE_OCPN1464_n1),
	.Z(FE_OCPN1374_FE_OFN752_n1));
   DFQD4BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ (.CP(CLK),
	.D(N35),
	.Q(wire_tree_level_0__i_valid_latch_0_));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ (.CP(CLK),
	.D(N34),
	.Q(wire_tree_level_0__i_data_latch[31]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ (.CP(CLK),
	.D(N33),
	.Q(wire_tree_level_0__i_data_latch[30]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ (.CP(CLK),
	.D(N32),
	.Q(wire_tree_level_0__i_data_latch[29]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ (.CP(CLK),
	.D(N31),
	.Q(wire_tree_level_0__i_data_latch[28]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ (.CP(CLK),
	.D(N30),
	.Q(wire_tree_level_0__i_data_latch[27]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ (.CP(CLK),
	.D(N29),
	.Q(wire_tree_level_0__i_data_latch[26]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ (.CP(CLK),
	.D(N28),
	.Q(wire_tree_level_0__i_data_latch[25]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ (.CP(CLK),
	.D(N27),
	.Q(wire_tree_level_0__i_data_latch[24]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ (.CP(CLK),
	.D(N26),
	.Q(wire_tree_level_0__i_data_latch[23]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ (.CP(CLK),
	.D(N25),
	.Q(wire_tree_level_0__i_data_latch[22]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ (.CP(CLK),
	.D(N24),
	.Q(wire_tree_level_0__i_data_latch[21]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ (.CP(CLK),
	.D(N23),
	.Q(wire_tree_level_0__i_data_latch[20]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ (.CP(CLK),
	.D(N22),
	.Q(wire_tree_level_0__i_data_latch[19]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ (.CP(CLK),
	.D(N21),
	.Q(wire_tree_level_0__i_data_latch[18]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ (.CP(CLK),
	.D(N20),
	.Q(wire_tree_level_0__i_data_latch[17]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ (.CP(CLK),
	.D(N19),
	.Q(wire_tree_level_0__i_data_latch[16]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ (.CP(CLK),
	.D(N18),
	.Q(wire_tree_level_0__i_data_latch[15]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ (.CP(CLK),
	.D(N17),
	.Q(wire_tree_level_0__i_data_latch[14]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ (.CP(CLK),
	.D(N16),
	.Q(wire_tree_level_0__i_data_latch[13]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ (.CP(CLK),
	.D(N15),
	.Q(wire_tree_level_0__i_data_latch[12]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ (.CP(CLK),
	.D(N14),
	.Q(wire_tree_level_0__i_data_latch[11]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ (.CP(CLK),
	.D(N13),
	.Q(wire_tree_level_0__i_data_latch[10]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ (.CP(CLK),
	.D(N12),
	.Q(wire_tree_level_0__i_data_latch[9]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ (.CP(CLK),
	.D(N11),
	.Q(wire_tree_level_0__i_data_latch[8]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ (.CP(CLK),
	.D(N10),
	.Q(wire_tree_level_0__i_data_latch[7]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ (.CP(CLK),
	.D(N9),
	.Q(wire_tree_level_0__i_data_latch[6]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ (.CP(CLK),
	.D(N8),
	.Q(wire_tree_level_0__i_data_latch[5]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ (.CP(CLK),
	.D(N7),
	.Q(wire_tree_level_0__i_data_latch[4]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ (.CP(CLK),
	.D(N6),
	.Q(wire_tree_level_0__i_data_latch[3]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ (.CP(CLK),
	.D(N5),
	.Q(wire_tree_level_0__i_data_latch[2]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ (.CP(CLK),
	.D(N4),
	.Q(wire_tree_level_0__i_data_latch[1]));
   DFQD4BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ (.CP(CLK),
	.D(N3),
	.Q(wire_tree_level_0__i_data_latch[0]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ (.CP(CLK_clone1),
	.D(N99),
	.Q(wire_tree_level_1__i_data_latch[63]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ (.CP(CLK_clone1),
	.D(N98),
	.Q(wire_tree_level_1__i_data_latch[62]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ (.CP(CLK_clone2),
	.D(N97),
	.Q(wire_tree_level_1__i_data_latch[61]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ (.CP(CLK_clone40),
	.D(N96),
	.Q(wire_tree_level_1__i_data_latch[60]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ (.CP(CLK_clone12),
	.D(N95),
	.Q(wire_tree_level_1__i_data_latch[59]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ (.CP(CLK_clone3),
	.D(N94),
	.Q(wire_tree_level_1__i_data_latch[58]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ (.CP(CLK_clone12),
	.D(N93),
	.Q(wire_tree_level_1__i_data_latch[57]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ (.CP(CLK_clone3),
	.D(N92),
	.Q(wire_tree_level_1__i_data_latch[56]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ (.CP(CLK_clone15),
	.D(N91),
	.Q(wire_tree_level_1__i_data_latch[55]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ (.CP(CLK_clone3),
	.D(N90),
	.Q(wire_tree_level_1__i_data_latch[54]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ (.CP(CLK_clone11),
	.D(N89),
	.Q(wire_tree_level_1__i_data_latch[53]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ (.CP(CLK_clone15),
	.D(N88),
	.Q(wire_tree_level_1__i_data_latch[52]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ (.CP(CLK_clone3),
	.D(N87),
	.Q(wire_tree_level_1__i_data_latch[51]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ (.CP(CLK_clone12),
	.D(N86),
	.Q(wire_tree_level_1__i_data_latch[50]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ (.CP(CLK_clone13),
	.D(N85),
	.Q(wire_tree_level_1__i_data_latch[49]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ (.CP(CLK_clone40),
	.D(N84),
	.Q(wire_tree_level_1__i_data_latch[48]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ (.CP(CLK_clone9),
	.D(N83),
	.Q(wire_tree_level_1__i_data_latch[47]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ (.CP(CLK_clone36),
	.D(N82),
	.Q(wire_tree_level_1__i_data_latch[46]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ (.CP(CLK_clone1),
	.D(N81),
	.Q(wire_tree_level_1__i_data_latch[45]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ (.CP(CLK_clone2),
	.D(N80),
	.Q(wire_tree_level_1__i_data_latch[44]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ (.CP(CLK_clone1),
	.D(N79),
	.Q(wire_tree_level_1__i_data_latch[43]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ (.CP(CLK_clone5),
	.D(N78),
	.Q(wire_tree_level_1__i_data_latch[42]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ (.CP(CLK_clone1),
	.D(N77),
	.Q(wire_tree_level_1__i_data_latch[41]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ (.CP(CLK_clone10),
	.D(N76),
	.Q(wire_tree_level_1__i_data_latch[40]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ (.CP(CLK_clone5),
	.D(N75),
	.Q(wire_tree_level_1__i_data_latch[39]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ (.CP(CLK_clone32),
	.D(N74),
	.Q(wire_tree_level_1__i_data_latch[38]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ (.CP(CLK_clone30),
	.D(N73),
	.Q(wire_tree_level_1__i_data_latch[37]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ (.CP(CLK_clone31),
	.D(N72),
	.Q(wire_tree_level_1__i_data_latch[36]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ (.CP(CLK_clone30),
	.D(N71),
	.Q(wire_tree_level_1__i_data_latch[35]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ (.CP(CLK_clone5),
	.D(N70),
	.Q(wire_tree_level_1__i_data_latch[34]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ (.CP(CLK_clone34),
	.D(N69),
	.Q(wire_tree_level_1__i_data_latch[33]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ (.CP(CLK_clone33),
	.D(N68),
	.Q(wire_tree_level_1__i_data_latch[32]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ (.CP(CLK_clone1),
	.D(N99),
	.Q(wire_tree_level_1__i_data_latch[31]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ (.CP(CLK_clone1),
	.D(N98),
	.Q(wire_tree_level_1__i_data_latch[30]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ (.CP(CLK_clone2),
	.D(N97),
	.Q(wire_tree_level_1__i_data_latch[29]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ (.CP(CLK_clone36),
	.D(N96),
	.Q(wire_tree_level_1__i_data_latch[28]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ (.CP(CLK_clone12),
	.D(N95),
	.Q(wire_tree_level_1__i_data_latch[27]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ (.CP(CLK_clone3),
	.D(N94),
	.Q(wire_tree_level_1__i_data_latch[26]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ (.CP(CLK_clone12),
	.D(N93),
	.Q(wire_tree_level_1__i_data_latch[25]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ (.CP(CLK_clone3),
	.D(N92),
	.Q(wire_tree_level_1__i_data_latch[24]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ (.CP(CLK_clone3),
	.D(N91),
	.Q(wire_tree_level_1__i_data_latch[23]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ (.CP(CLK_clone3),
	.D(N90),
	.Q(wire_tree_level_1__i_data_latch[22]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ (.CP(CLK_clone11),
	.D(N89),
	.Q(wire_tree_level_1__i_data_latch[21]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ (.CP(CLK_clone3),
	.D(N88),
	.Q(wire_tree_level_1__i_data_latch[20]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ (.CP(CLK_clone3),
	.D(N87),
	.Q(wire_tree_level_1__i_data_latch[19]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ (.CP(CLK_clone12),
	.D(N86),
	.Q(wire_tree_level_1__i_data_latch[18]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ (.CP(CLK_clone9),
	.D(N85),
	.Q(wire_tree_level_1__i_data_latch[17]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ (.CP(CLK_clone13),
	.D(N84),
	.Q(wire_tree_level_1__i_data_latch[16]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ (.CP(CLK_clone9),
	.D(N83),
	.Q(wire_tree_level_1__i_data_latch[15]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ (.CP(CLK_clone9),
	.D(N82),
	.Q(wire_tree_level_1__i_data_latch[14]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ (.CP(CLK_clone1),
	.D(N81),
	.Q(wire_tree_level_1__i_data_latch[13]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ (.CP(CLK_clone2),
	.D(N80),
	.Q(wire_tree_level_1__i_data_latch[12]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ (.CP(CLK_clone1),
	.D(N79),
	.Q(wire_tree_level_1__i_data_latch[11]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ (.CP(CLK_clone5),
	.D(N78),
	.Q(wire_tree_level_1__i_data_latch[10]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ (.CP(CLK_clone10),
	.D(N77),
	.Q(wire_tree_level_1__i_data_latch[9]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ (.CP(CLK_clone10),
	.D(N76),
	.Q(wire_tree_level_1__i_data_latch[8]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ (.CP(CLK_clone5),
	.D(N75),
	.Q(wire_tree_level_1__i_data_latch[7]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ (.CP(CLK_clone6),
	.D(N74),
	.Q(wire_tree_level_1__i_data_latch[6]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ (.CP(CLK_clone32),
	.D(N73),
	.Q(wire_tree_level_1__i_data_latch[5]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ (.CP(CLK_clone32),
	.D(N72),
	.Q(wire_tree_level_1__i_data_latch[4]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ (.CP(CLK_clone32),
	.D(N71),
	.Q(wire_tree_level_1__i_data_latch[3]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ (.CP(CLK_clone5),
	.D(N70),
	.Q(wire_tree_level_1__i_data_latch[2]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ (.CP(CLK_clone34),
	.D(N69),
	.Q(wire_tree_level_1__i_data_latch[1]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ (.CP(CLK_clone35),
	.D(N68),
	.Q(wire_tree_level_1__i_data_latch[0]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ (.CP(CLK_clone44),
	.D(N101),
	.Q(wire_tree_level_1__i_valid_latch[1]));
   DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ (.CP(CLK_clone44),
	.D(N101),
	.Q(wire_tree_level_1__i_valid_latch[0]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ (.CP(CLK_clone10),
	.D(N165),
	.Q(wire_tree_level_2__i_data_latch[63]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ (.CP(CLK_clone10),
	.D(N164),
	.Q(wire_tree_level_2__i_data_latch[62]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ (.CP(CLK_clone2),
	.D(N163),
	.Q(wire_tree_level_2__i_data_latch[61]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ (.CP(CLK_clone36),
	.D(N162),
	.Q(wire_tree_level_2__i_data_latch[60]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ (.CP(CLK_clone12),
	.D(N161),
	.Q(wire_tree_level_2__i_data_latch[59]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ (.CP(CLK_clone3),
	.D(N160),
	.Q(wire_tree_level_2__i_data_latch[58]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ (.CP(CLK_clone12),
	.D(N159),
	.Q(wire_tree_level_2__i_data_latch[57]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ (.CP(CLK_clone3),
	.D(N158),
	.Q(wire_tree_level_2__i_data_latch[56]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ (.CP(CLK_clone16),
	.D(N157),
	.Q(wire_tree_level_2__i_data_latch[55]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ (.CP(CLK_clone3),
	.D(N156),
	.Q(wire_tree_level_2__i_data_latch[54]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ (.CP(CLK_clone13),
	.D(N155),
	.Q(wire_tree_level_2__i_data_latch[53]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ (.CP(CLK_clone3),
	.D(N154),
	.Q(wire_tree_level_2__i_data_latch[52]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ (.CP(CLK_clone3),
	.D(N153),
	.Q(wire_tree_level_2__i_data_latch[51]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ (.CP(CLK_clone2),
	.D(N152),
	.Q(wire_tree_level_2__i_data_latch[50]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ (.CP(CLK_clone36),
	.D(N151),
	.Q(wire_tree_level_2__i_data_latch[49]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ (.CP(CLK_clone13),
	.D(N150),
	.Q(wire_tree_level_2__i_data_latch[48]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ (.CP(CLK_clone35),
	.D(N149),
	.Q(wire_tree_level_2__i_data_latch[47]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ (.CP(CLK_clone35),
	.D(N148),
	.Q(wire_tree_level_2__i_data_latch[46]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ (.CP(CLK_clone1),
	.D(N147),
	.Q(wire_tree_level_2__i_data_latch[45]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ (.CP(CLK_clone2),
	.D(N146),
	.Q(wire_tree_level_2__i_data_latch[44]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ (.CP(CLK_clone10),
	.D(N145),
	.Q(wire_tree_level_2__i_data_latch[43]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ (.CP(CLK_clone5),
	.D(N144),
	.Q(wire_tree_level_2__i_data_latch[42]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ (.CP(CLK_clone5),
	.D(N143),
	.Q(wire_tree_level_2__i_data_latch[41]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ (.CP(CLK_clone10),
	.D(N142),
	.Q(wire_tree_level_2__i_data_latch[40]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ (.CP(CLK_clone5),
	.D(N141),
	.Q(wire_tree_level_2__i_data_latch[39]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ (.CP(CLK_clone32),
	.D(N140),
	.Q(wire_tree_level_2__i_data_latch[38]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ (.CP(CLK_clone32),
	.D(N139),
	.Q(wire_tree_level_2__i_data_latch[37]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ (.CP(CLK_clone31),
	.D(N138),
	.Q(wire_tree_level_2__i_data_latch[36]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ (.CP(CLK_clone32),
	.D(N137),
	.Q(wire_tree_level_2__i_data_latch[35]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ (.CP(CLK_clone5),
	.D(N136),
	.Q(wire_tree_level_2__i_data_latch[34]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ (.CP(CLK_clone32),
	.D(N135),
	.Q(wire_tree_level_2__i_data_latch[33]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ (.CP(CLK_clone35),
	.D(N134),
	.Q(wire_tree_level_2__i_data_latch[32]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ (.CP(CLK_clone10),
	.D(N165),
	.Q(wire_tree_level_2__i_data_latch[31]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ (.CP(CLK_clone10),
	.D(N164),
	.Q(wire_tree_level_2__i_data_latch[30]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ (.CP(CLK_clone2),
	.D(N163),
	.Q(wire_tree_level_2__i_data_latch[29]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ (.CP(CLK_clone36),
	.D(N162),
	.Q(wire_tree_level_2__i_data_latch[28]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ (.CP(CLK_clone2),
	.D(N161),
	.Q(wire_tree_level_2__i_data_latch[27]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ (.CP(CLK_clone3),
	.D(N160),
	.Q(wire_tree_level_2__i_data_latch[26]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ (.CP(CLK_clone12),
	.D(N159),
	.Q(wire_tree_level_2__i_data_latch[25]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ (.CP(CLK_clone3),
	.D(N158),
	.Q(wire_tree_level_2__i_data_latch[24]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ (.CP(CLK_clone16),
	.D(N157),
	.Q(wire_tree_level_2__i_data_latch[23]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ (.CP(CLK_clone3),
	.D(N156),
	.Q(wire_tree_level_2__i_data_latch[22]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ (.CP(CLK_clone13),
	.D(N155),
	.Q(wire_tree_level_2__i_data_latch[21]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ (.CP(CLK_clone3),
	.D(N154),
	.Q(wire_tree_level_2__i_data_latch[20]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ (.CP(CLK_clone3),
	.D(N153),
	.Q(wire_tree_level_2__i_data_latch[19]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ (.CP(CLK_clone2),
	.D(N152),
	.Q(wire_tree_level_2__i_data_latch[18]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ (.CP(CLK_clone36),
	.D(N151),
	.Q(wire_tree_level_2__i_data_latch[17]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ (.CP(CLK_clone13),
	.D(N150),
	.Q(wire_tree_level_2__i_data_latch[16]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ (.CP(CLK_clone35),
	.D(N149),
	.Q(wire_tree_level_2__i_data_latch[15]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ (.CP(CLK_clone35),
	.D(N148),
	.Q(wire_tree_level_2__i_data_latch[14]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ (.CP(CLK_clone1),
	.D(N147),
	.Q(wire_tree_level_2__i_data_latch[13]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ (.CP(CLK_clone2),
	.D(N146),
	.Q(wire_tree_level_2__i_data_latch[12]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ (.CP(CLK_clone10),
	.D(N145),
	.Q(wire_tree_level_2__i_data_latch[11]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ (.CP(CLK_clone5),
	.D(N144),
	.Q(wire_tree_level_2__i_data_latch[10]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ (.CP(CLK_clone5),
	.D(N143),
	.Q(wire_tree_level_2__i_data_latch[9]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ (.CP(CLK_clone10),
	.D(N142),
	.Q(wire_tree_level_2__i_data_latch[8]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ (.CP(CLK_clone5),
	.D(N141),
	.Q(wire_tree_level_2__i_data_latch[7]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ (.CP(CLK_clone32),
	.D(N140),
	.Q(wire_tree_level_2__i_data_latch[6]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ (.CP(CLK_clone32),
	.D(N139),
	.Q(wire_tree_level_2__i_data_latch[5]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ (.CP(CLK_clone31),
	.D(N138),
	.Q(wire_tree_level_2__i_data_latch[4]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ (.CP(CLK_clone32),
	.D(N137),
	.Q(wire_tree_level_2__i_data_latch[3]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ (.CP(CLK_clone5),
	.D(N136),
	.Q(wire_tree_level_2__i_data_latch[2]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ (.CP(CLK_clone32),
	.D(N135),
	.Q(wire_tree_level_2__i_data_latch[1]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ (.CP(CLK_clone35),
	.D(N134),
	.Q(wire_tree_level_2__i_data_latch[0]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ (.CP(CLK_clone44),
	.D(N167),
	.Q(wire_tree_level_2__i_valid_latch[1]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ (.CP(CLK_clone44),
	.D(N167),
	.Q(wire_tree_level_2__i_valid_latch[0]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ (.CP(CLK_clone25),
	.D(N231),
	.Q(wire_tree_level_2__i_data_latch[127]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ (.CP(CLK_clone25),
	.D(N230),
	.Q(wire_tree_level_2__i_data_latch[126]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ (.CP(CLK_clone17),
	.D(N229),
	.Q(wire_tree_level_2__i_data_latch[125]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ (.CP(CLK_clone40),
	.D(N228),
	.Q(wire_tree_level_2__i_data_latch[124]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ (.CP(CLK_clone40),
	.D(N227),
	.Q(wire_tree_level_2__i_data_latch[123]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ (.CP(CLK_clone38),
	.D(N226),
	.Q(wire_tree_level_2__i_data_latch[122]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ (.CP(CLK_clone38),
	.D(N225),
	.Q(wire_tree_level_2__i_data_latch[121]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ (.CP(CLK_clone43),
	.D(N224),
	.Q(wire_tree_level_2__i_data_latch[120]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ (.CP(CLK_clone43),
	.D(N223),
	.Q(wire_tree_level_2__i_data_latch[119]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ (.CP(CLK_clone39),
	.D(N222),
	.Q(wire_tree_level_2__i_data_latch[118]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ (.CP(CLK_clone43),
	.D(N221),
	.Q(wire_tree_level_2__i_data_latch[117]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ (.CP(CLK_clone43),
	.D(N220),
	.Q(wire_tree_level_2__i_data_latch[116]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ (.CP(CLK_clone43),
	.D(N219),
	.Q(wire_tree_level_2__i_data_latch[115]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ (.CP(CLK_clone38),
	.D(N218),
	.Q(wire_tree_level_2__i_data_latch[114]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ (.CP(CLK_clone40),
	.D(N217),
	.Q(wire_tree_level_2__i_data_latch[113]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ (.CP(CLK_clone40),
	.D(N216),
	.Q(wire_tree_level_2__i_data_latch[112]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ (.CP(CLK_clone40),
	.D(N215),
	.Q(wire_tree_level_2__i_data_latch[111]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ (.CP(CLK_clone17),
	.D(N214),
	.Q(wire_tree_level_2__i_data_latch[110]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ (.CP(CLK_clone17),
	.D(N213),
	.Q(wire_tree_level_2__i_data_latch[109]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ (.CP(CLK_clone17),
	.D(N212),
	.Q(wire_tree_level_2__i_data_latch[108]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ (.CP(CLK_clone25),
	.D(N211),
	.Q(wire_tree_level_2__i_data_latch[107]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ (.CP(CLK_clone29),
	.D(N210),
	.Q(wire_tree_level_2__i_data_latch[106]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ (.CP(CLK_clone25),
	.D(N209),
	.Q(wire_tree_level_2__i_data_latch[105]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ (.CP(CLK_clone29),
	.D(N208),
	.Q(wire_tree_level_2__i_data_latch[104]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ (.CP(CLK_clone29),
	.D(N207),
	.Q(wire_tree_level_2__i_data_latch[103]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ (.CP(CLK_clone30),
	.D(N206),
	.Q(wire_tree_level_2__i_data_latch[102]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ (.CP(CLK_clone30),
	.D(N205),
	.Q(wire_tree_level_2__i_data_latch[101]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ (.CP(CLK_clone30),
	.D(N204),
	.Q(wire_tree_level_2__i_data_latch[100]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ (.CP(CLK_clone22),
	.D(N203),
	.Q(wire_tree_level_2__i_data_latch[99]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ (.CP(CLK_clone29),
	.D(N202),
	.Q(wire_tree_level_2__i_data_latch[98]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ (.CP(CLK_clone25),
	.D(N201),
	.Q(wire_tree_level_2__i_data_latch[97]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ (.CP(CLK_clone25),
	.D(N200),
	.Q(wire_tree_level_2__i_data_latch[96]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ (.CP(CLK_clone25),
	.D(N231),
	.Q(wire_tree_level_2__i_data_latch[95]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ (.CP(CLK_clone18),
	.D(N230),
	.Q(wire_tree_level_2__i_data_latch[94]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ (.CP(CLK_clone17),
	.D(N229),
	.Q(wire_tree_level_2__i_data_latch[93]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ (.CP(CLK_clone40),
	.D(N228),
	.Q(wire_tree_level_2__i_data_latch[92]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ (.CP(CLK_clone40),
	.D(N227),
	.Q(wire_tree_level_2__i_data_latch[91]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ (.CP(CLK_clone38),
	.D(N226),
	.Q(wire_tree_level_2__i_data_latch[90]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ (.CP(CLK_clone38),
	.D(N225),
	.Q(wire_tree_level_2__i_data_latch[89]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ (.CP(CLK_clone43),
	.D(N224),
	.Q(wire_tree_level_2__i_data_latch[88]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ (.CP(CLK_clone43),
	.D(N223),
	.Q(wire_tree_level_2__i_data_latch[87]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ (.CP(CLK_clone38),
	.D(N222),
	.Q(wire_tree_level_2__i_data_latch[86]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ (.CP(CLK_clone43),
	.D(N221),
	.Q(wire_tree_level_2__i_data_latch[85]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ (.CP(CLK_clone43),
	.D(N220),
	.Q(wire_tree_level_2__i_data_latch[84]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ (.CP(CLK_clone43),
	.D(N219),
	.Q(wire_tree_level_2__i_data_latch[83]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ (.CP(CLK_clone38),
	.D(N218),
	.Q(wire_tree_level_2__i_data_latch[82]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ (.CP(CLK_clone40),
	.D(N217),
	.Q(wire_tree_level_2__i_data_latch[81]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ (.CP(CLK_clone40),
	.D(N216),
	.Q(wire_tree_level_2__i_data_latch[80]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ (.CP(CLK_clone40),
	.D(N215),
	.Q(wire_tree_level_2__i_data_latch[79]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ (.CP(CLK_clone17),
	.D(N214),
	.Q(wire_tree_level_2__i_data_latch[78]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ (.CP(CLK_clone25),
	.D(N213),
	.Q(wire_tree_level_2__i_data_latch[77]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ (.CP(CLK_clone17),
	.D(N212),
	.Q(wire_tree_level_2__i_data_latch[76]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ (.CP(CLK_clone25),
	.D(N211),
	.Q(wire_tree_level_2__i_data_latch[75]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ (.CP(CLK_clone29),
	.D(N210),
	.Q(wire_tree_level_2__i_data_latch[74]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ (.CP(CLK_clone25),
	.D(N209),
	.Q(wire_tree_level_2__i_data_latch[73]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ (.CP(CLK_clone25),
	.D(N208),
	.Q(wire_tree_level_2__i_data_latch[72]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ (.CP(CLK_clone29),
	.D(N207),
	.Q(wire_tree_level_2__i_data_latch[71]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ (.CP(CLK_clone30),
	.D(N206),
	.Q(wire_tree_level_2__i_data_latch[70]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ (.CP(CLK_clone30),
	.D(N205),
	.Q(wire_tree_level_2__i_data_latch[69]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ (.CP(CLK_clone30),
	.D(N204),
	.Q(wire_tree_level_2__i_data_latch[68]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ (.CP(CLK_clone30),
	.D(N203),
	.Q(wire_tree_level_2__i_data_latch[67]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ (.CP(CLK_clone23),
	.D(N202),
	.Q(wire_tree_level_2__i_data_latch[66]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ (.CP(CLK_clone25),
	.D(N201),
	.Q(wire_tree_level_2__i_data_latch[65]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ (.CP(CLK_clone18),
	.D(N200),
	.Q(wire_tree_level_2__i_data_latch[64]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ (.CP(CLK_clone44),
	.D(N233),
	.Q(wire_tree_level_2__i_valid_latch[3]));
   DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ (.CP(CLK_clone41),
	.D(N233),
	.Q(wire_tree_level_2__i_valid_latch[2]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ (.CP(CLK_clone10),
	.D(N297),
	.Q(o_data_bus[63]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ (.CP(CLK_clone10),
	.D(N296),
	.Q(o_data_bus[62]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ (.CP(CLK_clone2),
	.D(N295),
	.Q(o_data_bus[61]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ (.CP(CLK_clone36),
	.D(N294),
	.Q(o_data_bus[60]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ (.CP(CLK_clone2),
	.D(N293),
	.Q(o_data_bus[59]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ (.CP(CLK_clone15),
	.D(N292),
	.Q(o_data_bus[58]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ (.CP(CLK_clone12),
	.D(N291),
	.Q(o_data_bus[57]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ (.CP(CLK_clone3),
	.D(N290),
	.Q(o_data_bus[56]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ (.CP(CLK_clone16),
	.D(N289),
	.Q(o_data_bus[55]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ (.CP(CLK_clone3),
	.D(N288),
	.Q(o_data_bus[54]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ (.CP(CLK_clone13),
	.D(N287),
	.Q(o_data_bus[53]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ (.CP(CLK_clone3),
	.D(N286),
	.Q(o_data_bus[52]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ (.CP(CLK_clone3),
	.D(N285),
	.Q(o_data_bus[51]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ (.CP(CLK_clone2),
	.D(N284),
	.Q(o_data_bus[50]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ (.CP(CLK_clone35),
	.D(N283),
	.Q(o_data_bus[49]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ (.CP(CLK_clone36),
	.D(N282),
	.Q(o_data_bus[48]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ (.CP(CLK_clone35),
	.D(N281),
	.Q(o_data_bus[47]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ (.CP(CLK_clone35),
	.D(N280),
	.Q(o_data_bus[46]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ (.CP(CLK_clone10),
	.D(N279),
	.Q(o_data_bus[45]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ (.CP(CLK_clone2),
	.D(N278),
	.Q(o_data_bus[44]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ (.CP(CLK_clone10),
	.D(N277),
	.Q(o_data_bus[43]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ (.CP(CLK_clone4),
	.D(N276),
	.Q(o_data_bus[42]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ (.CP(CLK_clone5),
	.D(N275),
	.Q(o_data_bus[41]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ (.CP(CLK_clone5),
	.D(N274),
	.Q(o_data_bus[40]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ (.CP(CLK_clone5),
	.D(N273),
	.Q(o_data_bus[39]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ (.CP(CLK_clone32),
	.D(N272),
	.Q(o_data_bus[38]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ (.CP(CLK_clone32),
	.D(N271),
	.Q(o_data_bus[37]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ (.CP(CLK_clone31),
	.D(N270),
	.Q(o_data_bus[36]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ (.CP(CLK_clone28),
	.D(N269),
	.Q(o_data_bus[35]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ (.CP(CLK_clone4),
	.D(N268),
	.Q(o_data_bus[34]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ (.CP(CLK_clone32),
	.D(N267),
	.Q(o_data_bus[33]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ (.CP(CLK_clone35),
	.D(N266),
	.Q(o_data_bus[32]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ (.CP(CLK_clone10),
	.D(N297),
	.Q(o_data_bus[31]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ (.CP(CLK_clone10),
	.D(N296),
	.Q(o_data_bus[30]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ (.CP(CLK_clone2),
	.D(N295),
	.Q(o_data_bus[29]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ (.CP(CLK_clone36),
	.D(N294),
	.Q(o_data_bus[28]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ (.CP(CLK_clone2),
	.D(N293),
	.Q(o_data_bus[27]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ (.CP(CLK_clone15),
	.D(N292),
	.Q(o_data_bus[26]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ (.CP(CLK_clone12),
	.D(N291),
	.Q(o_data_bus[25]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ (.CP(CLK_clone3),
	.D(N290),
	.Q(o_data_bus[24]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ (.CP(CLK_clone16),
	.D(N289),
	.Q(o_data_bus[23]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ (.CP(CLK_clone3),
	.D(N288),
	.Q(o_data_bus[22]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ (.CP(CLK_clone13),
	.D(N287),
	.Q(o_data_bus[21]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ (.CP(CLK_clone3),
	.D(N286),
	.Q(o_data_bus[20]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ (.CP(CLK_clone3),
	.D(N285),
	.Q(o_data_bus[19]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ (.CP(CLK_clone2),
	.D(N284),
	.Q(o_data_bus[18]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ (.CP(CLK_clone36),
	.D(N283),
	.Q(o_data_bus[17]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ (.CP(CLK_clone13),
	.D(N282),
	.Q(o_data_bus[16]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ (.CP(CLK_clone35),
	.D(N281),
	.Q(o_data_bus[15]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ (.CP(CLK_clone35),
	.D(N280),
	.Q(o_data_bus[14]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ (.CP(CLK_clone10),
	.D(N279),
	.Q(o_data_bus[13]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ (.CP(CLK_clone2),
	.D(N278),
	.Q(o_data_bus[12]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ (.CP(CLK_clone10),
	.D(N277),
	.Q(o_data_bus[11]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ (.CP(CLK_clone5),
	.D(N276),
	.Q(o_data_bus[10]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ (.CP(CLK_clone5),
	.D(N275),
	.Q(o_data_bus[9]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ (.CP(CLK_clone5),
	.D(N274),
	.Q(o_data_bus[8]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ (.CP(CLK_clone5),
	.D(N273),
	.Q(o_data_bus[7]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ (.CP(CLK_clone32),
	.D(N272),
	.Q(o_data_bus[6]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ (.CP(CLK_clone32),
	.D(N271),
	.Q(o_data_bus[5]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ (.CP(CLK_clone31),
	.D(N270),
	.Q(o_data_bus[4]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ (.CP(CLK_clone32),
	.D(N269),
	.Q(o_data_bus[3]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ (.CP(CLK_clone6),
	.D(N268),
	.Q(o_data_bus[2]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ (.CP(CLK_clone32),
	.D(N267),
	.Q(o_data_bus[1]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ (.CP(CLK_clone35),
	.D(N266),
	.Q(o_data_bus[0]));
   DFQD1BWP30P140LVT o_valid_reg_reg_1_ (.CP(CLK_clone14),
	.D(N299),
	.Q(o_valid[1]));
   DFQD1BWP30P140LVT o_valid_reg_reg_0_ (.CP(CLK_clone11),
	.D(N299),
	.Q(o_valid[0]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ (.CP(CLK_clone10),
	.D(N363),
	.Q(o_data_bus[127]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ (.CP(CLK_clone10),
	.D(N362),
	.Q(o_data_bus[126]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ (.CP(CLK_clone2),
	.D(N361),
	.Q(o_data_bus[125]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ (.CP(CLK_clone36),
	.D(N360),
	.Q(o_data_bus[124]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ (.CP(CLK_clone2),
	.D(N359),
	.Q(o_data_bus[123]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ (.CP(CLK_clone15),
	.D(N358),
	.Q(o_data_bus[122]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ (.CP(CLK_clone12),
	.D(N357),
	.Q(o_data_bus[121]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ (.CP(CLK_clone3),
	.D(N356),
	.Q(o_data_bus[120]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ (.CP(CLK_clone16),
	.D(N355),
	.Q(o_data_bus[119]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ (.CP(CLK_clone16),
	.D(N354),
	.Q(o_data_bus[118]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ (.CP(CLK_clone13),
	.D(N353),
	.Q(o_data_bus[117]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ (.CP(CLK_clone12),
	.D(N352),
	.Q(o_data_bus[116]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ (.CP(CLK_clone12),
	.D(N351),
	.Q(o_data_bus[115]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ (.CP(CLK_clone2),
	.D(N350),
	.Q(o_data_bus[114]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ (.CP(CLK_clone36),
	.D(N349),
	.Q(o_data_bus[113]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ (.CP(CLK_clone13),
	.D(N348),
	.Q(o_data_bus[112]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ (.CP(CLK_clone35),
	.D(N347),
	.Q(o_data_bus[111]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ (.CP(CLK_clone35),
	.D(N346),
	.Q(o_data_bus[110]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ (.CP(CLK_clone2),
	.D(N345),
	.Q(o_data_bus[109]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ (.CP(CLK_clone2),
	.D(N344),
	.Q(o_data_bus[108]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ (.CP(CLK_clone10),
	.D(N343),
	.Q(o_data_bus[107]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ (.CP(CLK_clone5),
	.D(N342),
	.Q(o_data_bus[106]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ (.CP(CLK_clone5),
	.D(N341),
	.Q(o_data_bus[105]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ (.CP(CLK_clone10),
	.D(N340),
	.Q(o_data_bus[104]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ (.CP(CLK_clone5),
	.D(N339),
	.Q(o_data_bus[103]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ (.CP(CLK_clone32),
	.D(N338),
	.Q(o_data_bus[102]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ (.CP(CLK_clone32),
	.D(N337),
	.Q(o_data_bus[101]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ (.CP(CLK_clone31),
	.D(N336),
	.Q(o_data_bus[100]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ (.CP(CLK_clone31),
	.D(N335),
	.Q(o_data_bus[99]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ (.CP(CLK_clone6),
	.D(N334),
	.Q(o_data_bus[98]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ (.CP(CLK_clone32),
	.D(N333),
	.Q(o_data_bus[97]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ (.CP(CLK_clone31),
	.D(N332),
	.Q(o_data_bus[96]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ (.CP(CLK_clone10),
	.D(N363),
	.Q(o_data_bus[95]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ (.CP(CLK_clone10),
	.D(N362),
	.Q(o_data_bus[94]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ (.CP(CLK_clone2),
	.D(N361),
	.Q(o_data_bus[93]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ (.CP(CLK_clone36),
	.D(N360),
	.Q(o_data_bus[92]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ (.CP(CLK_clone2),
	.D(N359),
	.Q(o_data_bus[91]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ (.CP(CLK_clone15),
	.D(N358),
	.Q(o_data_bus[90]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ (.CP(CLK_clone12),
	.D(N357),
	.Q(o_data_bus[89]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ (.CP(CLK_clone3),
	.D(N356),
	.Q(o_data_bus[88]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ (.CP(CLK_clone16),
	.D(N355),
	.Q(o_data_bus[87]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ (.CP(CLK_clone15),
	.D(N354),
	.Q(o_data_bus[86]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ (.CP(CLK_clone13),
	.D(N353),
	.Q(o_data_bus[85]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ (.CP(CLK_clone12),
	.D(N352),
	.Q(o_data_bus[84]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ (.CP(CLK_clone12),
	.D(N351),
	.Q(o_data_bus[83]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ (.CP(CLK_clone2),
	.D(N350),
	.Q(o_data_bus[82]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ (.CP(CLK_clone36),
	.D(N349),
	.Q(o_data_bus[81]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ (.CP(CLK_clone13),
	.D(N348),
	.Q(o_data_bus[80]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ (.CP(CLK_clone35),
	.D(N347),
	.Q(o_data_bus[79]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ (.CP(CLK_clone35),
	.D(N346),
	.Q(o_data_bus[78]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ (.CP(CLK_clone2),
	.D(N345),
	.Q(o_data_bus[77]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ (.CP(CLK_clone2),
	.D(N344),
	.Q(o_data_bus[76]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ (.CP(CLK_clone10),
	.D(N343),
	.Q(o_data_bus[75]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ (.CP(CLK_clone5),
	.D(N342),
	.Q(o_data_bus[74]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ (.CP(CLK_clone5),
	.D(N341),
	.Q(o_data_bus[73]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ (.CP(CLK_clone10),
	.D(N340),
	.Q(o_data_bus[72]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ (.CP(CLK_clone5),
	.D(N339),
	.Q(o_data_bus[71]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ (.CP(CLK_clone32),
	.D(N338),
	.Q(o_data_bus[70]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ (.CP(CLK_clone32),
	.D(N337),
	.Q(o_data_bus[69]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ (.CP(CLK_clone31),
	.D(N336),
	.Q(o_data_bus[68]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ (.CP(CLK_clone31),
	.D(N335),
	.Q(o_data_bus[67]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ (.CP(CLK_clone6),
	.D(N334),
	.Q(o_data_bus[66]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ (.CP(CLK_clone32),
	.D(N333),
	.Q(o_data_bus[65]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ (.CP(CLK_clone31),
	.D(N332),
	.Q(o_data_bus[64]));
   DFQD1BWP30P140LVT o_valid_reg_reg_3_ (.CP(CLK_clone11),
	.D(N365),
	.Q(o_valid[3]));
   DFQD1BWP30P140LVT o_valid_reg_reg_2_ (.CP(CLK_clone11),
	.D(N365),
	.Q(o_valid[2]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ (.CP(CLK_clone24),
	.D(N429),
	.Q(o_data_bus[191]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ (.CP(CLK_clone26),
	.D(N428),
	.Q(o_data_bus[190]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ (.CP(CLK_clone21),
	.D(N427),
	.Q(o_data_bus[189]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ (.CP(CLK_clone19),
	.D(N426),
	.Q(o_data_bus[188]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ (.CP(CLK_clone37),
	.D(N425),
	.Q(o_data_bus[187]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ (.CP(CLK_clone37),
	.D(N424),
	.Q(o_data_bus[186]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ (.CP(CLK_clone20),
	.D(N423),
	.Q(o_data_bus[185]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ (.CP(CLK_clone20),
	.D(N422),
	.Q(o_data_bus[184]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ (.CP(CLK_clone42),
	.D(N421),
	.Q(o_data_bus[183]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ (.CP(CLK_clone42),
	.D(N420),
	.Q(o_data_bus[182]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ (.CP(CLK_clone42),
	.D(N419),
	.Q(o_data_bus[181]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ (.CP(CLK_clone20),
	.D(N418),
	.Q(o_data_bus[180]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ (.CP(CLK_clone7),
	.D(N417),
	.Q(o_data_bus[179]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ (.CP(CLK_clone20),
	.D(N416),
	.Q(o_data_bus[178]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ (.CP(CLK_clone21),
	.D(N415),
	.Q(o_data_bus[177]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ (.CP(CLK_clone21),
	.D(N414),
	.Q(o_data_bus[176]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ (.CP(CLK_clone21),
	.D(N413),
	.Q(o_data_bus[175]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ (.CP(CLK_clone21),
	.D(N412),
	.Q(o_data_bus[174]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ (.CP(CLK_clone8),
	.D(N411),
	.Q(o_data_bus[173]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ (.CP(CLK_clone21),
	.D(N410),
	.Q(o_data_bus[172]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ (.CP(CLK_clone8),
	.D(N409),
	.Q(o_data_bus[171]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ (.CP(CLK_clone26),
	.D(N408),
	.Q(o_data_bus[170]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ (.CP(CLK_clone26),
	.D(N407),
	.Q(o_data_bus[169]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ (.CP(CLK_clone26),
	.D(N406),
	.Q(o_data_bus[168]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ (.CP(CLK_clone26),
	.D(N405),
	.Q(o_data_bus[167]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ (.CP(CLK_clone27),
	.D(N404),
	.Q(o_data_bus[166]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ (.CP(CLK_clone26),
	.D(N403),
	.Q(o_data_bus[165]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ (.CP(CLK_clone26),
	.D(N402),
	.Q(o_data_bus[164]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ (.CP(CLK_clone27),
	.D(N401),
	.Q(o_data_bus[163]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ (.CP(CLK_clone26),
	.D(N400),
	.Q(o_data_bus[162]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ (.CP(CLK_clone26),
	.D(N399),
	.Q(o_data_bus[161]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ (.CP(CLK_clone26),
	.D(N398),
	.Q(o_data_bus[160]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ (.CP(CLK_clone24),
	.D(N429),
	.Q(o_data_bus[159]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ (.CP(CLK_clone26),
	.D(N428),
	.Q(o_data_bus[158]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ (.CP(CLK_clone21),
	.D(N427),
	.Q(o_data_bus[157]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ (.CP(CLK_clone21),
	.D(N426),
	.Q(o_data_bus[156]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ (.CP(CLK_clone20),
	.D(N425),
	.Q(o_data_bus[155]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ (.CP(CLK_clone37),
	.D(N424),
	.Q(o_data_bus[154]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ (.CP(CLK_clone20),
	.D(N423),
	.Q(o_data_bus[153]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ (.CP(CLK_clone42),
	.D(N422),
	.Q(o_data_bus[152]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ (.CP(CLK_clone42),
	.D(N421),
	.Q(o_data_bus[151]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ (.CP(CLK_clone42),
	.D(N420),
	.Q(o_data_bus[150]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ (.CP(CLK_clone42),
	.D(N419),
	.Q(o_data_bus[149]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ (.CP(CLK_clone20),
	.D(N418),
	.Q(o_data_bus[148]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ (.CP(CLK_clone7),
	.D(N417),
	.Q(o_data_bus[147]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ (.CP(CLK_clone37),
	.D(N416),
	.Q(o_data_bus[146]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ (.CP(CLK_clone21),
	.D(N415),
	.Q(o_data_bus[145]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ (.CP(CLK_clone21),
	.D(N414),
	.Q(o_data_bus[144]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ (.CP(CLK_clone21),
	.D(N413),
	.Q(o_data_bus[143]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ (.CP(CLK_clone21),
	.D(N412),
	.Q(o_data_bus[142]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ (.CP(CLK_clone8),
	.D(N411),
	.Q(o_data_bus[141]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ (.CP(CLK_clone21),
	.D(N410),
	.Q(o_data_bus[140]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ (.CP(CLK_clone8),
	.D(N409),
	.Q(o_data_bus[139]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ (.CP(CLK_clone26),
	.D(N408),
	.Q(o_data_bus[138]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ (.CP(CLK_clone26),
	.D(N407),
	.Q(o_data_bus[137]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ (.CP(CLK_clone26),
	.D(N406),
	.Q(o_data_bus[136]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ (.CP(CLK_clone26),
	.D(N405),
	.Q(o_data_bus[135]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ (.CP(CLK_clone27),
	.D(N404),
	.Q(o_data_bus[134]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ (.CP(CLK_clone26),
	.D(N403),
	.Q(o_data_bus[133]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ (.CP(CLK_clone26),
	.D(N402),
	.Q(o_data_bus[132]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ (.CP(CLK_clone27),
	.D(N401),
	.Q(o_data_bus[131]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ (.CP(CLK_clone26),
	.D(N400),
	.Q(o_data_bus[130]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ (.CP(CLK_clone26),
	.D(N399),
	.Q(o_data_bus[129]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ (.CP(CLK_clone26),
	.D(N398),
	.Q(o_data_bus[128]));
   DFQD1BWP30P140LVT o_valid_reg_reg_5_ (.CP(CLK_clone7),
	.D(N431),
	.Q(o_valid[5]));
   DFQD1BWP30P140LVT o_valid_reg_reg_4_ (.CP(CLK_clone7),
	.D(N431),
	.Q(o_valid[4]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ (.CP(CLK_clone25),
	.D(N495),
	.Q(o_data_bus[255]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ (.CP(CLK_clone25),
	.D(N494),
	.Q(o_data_bus[254]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ (.CP(CLK_clone17),
	.D(N493),
	.Q(o_data_bus[253]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ (.CP(CLK_clone17),
	.D(N492),
	.Q(o_data_bus[252]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ (.CP(CLK_clone40),
	.D(N491),
	.Q(o_data_bus[251]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ (.CP(CLK_clone38),
	.D(N490),
	.Q(o_data_bus[250]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ (.CP(CLK_clone38),
	.D(N489),
	.Q(o_data_bus[249]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ (.CP(CLK_clone43),
	.D(N488),
	.Q(o_data_bus[248]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ (.CP(CLK_clone38),
	.D(N487),
	.Q(o_data_bus[247]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ (.CP(CLK_clone38),
	.D(N486),
	.Q(o_data_bus[246]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ (.CP(CLK_clone43),
	.D(N485),
	.Q(o_data_bus[245]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ (.CP(CLK_clone43),
	.D(N484),
	.Q(o_data_bus[244]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ (.CP(CLK_clone43),
	.D(N483),
	.Q(o_data_bus[243]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ (.CP(CLK_clone40),
	.D(N482),
	.Q(o_data_bus[242]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ (.CP(CLK_clone40),
	.D(N481),
	.Q(o_data_bus[241]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ (.CP(CLK_clone40),
	.D(N480),
	.Q(o_data_bus[240]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ (.CP(CLK_clone40),
	.D(N479),
	.Q(o_data_bus[239]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ (.CP(CLK_clone17),
	.D(N478),
	.Q(o_data_bus[238]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ (.CP(CLK_clone17),
	.D(N477),
	.Q(o_data_bus[237]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ (.CP(CLK_clone17),
	.D(N476),
	.Q(o_data_bus[236]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ (.CP(CLK_clone25),
	.D(N475),
	.Q(o_data_bus[235]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ (.CP(CLK_clone29),
	.D(N474),
	.Q(o_data_bus[234]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ (.CP(CLK_clone25),
	.D(N473),
	.Q(o_data_bus[233]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ (.CP(CLK_clone29),
	.D(N472),
	.Q(o_data_bus[232]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ (.CP(CLK_clone29),
	.D(N471),
	.Q(o_data_bus[231]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ (.CP(CLK_clone29),
	.D(N470),
	.Q(o_data_bus[230]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ (.CP(CLK_clone22),
	.D(N469),
	.Q(o_data_bus[229]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ (.CP(CLK_clone29),
	.D(N468),
	.Q(o_data_bus[228]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ (.CP(CLK_clone22),
	.D(N467),
	.Q(o_data_bus[227]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ (.CP(CLK_clone29),
	.D(N466),
	.Q(o_data_bus[226]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ (.CP(CLK_clone29),
	.D(N465),
	.Q(o_data_bus[225]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ (.CP(CLK_clone25),
	.D(N464),
	.Q(o_data_bus[224]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ (.CP(CLK_clone25),
	.D(N495),
	.Q(o_data_bus[223]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ (.CP(CLK_clone25),
	.D(N494),
	.Q(o_data_bus[222]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ (.CP(CLK_clone17),
	.D(N493),
	.Q(o_data_bus[221]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ (.CP(CLK_clone17),
	.D(N492),
	.Q(o_data_bus[220]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ (.CP(CLK_clone40),
	.D(N491),
	.Q(o_data_bus[219]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ (.CP(CLK_clone38),
	.D(N490),
	.Q(o_data_bus[218]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ (.CP(CLK_clone38),
	.D(N489),
	.Q(o_data_bus[217]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ (.CP(CLK_clone43),
	.D(N488),
	.Q(o_data_bus[216]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ (.CP(CLK_clone38),
	.D(N487),
	.Q(o_data_bus[215]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ (.CP(CLK_clone38),
	.D(N486),
	.Q(o_data_bus[214]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ (.CP(CLK_clone43),
	.D(N485),
	.Q(o_data_bus[213]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ (.CP(CLK_clone43),
	.D(N484),
	.Q(o_data_bus[212]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ (.CP(CLK_clone43),
	.D(N483),
	.Q(o_data_bus[211]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ (.CP(CLK_clone38),
	.D(N482),
	.Q(o_data_bus[210]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ (.CP(CLK_clone40),
	.D(N481),
	.Q(o_data_bus[209]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ (.CP(CLK_clone40),
	.D(N480),
	.Q(o_data_bus[208]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ (.CP(CLK_clone40),
	.D(N479),
	.Q(o_data_bus[207]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ (.CP(CLK_clone17),
	.D(N478),
	.Q(o_data_bus[206]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ (.CP(CLK_clone17),
	.D(N477),
	.Q(o_data_bus[205]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ (.CP(CLK_clone17),
	.D(N476),
	.Q(o_data_bus[204]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ (.CP(CLK_clone25),
	.D(N475),
	.Q(o_data_bus[203]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ (.CP(CLK_clone29),
	.D(N474),
	.Q(o_data_bus[202]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ (.CP(CLK_clone25),
	.D(N473),
	.Q(o_data_bus[201]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ (.CP(CLK_clone29),
	.D(N472),
	.Q(o_data_bus[200]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ (.CP(CLK_clone29),
	.D(N471),
	.Q(o_data_bus[199]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ (.CP(CLK_clone29),
	.D(N470),
	.Q(o_data_bus[198]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ (.CP(CLK_clone30),
	.D(N469),
	.Q(o_data_bus[197]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ (.CP(CLK_clone29),
	.D(N468),
	.Q(o_data_bus[196]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ (.CP(CLK_clone30),
	.D(N467),
	.Q(o_data_bus[195]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ (.CP(CLK_clone29),
	.D(N466),
	.Q(o_data_bus[194]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ (.CP(CLK_clone29),
	.D(N465),
	.Q(o_data_bus[193]));
   DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ (.CP(CLK_clone25),
	.D(N464),
	.Q(o_data_bus[192]));
   DFQD1BWP30P140LVT o_valid_reg_reg_7_ (.CP(CLK_clone41),
	.D(N497),
	.Q(o_valid[7]));
   DFQD1BWP30P140LVT o_valid_reg_reg_6_ (.CP(CLK_clone41),
	.D(N497),
	.Q(o_valid[6]));
   INR2D4BWP30P140LVT U3 (.A1(i_en),
	.B1(rst),
	.ZN(n1));
   AN2D4BWP30P140LVT U5 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.A2(i_data_bus[31]),
	.Z(N34));
   AN2D4BWP30P140LVT U6 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.A2(i_data_bus[0]),
	.Z(N3));
   AN2D4BWP30P140LVT U7 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.A2(i_data_bus[1]),
	.Z(N4));
   CKAN2D1BWP30P140LVT U8 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.A2(i_data_bus[2]),
	.Z(N5));
   AN2D4BWP30P140LVT U9 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.A2(i_data_bus[3]),
	.Z(N6));
   CKAN2D1BWP30P140LVT U10 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.A2(i_data_bus[4]),
	.Z(N7));
   AN2D4BWP30P140LVT U11 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.A2(i_data_bus[5]),
	.Z(N8));
   CKAN2D1BWP30P140LVT U12 (.A1(FE_OCPN1375_FE_OFN344_n1),
	.A2(i_data_bus[6]),
	.Z(N9));
   CKAN2D1BWP30P140LVT U13 (.A1(FE_OCPN1375_FE_OFN344_n1),
	.A2(i_data_bus[7]),
	.Z(N10));
   AN2D4BWP30P140LVT U14 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.A2(i_data_bus[8]),
	.Z(N11));
   AN2D4BWP30P140LVT U15 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.A2(i_data_bus[9]),
	.Z(N12));
   AN2D4BWP30P140LVT U16 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.A2(i_data_bus[10]),
	.Z(N13));
   AN2D4BWP30P140LVT U17 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.A2(i_data_bus[11]),
	.Z(N14));
   AN2D4BWP30P140LVT U18 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.A2(i_data_bus[12]),
	.Z(N15));
   AN2D4BWP30P140LVT U22 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.A2(i_data_bus[16]),
	.Z(N19));
   CKAN2D1BWP30P140LVT U23 (.A1(FE_OCPN1375_FE_OFN344_n1),
	.A2(i_data_bus[17]),
	.Z(N20));
   AN2D4BWP30P140LVT U24 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.A2(i_data_bus[18]),
	.Z(N21));
   AN2D4BWP30P140LVT U25 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.A2(i_data_bus[19]),
	.Z(N22));
   AN2D4BWP30P140LVT U26 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.A2(i_data_bus[20]),
	.Z(N23));
   AN2D4BWP30P140LVT U27 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.A2(i_data_bus[21]),
	.Z(N24));
   AN2D4BWP30P140LVT U29 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.A2(i_data_bus[23]),
	.Z(N26));
   AN2D4BWP30P140LVT U30 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.A2(i_data_bus[24]),
	.Z(N27));
   AN2D4BWP30P140LVT U31 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.A2(i_data_bus[25]),
	.Z(N28));
   CKAN2D1BWP30P140LVT U32 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.A2(i_data_bus[26]),
	.Z(N29));
   AN2D4BWP30P140LVT U34 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.A2(i_data_bus[28]),
	.Z(N31));
   AN2D4BWP30P140LVT U35 (.A1(FE_OCPN1376_FE_OFN344_n1),
	.A2(i_data_bus[29]),
	.Z(N32));
   CKAN2D1BWP30P140LVT U37 (.A1(FE_OCPN1467_n1),
	.A2(wire_tree_level_0__i_data_latch[31]),
	.Z(N99));
   CKAN2D1BWP30P140LVT U38 (.A1(FE_OCPN1467_n1),
	.A2(wire_tree_level_0__i_data_latch[30]),
	.Z(N98));
   CKAN2D1BWP30P140LVT U39 (.A1(FE_OCPN1466_n1),
	.A2(wire_tree_level_0__i_data_latch[23]),
	.Z(N91));
   CKAN2D0BWP30P140LVT U40 (.A1(FE_OCPN1375_FE_OFN344_n1),
	.A2(wire_tree_level_0__i_data_latch[22]),
	.Z(N90));
   CKAN2D1BWP30P140LVT U41 (.A1(FE_OCPN1469_n1),
	.A2(wire_tree_level_0__i_data_latch[21]),
	.Z(N89));
   CKAN2D1BWP30P140LVT U42 (.A1(FE_OCPN1375_FE_OFN344_n1),
	.A2(wire_tree_level_0__i_data_latch[20]),
	.Z(N88));
   CKAN2D1BWP30P140LVT U43 (.A1(FE_OCPN1375_FE_OFN344_n1),
	.A2(wire_tree_level_0__i_data_latch[19]),
	.Z(N87));
   CKAN2D1BWP30P140LVT U44 (.A1(FE_OCPN1375_FE_OFN344_n1),
	.A2(wire_tree_level_0__i_data_latch[18]),
	.Z(N86));
   CKAN2D1BWP30P140LVT U45 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_0__i_data_latch[17]),
	.Z(N85));
   CKAN2D1BWP30P140LVT U46 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_0__i_data_latch[16]),
	.Z(N84));
   CKAN2D0BWP30P140LVT U47 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_0__i_data_latch[15]),
	.Z(N83));
   CKAN2D1BWP30P140LVT U48 (.A1(FE_OCPN1374_FE_OFN752_n1),
	.A2(wire_tree_level_0__i_data_latch[14]),
	.Z(N82));
   CKAN2D1BWP30P140LVT U49 (.A1(FE_OCPN1467_n1),
	.A2(wire_tree_level_0__i_data_latch[13]),
	.Z(N81));
   CKAN2D1BWP30P140LVT U50 (.A1(FE_OCPN1467_n1),
	.A2(wire_tree_level_0__i_data_latch[12]),
	.Z(N80));
   CKAN2D1BWP30P140LVT U51 (.A1(FE_OCPN1467_n1),
	.A2(wire_tree_level_0__i_data_latch[11]),
	.Z(N79));
   CKAN2D1BWP30P140LVT U52 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_0__i_data_latch[10]),
	.Z(N78));
   CKAN2D1BWP30P140LVT U53 (.A1(FE_OCPN1467_n1),
	.A2(wire_tree_level_0__i_data_latch[9]),
	.Z(N77));
   CKAN2D1BWP30P140LVT U54 (.A1(FE_OCPN1467_n1),
	.A2(wire_tree_level_0__i_data_latch[8]),
	.Z(N76));
   CKAN2D1BWP30P140LVT U55 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_0__i_data_latch[7]),
	.Z(N75));
   CKAN2D1BWP30P140LVT U56 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_0__i_data_latch[6]),
	.Z(N74));
   CKAN2D1BWP30P140LVT U57 (.A1(FE_OCPN1374_FE_OFN752_n1),
	.A2(wire_tree_level_0__i_data_latch[5]),
	.Z(N73));
   CKAN2D1BWP30P140LVT U58 (.A1(FE_OCPN1374_FE_OFN752_n1),
	.A2(wire_tree_level_0__i_data_latch[4]),
	.Z(N72));
   CKAN2D1BWP30P140LVT U59 (.A1(FE_OCPN1374_FE_OFN752_n1),
	.A2(wire_tree_level_0__i_data_latch[3]),
	.Z(N71));
   CKAN2D0BWP30P140LVT U60 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_0__i_data_latch[2]),
	.Z(N70));
   CKAN2D1BWP30P140LVT U61 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_0__i_data_latch[1]),
	.Z(N69));
   CKAN2D1BWP30P140LVT U62 (.A1(FE_OCPN1374_FE_OFN752_n1),
	.A2(wire_tree_level_0__i_data_latch[0]),
	.Z(N68));
   CKAN2D1BWP30P140LVT U63 (.A1(FE_OCPN1469_n1),
	.A2(wire_tree_level_0__i_valid_latch_0_),
	.Z(N101));
   CKAN2D1BWP30P140LVT U64 (.A1(FE_OCPN1467_n1),
	.A2(wire_tree_level_0__i_data_latch[29]),
	.Z(N97));
   CKAN2D1BWP30P140LVT U65 (.A1(FE_OCPN1374_FE_OFN752_n1),
	.A2(wire_tree_level_0__i_data_latch[28]),
	.Z(N96));
   CKAN2D1BWP30P140LVT U66 (.A1(FE_OCPN1375_FE_OFN344_n1),
	.A2(wire_tree_level_0__i_data_latch[27]),
	.Z(N95));
   CKAN2D0BWP30P140LVT U67 (.A1(FE_OCPN1375_FE_OFN344_n1),
	.A2(wire_tree_level_0__i_data_latch[26]),
	.Z(N94));
   CKAN2D1BWP30P140LVT U68 (.A1(FE_OCPN1375_FE_OFN344_n1),
	.A2(wire_tree_level_0__i_data_latch[25]),
	.Z(N93));
   CKAN2D1BWP30P140LVT U69 (.A1(FE_OCPN1375_FE_OFN344_n1),
	.A2(wire_tree_level_0__i_data_latch[24]),
	.Z(N92));
   CKAN2D1BWP30P140LVT U70 (.A1(FE_OCPN1469_n1),
	.A2(wire_tree_level_1__i_valid_latch[1]),
	.Z(N233));
   CKAN2D0BWP30P140LVT U71 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_2__i_data_latch[31]),
	.Z(N297));
   CKAN2D0BWP30P140LVT U72 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_2__i_data_latch[30]),
	.Z(N296));
   CKAN2D1BWP30P140LVT U73 (.A1(FE_OCPN1467_n1),
	.A2(wire_tree_level_2__i_data_latch[29]),
	.Z(N295));
   CKAN2D0BWP30P140LVT U74 (.A1(FE_OCPN1374_FE_OFN752_n1),
	.A2(wire_tree_level_2__i_data_latch[28]),
	.Z(N294));
   CKAN2D0BWP30P140LVT U75 (.A1(FE_OCPN1466_n1),
	.A2(wire_tree_level_2__i_data_latch[27]),
	.Z(N293));
   CKAN2D0BWP30P140LVT U76 (.A1(FE_OCPN1466_n1),
	.A2(wire_tree_level_2__i_data_latch[26]),
	.Z(N292));
   CKAN2D0BWP30P140LVT U77 (.A1(FE_OCPN1466_n1),
	.A2(wire_tree_level_2__i_data_latch[25]),
	.Z(N291));
   CKAN2D0BWP30P140LVT U78 (.A1(FE_OCPN1466_n1),
	.A2(wire_tree_level_2__i_data_latch[24]),
	.Z(N290));
   CKAN2D0BWP30P140LVT U79 (.A1(FE_OCPN1466_n1),
	.A2(wire_tree_level_2__i_data_latch[23]),
	.Z(N289));
   CKAN2D0BWP30P140LVT U80 (.A1(FE_OCPN1466_n1),
	.A2(wire_tree_level_2__i_data_latch[22]),
	.Z(N288));
   CKAN2D0BWP30P140LVT U81 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_2__i_data_latch[21]),
	.Z(N287));
   CKAN2D0BWP30P140LVT U82 (.A1(FE_OCPN1466_n1),
	.A2(wire_tree_level_2__i_data_latch[20]),
	.Z(N286));
   CKAN2D0BWP30P140LVT U83 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_1__i_data_latch[31]),
	.Z(N165));
   CKAN2D0BWP30P140LVT U84 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_1__i_data_latch[30]),
	.Z(N164));
   CKAN2D0BWP30P140LVT U85 (.A1(FE_OCPN1467_n1),
	.A2(wire_tree_level_1__i_data_latch[29]),
	.Z(N163));
   CKAN2D0BWP30P140LVT U86 (.A1(FE_OCPN1374_FE_OFN752_n1),
	.A2(wire_tree_level_1__i_data_latch[28]),
	.Z(N162));
   CKAN2D0BWP30P140LVT U87 (.A1(FE_OCPN1466_n1),
	.A2(wire_tree_level_1__i_data_latch[27]),
	.Z(N161));
   CKAN2D0BWP30P140LVT U88 (.A1(FE_OCPN1466_n1),
	.A2(wire_tree_level_1__i_data_latch[26]),
	.Z(N160));
   CKAN2D0BWP30P140LVT U89 (.A1(FE_OCPN1466_n1),
	.A2(wire_tree_level_1__i_data_latch[25]),
	.Z(N159));
   CKAN2D0BWP30P140LVT U90 (.A1(FE_OCPN1466_n1),
	.A2(wire_tree_level_1__i_data_latch[24]),
	.Z(N158));
   CKAN2D0BWP30P140LVT U91 (.A1(FE_OCPN1466_n1),
	.A2(wire_tree_level_1__i_data_latch[23]),
	.Z(N157));
   CKAN2D0BWP30P140LVT U92 (.A1(FE_OCPN1466_n1),
	.A2(wire_tree_level_1__i_data_latch[22]),
	.Z(N156));
   CKAN2D0BWP30P140LVT U93 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_1__i_data_latch[21]),
	.Z(N155));
   CKAN2D0BWP30P140LVT U94 (.A1(FE_OCPN1466_n1),
	.A2(wire_tree_level_1__i_data_latch[20]),
	.Z(N154));
   CKAN2D0BWP30P140LVT U95 (.A1(FE_OCPN1466_n1),
	.A2(wire_tree_level_1__i_data_latch[19]),
	.Z(N153));
   CKAN2D0BWP30P140LVT U96 (.A1(FE_OCPN1467_n1),
	.A2(wire_tree_level_1__i_data_latch[18]),
	.Z(N152));
   CKAN2D0BWP30P140LVT U97 (.A1(FE_OCPN1374_FE_OFN752_n1),
	.A2(wire_tree_level_1__i_data_latch[17]),
	.Z(N151));
   CKAN2D0BWP30P140LVT U98 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_1__i_data_latch[16]),
	.Z(N150));
   CKAN2D0BWP30P140LVT U99 (.A1(FE_OCPN1374_FE_OFN752_n1),
	.A2(wire_tree_level_1__i_data_latch[15]),
	.Z(N149));
   CKAN2D1BWP30P140LVT U100 (.A1(FE_OCPN1374_FE_OFN752_n1),
	.A2(wire_tree_level_1__i_data_latch[14]),
	.Z(N148));
   CKAN2D0BWP30P140LVT U101 (.A1(FE_OCPN1467_n1),
	.A2(wire_tree_level_1__i_data_latch[13]),
	.Z(N147));
   CKAN2D0BWP30P140LVT U102 (.A1(FE_OCPN1467_n1),
	.A2(wire_tree_level_1__i_data_latch[12]),
	.Z(N146));
   CKAN2D0BWP30P140LVT U103 (.A1(FE_OCPN1467_n1),
	.A2(wire_tree_level_1__i_data_latch[11]),
	.Z(N145));
   CKAN2D0BWP30P140LVT U104 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_1__i_data_latch[10]),
	.Z(N144));
   CKAN2D0BWP30P140LVT U105 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_1__i_data_latch[9]),
	.Z(N143));
   CKAN2D0BWP30P140LVT U106 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_1__i_data_latch[8]),
	.Z(N142));
   CKAN2D0BWP30P140LVT U107 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_1__i_data_latch[7]),
	.Z(N141));
   CKAN2D0BWP30P140LVT U108 (.A1(FE_OCPN1464_n1),
	.A2(wire_tree_level_1__i_data_latch[6]),
	.Z(N140));
   CKAN2D0BWP30P140LVT U109 (.A1(FE_OCPN1464_n1),
	.A2(wire_tree_level_1__i_data_latch[5]),
	.Z(N139));
   CKAN2D0BWP30P140LVT U110 (.A1(FE_OCPN1464_n1),
	.A2(wire_tree_level_1__i_data_latch[4]),
	.Z(N138));
   CKAN2D0BWP30P140LVT U111 (.A1(FE_OCPN1464_n1),
	.A2(wire_tree_level_1__i_data_latch[3]),
	.Z(N137));
   CKAN2D0BWP30P140LVT U112 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_1__i_data_latch[2]),
	.Z(N136));
   CKAN2D0BWP30P140LVT U113 (.A1(FE_OCPN1374_FE_OFN752_n1),
	.A2(wire_tree_level_1__i_data_latch[1]),
	.Z(N135));
   CKAN2D0BWP30P140LVT U114 (.A1(FE_OCPN1374_FE_OFN752_n1),
	.A2(wire_tree_level_1__i_data_latch[0]),
	.Z(N134));
   CKAN2D0BWP30P140LVT U115 (.A1(FE_OCPN1469_n1),
	.A2(wire_tree_level_1__i_valid_latch[0]),
	.Z(N167));
   CKAN2D1BWP30P140LVT U116 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_1__i_data_latch[60]),
	.Z(N228));
   CKAN2D1BWP30P140LVT U117 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_1__i_data_latch[59]),
	.Z(N227));
   CKAN2D1BWP30P140LVT U118 (.A1(FE_OCPN1469_n1),
	.A2(wire_tree_level_1__i_data_latch[58]),
	.Z(N226));
   CKAN2D1BWP30P140LVT U119 (.A1(FE_OCPN1469_n1),
	.A2(wire_tree_level_1__i_data_latch[57]),
	.Z(N225));
   CKAN2D1BWP30P140LVT U120 (.A1(FE_OCPN1469_n1),
	.A2(wire_tree_level_1__i_data_latch[56]),
	.Z(N224));
   CKAN2D1BWP30P140LVT U121 (.A1(FE_OCPN1469_n1),
	.A2(wire_tree_level_1__i_data_latch[55]),
	.Z(N223));
   CKAN2D1BWP30P140LVT U122 (.A1(FE_OCPN1469_n1),
	.A2(wire_tree_level_1__i_data_latch[54]),
	.Z(N222));
   CKAN2D1BWP30P140LVT U123 (.A1(FE_OCPN1469_n1),
	.A2(wire_tree_level_1__i_data_latch[53]),
	.Z(N221));
   CKAN2D1BWP30P140LVT U124 (.A1(FE_OCPN1469_n1),
	.A2(wire_tree_level_1__i_data_latch[52]),
	.Z(N220));
   CKAN2D1BWP30P140LVT U125 (.A1(FE_OCPN1469_n1),
	.A2(wire_tree_level_1__i_data_latch[51]),
	.Z(N219));
   CKAN2D0BWP30P140LVT U126 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_1__i_data_latch[50]),
	.Z(N218));
   CKAN2D1BWP30P140LVT U127 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_1__i_data_latch[49]),
	.Z(N217));
   CKAN2D1BWP30P140LVT U128 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_1__i_data_latch[48]),
	.Z(N216));
   CKAN2D1BWP30P140LVT U129 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_1__i_data_latch[47]),
	.Z(N215));
   CKAN2D1BWP30P140LVT U130 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_1__i_data_latch[46]),
	.Z(N214));
   CKAN2D1BWP30P140LVT U131 (.A1(FE_OCPN1470_n1),
	.A2(wire_tree_level_1__i_data_latch[45]),
	.Z(N213));
   CKAN2D1BWP30P140LVT U132 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_1__i_data_latch[44]),
	.Z(N212));
   CKAN2D1BWP30P140LVT U133 (.A1(FE_OCPN1470_n1),
	.A2(wire_tree_level_1__i_data_latch[43]),
	.Z(N211));
   CKAN2D1BWP30P140LVT U134 (.A1(FE_OCPN1465_n1),
	.A2(wire_tree_level_1__i_data_latch[42]),
	.Z(N210));
   CKAN2D1BWP30P140LVT U135 (.A1(FE_OCPN1470_n1),
	.A2(wire_tree_level_1__i_data_latch[41]),
	.Z(N209));
   CKAN2D1BWP30P140LVT U136 (.A1(FE_OCPN1470_n1),
	.A2(wire_tree_level_1__i_data_latch[40]),
	.Z(N208));
   CKAN2D1BWP30P140LVT U137 (.A1(FE_OCPN1464_n1),
	.A2(wire_tree_level_1__i_data_latch[39]),
	.Z(N207));
   CKAN2D0BWP30P140LVT U138 (.A1(FE_OCPN1465_n1),
	.A2(wire_tree_level_1__i_data_latch[38]),
	.Z(N206));
   CKAN2D0BWP30P140LVT U139 (.A1(FE_OCPN1465_n1),
	.A2(wire_tree_level_1__i_data_latch[37]),
	.Z(N205));
   CKAN2D0BWP30P140LVT U140 (.A1(FE_OCPN1465_n1),
	.A2(wire_tree_level_1__i_data_latch[36]),
	.Z(N204));
   CKAN2D0BWP30P140LVT U141 (.A1(FE_OCPN1465_n1),
	.A2(wire_tree_level_1__i_data_latch[35]),
	.Z(N203));
   CKAN2D1BWP30P140LVT U142 (.A1(FE_OCPN1465_n1),
	.A2(wire_tree_level_1__i_data_latch[34]),
	.Z(N202));
   CKAN2D1BWP30P140LVT U143 (.A1(FE_OCPN1470_n1),
	.A2(wire_tree_level_1__i_data_latch[33]),
	.Z(N201));
   CKAN2D1BWP30P140LVT U144 (.A1(FE_OCPN1470_n1),
	.A2(wire_tree_level_1__i_data_latch[32]),
	.Z(N200));
   CKAN2D1BWP30P140LVT U145 (.A1(FE_OCPN1470_n1),
	.A2(wire_tree_level_1__i_data_latch[63]),
	.Z(N231));
   CKAN2D1BWP30P140LVT U146 (.A1(FE_OCPN1470_n1),
	.A2(wire_tree_level_1__i_data_latch[62]),
	.Z(N230));
   CKAN2D1BWP30P140LVT U147 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_1__i_data_latch[61]),
	.Z(N229));
   CKAN2D0BWP30P140LVT U148 (.A1(FE_OCPN1469_n1),
	.A2(wire_tree_level_2__i_data_latch[118]),
	.Z(N486));
   CKAN2D0BWP30P140LVT U149 (.A1(FE_OCPN1469_n1),
	.A2(wire_tree_level_2__i_data_latch[117]),
	.Z(N485));
   CKAN2D0BWP30P140LVT U150 (.A1(FE_OCPN1469_n1),
	.A2(wire_tree_level_2__i_data_latch[116]),
	.Z(N484));
   CKAN2D0BWP30P140LVT U151 (.A1(FE_OCPN1469_n1),
	.A2(wire_tree_level_2__i_data_latch[115]),
	.Z(N483));
   CKAN2D0BWP30P140LVT U152 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_2__i_data_latch[114]),
	.Z(N482));
   CKAN2D0BWP30P140LVT U153 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_2__i_data_latch[113]),
	.Z(N481));
   CKAN2D0BWP30P140LVT U154 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_2__i_data_latch[112]),
	.Z(N480));
   CKAN2D0BWP30P140LVT U155 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_2__i_data_latch[111]),
	.Z(N479));
   CKAN2D0BWP30P140LVT U156 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_2__i_data_latch[110]),
	.Z(N478));
   CKAN2D0BWP30P140LVT U157 (.A1(FE_OCPN1470_n1),
	.A2(wire_tree_level_2__i_data_latch[109]),
	.Z(N477));
   CKAN2D0BWP30P140LVT U158 (.A1(FE_OCPN1470_n1),
	.A2(wire_tree_level_2__i_data_latch[108]),
	.Z(N476));
   CKAN2D0BWP30P140LVT U159 (.A1(FE_OCPN1470_n1),
	.A2(wire_tree_level_2__i_data_latch[107]),
	.Z(N475));
   CKAN2D0BWP30P140LVT U160 (.A1(FE_OCPN1470_n1),
	.A2(wire_tree_level_2__i_data_latch[106]),
	.Z(N474));
   CKAN2D0BWP30P140LVT U161 (.A1(FE_OCPN1470_n1),
	.A2(wire_tree_level_2__i_data_latch[105]),
	.Z(N473));
   CKAN2D0BWP30P140LVT U162 (.A1(FE_OCPN1470_n1),
	.A2(wire_tree_level_2__i_data_latch[104]),
	.Z(N472));
   CKAN2D0BWP30P140LVT U163 (.A1(FE_OCPN1465_n1),
	.A2(wire_tree_level_2__i_data_latch[103]),
	.Z(N471));
   CKAN2D0BWP30P140LVT U164 (.A1(FE_OCPN1465_n1),
	.A2(wire_tree_level_2__i_data_latch[102]),
	.Z(N470));
   CKAN2D0BWP30P140LVT U165 (.A1(FE_OCPN1465_n1),
	.A2(wire_tree_level_2__i_data_latch[101]),
	.Z(N469));
   CKAN2D0BWP30P140LVT U166 (.A1(FE_OCPN1465_n1),
	.A2(wire_tree_level_2__i_data_latch[100]),
	.Z(N468));
   CKAN2D0BWP30P140LVT U167 (.A1(FE_OCPN1465_n1),
	.A2(wire_tree_level_2__i_data_latch[99]),
	.Z(N467));
   CKAN2D0BWP30P140LVT U168 (.A1(FE_OCPN1465_n1),
	.A2(wire_tree_level_2__i_data_latch[98]),
	.Z(N466));
   CKAN2D0BWP30P140LVT U169 (.A1(FE_OCPN1470_n1),
	.A2(wire_tree_level_2__i_data_latch[97]),
	.Z(N465));
   CKAN2D0BWP30P140LVT U170 (.A1(FE_OCPN1470_n1),
	.A2(wire_tree_level_2__i_data_latch[96]),
	.Z(N464));
   CKAN2D0BWP30P140LVT U171 (.A1(FE_OCPN1469_n1),
	.A2(wire_tree_level_2__i_valid_latch[3]),
	.Z(N497));
   CKAN2D0BWP30P140LVT U172 (.A1(FE_OCPN1469_n1),
	.A2(wire_tree_level_2__i_valid_latch[0]),
	.Z(N299));
   CKAN2D0BWP30P140LVT U173 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_2__i_data_latch[63]),
	.Z(N363));
   CKAN2D0BWP30P140LVT U174 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_2__i_data_latch[62]),
	.Z(N362));
   CKAN2D0BWP30P140LVT U175 (.A1(FE_OCPN1467_n1),
	.A2(wire_tree_level_2__i_data_latch[61]),
	.Z(N361));
   CKAN2D0BWP30P140LVT U176 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_2__i_data_latch[9]),
	.Z(N275));
   CKAN2D0BWP30P140LVT U177 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_2__i_data_latch[8]),
	.Z(N274));
   CKAN2D0BWP30P140LVT U178 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_2__i_data_latch[7]),
	.Z(N273));
   CKAN2D0BWP30P140LVT U179 (.A1(FE_OCPN1464_n1),
	.A2(wire_tree_level_2__i_data_latch[6]),
	.Z(N272));
   CKAN2D0BWP30P140LVT U180 (.A1(FE_OCPN1464_n1),
	.A2(wire_tree_level_2__i_data_latch[5]),
	.Z(N271));
   CKAN2D0BWP30P140LVT U181 (.A1(FE_OCPN1464_n1),
	.A2(wire_tree_level_2__i_data_latch[4]),
	.Z(N270));
   CKAN2D0BWP30P140LVT U182 (.A1(FE_OCPN1464_n1),
	.A2(wire_tree_level_2__i_data_latch[3]),
	.Z(N269));
   CKAN2D1BWP30P140LVT U183 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_2__i_data_latch[2]),
	.Z(N268));
   CKAN2D0BWP30P140LVT U184 (.A1(FE_OCPN1374_FE_OFN752_n1),
	.A2(wire_tree_level_2__i_data_latch[1]),
	.Z(N267));
   CKAN2D0BWP30P140LVT U185 (.A1(FE_OCPN1374_FE_OFN752_n1),
	.A2(wire_tree_level_2__i_data_latch[0]),
	.Z(N266));
   CKAN2D0BWP30P140LVT U186 (.A1(FE_OCPN1466_n1),
	.A2(wire_tree_level_2__i_data_latch[19]),
	.Z(N285));
   CKAN2D0BWP30P140LVT U187 (.A1(FE_OCPN1467_n1),
	.A2(wire_tree_level_2__i_data_latch[18]),
	.Z(N284));
   CKAN2D0BWP30P140LVT U188 (.A1(FE_OCPN1374_FE_OFN752_n1),
	.A2(wire_tree_level_2__i_data_latch[17]),
	.Z(N283));
   CKAN2D0BWP30P140LVT U189 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_2__i_data_latch[16]),
	.Z(N282));
   CKAN2D0BWP30P140LVT U190 (.A1(FE_OCPN1374_FE_OFN752_n1),
	.A2(wire_tree_level_2__i_data_latch[15]),
	.Z(N281));
   CKAN2D0BWP30P140LVT U191 (.A1(FE_OCPN1374_FE_OFN752_n1),
	.A2(wire_tree_level_2__i_data_latch[14]),
	.Z(N280));
   CKAN2D0BWP30P140LVT U192 (.A1(FE_OCPN1467_n1),
	.A2(wire_tree_level_2__i_data_latch[13]),
	.Z(N279));
   CKAN2D0BWP30P140LVT U193 (.A1(FE_OCPN1467_n1),
	.A2(wire_tree_level_2__i_data_latch[12]),
	.Z(N278));
   CKAN2D0BWP30P140LVT U194 (.A1(FE_OCPN1467_n1),
	.A2(wire_tree_level_2__i_data_latch[11]),
	.Z(N277));
   CKAN2D0BWP30P140LVT U195 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_2__i_data_latch[10]),
	.Z(N276));
   CKAN2D0BWP30P140LVT U196 (.A1(FE_OCPN1466_n1),
	.A2(wire_tree_level_2__i_data_latch[59]),
	.Z(N359));
   CKAN2D1BWP30P140LVT U197 (.A1(FE_OCPN1466_n1),
	.A2(wire_tree_level_2__i_data_latch[58]),
	.Z(N358));
   CKAN2D0BWP30P140LVT U198 (.A1(FE_OCPN1466_n1),
	.A2(wire_tree_level_2__i_data_latch[57]),
	.Z(N357));
   CKAN2D0BWP30P140LVT U199 (.A1(FE_OCPN1466_n1),
	.A2(wire_tree_level_2__i_data_latch[56]),
	.Z(N356));
   CKAN2D0BWP30P140LVT U200 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_2__i_data_latch[55]),
	.Z(N355));
   CKAN2D0BWP30P140LVT U201 (.A1(FE_OCPN1466_n1),
	.A2(wire_tree_level_2__i_data_latch[54]),
	.Z(N354));
   CKAN2D0BWP30P140LVT U202 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_2__i_data_latch[53]),
	.Z(N353));
   CKAN2D1BWP30P140LVT U203 (.A1(FE_OCPN1466_n1),
	.A2(wire_tree_level_2__i_data_latch[52]),
	.Z(N352));
   CKAN2D1BWP30P140LVT U204 (.A1(FE_OCPN1466_n1),
	.A2(wire_tree_level_2__i_data_latch[51]),
	.Z(N351));
   CKAN2D0BWP30P140LVT U205 (.A1(FE_OCPN1467_n1),
	.A2(wire_tree_level_2__i_data_latch[50]),
	.Z(N350));
   CKAN2D0BWP30P140LVT U206 (.A1(FE_OCPN1374_FE_OFN752_n1),
	.A2(wire_tree_level_2__i_data_latch[49]),
	.Z(N349));
   CKAN2D0BWP30P140LVT U207 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_2__i_data_latch[48]),
	.Z(N348));
   CKAN2D0BWP30P140LVT U208 (.A1(FE_OCPN1374_FE_OFN752_n1),
	.A2(wire_tree_level_2__i_data_latch[47]),
	.Z(N347));
   CKAN2D0BWP30P140LVT U209 (.A1(FE_OCPN1374_FE_OFN752_n1),
	.A2(wire_tree_level_2__i_data_latch[46]),
	.Z(N346));
   CKAN2D0BWP30P140LVT U210 (.A1(FE_OCPN1467_n1),
	.A2(wire_tree_level_2__i_data_latch[45]),
	.Z(N345));
   CKAN2D0BWP30P140LVT U211 (.A1(FE_OCPN1467_n1),
	.A2(wire_tree_level_2__i_data_latch[44]),
	.Z(N344));
   CKAN2D0BWP30P140LVT U212 (.A1(FE_OCPN1467_n1),
	.A2(wire_tree_level_2__i_data_latch[43]),
	.Z(N343));
   CKAN2D0BWP30P140LVT U213 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_2__i_data_latch[42]),
	.Z(N342));
   CKAN2D0BWP30P140LVT U214 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_2__i_data_latch[41]),
	.Z(N341));
   CKAN2D0BWP30P140LVT U215 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_2__i_data_latch[40]),
	.Z(N340));
   CKAN2D0BWP30P140LVT U216 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_2__i_data_latch[39]),
	.Z(N339));
   CKAN2D0BWP30P140LVT U217 (.A1(FE_OCPN1464_n1),
	.A2(wire_tree_level_2__i_data_latch[38]),
	.Z(N338));
   CKAN2D0BWP30P140LVT U218 (.A1(FE_OCPN1464_n1),
	.A2(wire_tree_level_2__i_data_latch[37]),
	.Z(N337));
   CKAN2D0BWP30P140LVT U219 (.A1(FE_OCPN1464_n1),
	.A2(wire_tree_level_2__i_data_latch[36]),
	.Z(N336));
   CKAN2D1BWP30P140LVT U220 (.A1(FE_OFN344_n1),
	.A2(wire_tree_level_2__i_data_latch[34]),
	.Z(N334));
   CKAN2D0BWP30P140LVT U221 (.A1(FE_OCPN1374_FE_OFN752_n1),
	.A2(wire_tree_level_2__i_data_latch[33]),
	.Z(N333));
   CKAN2D1BWP30P140LVT U222 (.A1(FE_OCPN1374_FE_OFN752_n1),
	.A2(wire_tree_level_2__i_data_latch[32]),
	.Z(N332));
   CKAN2D1BWP30P140LVT U223 (.A1(FE_OCPN1469_n1),
	.A2(wire_tree_level_2__i_valid_latch[1]),
	.Z(N365));
   CKAN2D0BWP30P140LVT U224 (.A1(FE_OCPN1374_FE_OFN752_n1),
	.A2(wire_tree_level_2__i_data_latch[60]),
	.Z(N360));
   CKAN2D0BWP30P140LVT U225 (.A1(FE_OFN343_n1),
	.A2(wire_tree_level_2__i_data_latch[95]),
	.Z(N429));
   CKAN2D1BWP30P140LVT U226 (.A1(FE_OFN343_n1),
	.A2(wire_tree_level_2__i_data_latch[94]),
	.Z(N428));
   CKAN2D1BWP30P140LVT U227 (.A1(FE_OFN343_n1),
	.A2(wire_tree_level_2__i_data_latch[93]),
	.Z(N427));
   CKAN2D1BWP30P140LVT U228 (.A1(FE_OFN343_n1),
	.A2(wire_tree_level_2__i_data_latch[92]),
	.Z(N426));
   CKAN2D1BWP30P140LVT U229 (.A1(FE_OCPN1468_n1),
	.A2(wire_tree_level_2__i_data_latch[91]),
	.Z(N425));
   CKAN2D1BWP30P140LVT U230 (.A1(FE_OCPN1468_n1),
	.A2(wire_tree_level_2__i_data_latch[90]),
	.Z(N424));
   CKAN2D1BWP30P140LVT U231 (.A1(FE_OCPN1468_n1),
	.A2(wire_tree_level_2__i_data_latch[89]),
	.Z(N423));
   CKAN2D1BWP30P140LVT U232 (.A1(FE_OCPN1468_n1),
	.A2(wire_tree_level_2__i_data_latch[88]),
	.Z(N422));
   CKAN2D1BWP30P140LVT U233 (.A1(FE_OCPN1468_n1),
	.A2(wire_tree_level_2__i_data_latch[87]),
	.Z(N421));
   CKAN2D1BWP30P140LVT U234 (.A1(FE_OCPN1468_n1),
	.A2(wire_tree_level_2__i_data_latch[86]),
	.Z(N420));
   CKAN2D1BWP30P140LVT U235 (.A1(FE_OCPN1468_n1),
	.A2(wire_tree_level_2__i_data_latch[85]),
	.Z(N419));
   CKAN2D1BWP30P140LVT U236 (.A1(FE_OCPN1468_n1),
	.A2(wire_tree_level_2__i_data_latch[84]),
	.Z(N418));
   CKAN2D1BWP30P140LVT U237 (.A1(FE_OCPN1469_n1),
	.A2(wire_tree_level_2__i_data_latch[83]),
	.Z(N417));
   CKAN2D1BWP30P140LVT U238 (.A1(FE_OCPN1468_n1),
	.A2(wire_tree_level_2__i_data_latch[82]),
	.Z(N416));
   CKAN2D1BWP30P140LVT U239 (.A1(FE_OFN343_n1),
	.A2(wire_tree_level_2__i_data_latch[81]),
	.Z(N415));
   CKAN2D1BWP30P140LVT U240 (.A1(FE_OFN343_n1),
	.A2(wire_tree_level_2__i_data_latch[80]),
	.Z(N414));
   CKAN2D1BWP30P140LVT U241 (.A1(FE_OFN343_n1),
	.A2(wire_tree_level_2__i_data_latch[79]),
	.Z(N413));
   CKAN2D1BWP30P140LVT U242 (.A1(FE_OFN343_n1),
	.A2(wire_tree_level_2__i_data_latch[78]),
	.Z(N412));
   CKAN2D1BWP30P140LVT U243 (.A1(FE_OFN343_n1),
	.A2(wire_tree_level_2__i_data_latch[77]),
	.Z(N411));
   CKAN2D1BWP30P140LVT U244 (.A1(FE_OFN343_n1),
	.A2(wire_tree_level_2__i_data_latch[76]),
	.Z(N410));
   CKAN2D1BWP30P140LVT U245 (.A1(FE_OFN343_n1),
	.A2(wire_tree_level_2__i_data_latch[75]),
	.Z(N409));
   CKAN2D1BWP30P140LVT U246 (.A1(FE_OFN343_n1),
	.A2(wire_tree_level_2__i_data_latch[74]),
	.Z(N408));
   CKAN2D1BWP30P140LVT U247 (.A1(FE_OFN343_n1),
	.A2(wire_tree_level_2__i_data_latch[73]),
	.Z(N407));
   CKAN2D1BWP30P140LVT U248 (.A1(FE_OFN343_n1),
	.A2(wire_tree_level_2__i_data_latch[72]),
	.Z(N406));
   CKAN2D1BWP30P140LVT U249 (.A1(FE_OFN343_n1),
	.A2(wire_tree_level_2__i_data_latch[71]),
	.Z(N405));
   CKAN2D1BWP30P140LVT U250 (.A1(FE_OFN343_n1),
	.A2(wire_tree_level_2__i_data_latch[70]),
	.Z(N404));
   CKAN2D1BWP30P140LVT U251 (.A1(FE_OFN343_n1),
	.A2(wire_tree_level_2__i_data_latch[69]),
	.Z(N403));
   CKAN2D1BWP30P140LVT U252 (.A1(FE_OFN343_n1),
	.A2(wire_tree_level_2__i_data_latch[68]),
	.Z(N402));
   CKAN2D1BWP30P140LVT U253 (.A1(FE_OFN343_n1),
	.A2(wire_tree_level_2__i_data_latch[67]),
	.Z(N401));
   CKAN2D1BWP30P140LVT U254 (.A1(FE_OFN343_n1),
	.A2(wire_tree_level_2__i_data_latch[66]),
	.Z(N400));
   CKAN2D1BWP30P140LVT U255 (.A1(FE_OFN343_n1),
	.A2(wire_tree_level_2__i_data_latch[65]),
	.Z(N399));
   CKAN2D1BWP30P140LVT U256 (.A1(FE_OFN343_n1),
	.A2(wire_tree_level_2__i_data_latch[64]),
	.Z(N398));
   CKAN2D1BWP30P140LVT U257 (.A1(FE_OCPN1469_n1),
	.A2(wire_tree_level_2__i_valid_latch[2]),
	.Z(N431));
   CKAN2D0BWP30P140LVT U258 (.A1(FE_OCPN1470_n1),
	.A2(wire_tree_level_2__i_data_latch[127]),
	.Z(N495));
   CKAN2D0BWP30P140LVT U259 (.A1(FE_OCPN1470_n1),
	.A2(wire_tree_level_2__i_data_latch[126]),
	.Z(N494));
   CKAN2D0BWP30P140LVT U260 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_2__i_data_latch[125]),
	.Z(N493));
   CKAN2D0BWP30P140LVT U261 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_2__i_data_latch[124]),
	.Z(N492));
   CKAN2D0BWP30P140LVT U262 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_2__i_data_latch[123]),
	.Z(N491));
   CKAN2D0BWP30P140LVT U263 (.A1(FE_OFN341_n1),
	.A2(wire_tree_level_2__i_data_latch[122]),
	.Z(N490));
   CKAN2D0BWP30P140LVT U264 (.A1(FE_OCPN1469_n1),
	.A2(wire_tree_level_2__i_data_latch[121]),
	.Z(N489));
   CKAN2D0BWP30P140LVT U265 (.A1(FE_OCPN1469_n1),
	.A2(wire_tree_level_2__i_data_latch[120]),
	.Z(N488));
   CKAN2D0BWP30P140LVT U266 (.A1(FE_OCPN1469_n1),
	.A2(wire_tree_level_2__i_data_latch[119]),
	.Z(N487));
   CKAN2D0BWP30P140LVT U267 (.A1(FE_OCPN1464_n1),
	.A2(wire_tree_level_2__i_data_latch[35]),
	.Z(N335));
endmodule
