
module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_0 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  BUFFD2BWP30P140 U3 ( .I(n41), .Z(n1) );
  INVD2BWP30P140 U4 ( .I(n41), .ZN(n39) );
  ND2D1BWP30P140 U5 ( .A1(n22), .A2(i_cmd[1]), .ZN(n9) );
  ND2D2BWP30P140 U6 ( .A1(n33), .A2(n23), .ZN(n6) );
  INVD3BWP30P140 U7 ( .I(n2), .ZN(n32) );
  CKND2D4BWP30P140 U8 ( .A1(i_cmd[0]), .A2(n21), .ZN(n5) );
  OAI22D1BWP30P140 U9 ( .A1(n95), .A2(n10), .B1(n36), .B2(n28), .ZN(N291) );
  CKND2D2BWP30P140 U10 ( .A1(i_valid[0]), .A2(n21), .ZN(n2) );
  INR2D6BWP30P140 U11 ( .A1(n9), .B1(n8), .ZN(n29) );
  INVD3BWP30P140 U12 ( .I(i_valid[1]), .ZN(n22) );
  ND2OPTPAD4BWP30P140 U13 ( .A1(n3), .A2(n24), .ZN(n41) );
  ND2D1BWP30P140 U14 ( .A1(n31), .A2(n30), .ZN(N290) );
  ND2OPTIBD1BWP30P140 U15 ( .A1(n29), .A2(i_data_bus[35]), .ZN(n31) );
  ND2OPTIBD1BWP30P140 U16 ( .A1(n93), .A2(i_data_bus[3]), .ZN(n30) );
  OAI22D1BWP30P140 U17 ( .A1(n95), .A2(n19), .B1(n36), .B2(n49), .ZN(N292) );
  OAI22D1BWP30P140 U18 ( .A1(n95), .A2(n18), .B1(n36), .B2(n62), .ZN(N293) );
  OAI22D1BWP30P140 U19 ( .A1(n95), .A2(n17), .B1(n36), .B2(n46), .ZN(N294) );
  OAI22D1BWP30P140 U20 ( .A1(n95), .A2(n16), .B1(n36), .B2(n60), .ZN(N304) );
  OAI22D1BWP30P140 U21 ( .A1(n95), .A2(n12), .B1(n36), .B2(n65), .ZN(N305) );
  OAI22D1BWP30P140 U22 ( .A1(n95), .A2(n13), .B1(n36), .B2(n69), .ZN(N306) );
  OAI22D1BWP30P140 U23 ( .A1(n95), .A2(n14), .B1(n36), .B2(n47), .ZN(N316) );
  OAI22D1BWP30P140 U24 ( .A1(n95), .A2(n11), .B1(n36), .B2(n45), .ZN(N317) );
  OAI22D1BWP30P140 U25 ( .A1(n95), .A2(n15), .B1(n36), .B2(n43), .ZN(N318) );
  OAI22D1BWP30P140 U26 ( .A1(n26), .A2(n10), .B1(n1), .B2(n28), .ZN(N323) );
  OAI22D1BWP30P140 U27 ( .A1(n26), .A2(n90), .B1(n1), .B2(n27), .ZN(N340) );
  OAI22D1BWP30P140 U28 ( .A1(n26), .A2(n79), .B1(n1), .B2(n25), .ZN(N345) );
  INVD3BWP30P140 U29 ( .I(n33), .ZN(n35) );
  NR2OPTPAD2BWP30P140 U30 ( .A1(n35), .A2(n38), .ZN(n3) );
  INVD4BWP30P140 U31 ( .I(i_cmd[1]), .ZN(n33) );
  INVD2BWP30P140 U32 ( .I(n70), .ZN(n26) );
  ND2OPTPAD4BWP30P140 U33 ( .A1(n20), .A2(n21), .ZN(n34) );
  INVD1BWP30P140 U34 ( .I(n38), .ZN(n21) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n4) );
  ND2D1BWP30P140 U36 ( .A1(n4), .A2(i_en), .ZN(n38) );
  INVD2BWP30P140 U37 ( .I(i_cmd[0]), .ZN(n37) );
  ND2OPTIBD8BWP30P140 U38 ( .A1(n32), .A2(n37), .ZN(n36) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[4]), .ZN(n28) );
  INVD2BWP30P140 U40 ( .I(n5), .ZN(n7) );
  INVD2BWP30P140 U41 ( .I(i_valid[0]), .ZN(n23) );
  ND2OPTIBD4BWP30P140 U42 ( .A1(n7), .A2(n6), .ZN(n8) );
  INVD12BWP30P140 U43 ( .I(n29), .ZN(n95) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[36]), .ZN(n10) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[62]), .ZN(n11) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[30]), .ZN(n45) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[50]), .ZN(n12) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[18]), .ZN(n65) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[51]), .ZN(n13) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[19]), .ZN(n69) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[61]), .ZN(n14) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[29]), .ZN(n47) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[63]), .ZN(n15) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[31]), .ZN(n43) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[49]), .ZN(n16) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[17]), .ZN(n60) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[39]), .ZN(n17) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[7]), .ZN(n46) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[38]), .ZN(n18) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[6]), .ZN(n62) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[37]), .ZN(n19) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[5]), .ZN(n49) );
  INR2D4BWP30P140 U63 ( .A1(i_valid[1]), .B1(n33), .ZN(n20) );
  INVD8BWP30P140 U64 ( .I(n34), .ZN(n70) );
  MUX2NOPTD4BWP30P140 U65 ( .I0(n23), .I1(n22), .S(i_cmd[0]), .ZN(n24) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[26]), .ZN(n25) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[21]), .ZN(n27) );
  INVD8BWP30P140 U68 ( .I(n36), .ZN(n93) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[3]), .ZN(n40) );
  OAI21D1BWP30P140 U70 ( .A1(n2), .A2(n35), .B(n26), .ZN(N354) );
  OAI31D1BWP30P140 U71 ( .A1(n38), .A2(n22), .A3(n37), .B(n36), .ZN(N353) );
  INVD4BWP30P140 U72 ( .I(n39), .ZN(n71) );
  MOAI22D1BWP30P140 U73 ( .A1(n40), .A2(n71), .B1(i_data_bus[35]), .B2(n70), 
        .ZN(N322) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[27]), .ZN(n42) );
  BUFFD4BWP30P140 U75 ( .I(n41), .Z(n67) );
  MOAI22D1BWP30P140 U76 ( .A1(n42), .A2(n67), .B1(i_data_bus[59]), .B2(n70), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U77 ( .A1(n43), .A2(n67), .B1(i_data_bus[63]), .B2(n70), 
        .ZN(N350) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[1]), .ZN(n44) );
  MOAI22D1BWP30P140 U79 ( .A1(n44), .A2(n71), .B1(i_data_bus[33]), .B2(n70), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U80 ( .A1(n45), .A2(n67), .B1(i_data_bus[62]), .B2(n70), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U81 ( .A1(n46), .A2(n71), .B1(i_data_bus[39]), .B2(n70), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U82 ( .A1(n47), .A2(n67), .B1(i_data_bus[61]), .B2(n70), 
        .ZN(N348) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[0]), .ZN(n48) );
  MOAI22D1BWP30P140 U84 ( .A1(n48), .A2(n71), .B1(i_data_bus[32]), .B2(n70), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U85 ( .A1(n49), .A2(n71), .B1(i_data_bus[37]), .B2(n70), 
        .ZN(N324) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[9]), .ZN(n50) );
  MOAI22D1BWP30P140 U87 ( .A1(n50), .A2(n67), .B1(i_data_bus[41]), .B2(n70), 
        .ZN(N328) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[22]), .ZN(n51) );
  MOAI22D1BWP30P140 U89 ( .A1(n51), .A2(n67), .B1(i_data_bus[54]), .B2(n70), 
        .ZN(N341) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[10]), .ZN(n52) );
  MOAI22D1BWP30P140 U91 ( .A1(n52), .A2(n71), .B1(i_data_bus[42]), .B2(n70), 
        .ZN(N329) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[11]), .ZN(n53) );
  MOAI22D1BWP30P140 U93 ( .A1(n53), .A2(n67), .B1(i_data_bus[43]), .B2(n70), 
        .ZN(N330) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[24]), .ZN(n54) );
  MOAI22D1BWP30P140 U95 ( .A1(n54), .A2(n67), .B1(i_data_bus[56]), .B2(n70), 
        .ZN(N343) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[12]), .ZN(n55) );
  MOAI22D1BWP30P140 U97 ( .A1(n55), .A2(n71), .B1(i_data_bus[44]), .B2(n70), 
        .ZN(N331) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[13]), .ZN(n56) );
  MOAI22D1BWP30P140 U99 ( .A1(n56), .A2(n67), .B1(i_data_bus[45]), .B2(n70), 
        .ZN(N332) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[14]), .ZN(n57) );
  MOAI22D1BWP30P140 U101 ( .A1(n57), .A2(n71), .B1(i_data_bus[46]), .B2(n70), 
        .ZN(N333) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[15]), .ZN(n58) );
  MOAI22D1BWP30P140 U103 ( .A1(n58), .A2(n67), .B1(i_data_bus[47]), .B2(n70), 
        .ZN(N334) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[16]), .ZN(n59) );
  MOAI22D1BWP30P140 U105 ( .A1(n59), .A2(n71), .B1(i_data_bus[48]), .B2(n70), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U106 ( .A1(n60), .A2(n71), .B1(i_data_bus[49]), .B2(n70), 
        .ZN(N336) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[23]), .ZN(n61) );
  MOAI22D1BWP30P140 U108 ( .A1(n61), .A2(n67), .B1(i_data_bus[55]), .B2(n70), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U109 ( .A1(n62), .A2(n71), .B1(i_data_bus[38]), .B2(n70), 
        .ZN(N325) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[2]), .ZN(n63) );
  MOAI22D1BWP30P140 U111 ( .A1(n63), .A2(n71), .B1(i_data_bus[34]), .B2(n70), 
        .ZN(N321) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[8]), .ZN(n64) );
  MOAI22D1BWP30P140 U113 ( .A1(n64), .A2(n71), .B1(i_data_bus[40]), .B2(n70), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U114 ( .A1(n65), .A2(n71), .B1(i_data_bus[50]), .B2(n70), 
        .ZN(N337) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[20]), .ZN(n66) );
  MOAI22D1BWP30P140 U116 ( .A1(n66), .A2(n67), .B1(i_data_bus[52]), .B2(n70), 
        .ZN(N339) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[28]), .ZN(n68) );
  MOAI22D1BWP30P140 U118 ( .A1(n68), .A2(n67), .B1(i_data_bus[60]), .B2(n70), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U119 ( .A1(n69), .A2(n71), .B1(i_data_bus[51]), .B2(n70), 
        .ZN(N338) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[25]), .ZN(n72) );
  MOAI22D1BWP30P140 U121 ( .A1(n72), .A2(n71), .B1(i_data_bus[57]), .B2(n70), 
        .ZN(N344) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[60]), .ZN(n73) );
  MOAI22D1BWP30P140 U123 ( .A1(n95), .A2(n73), .B1(n93), .B2(i_data_bus[28]), 
        .ZN(N315) );
  INVD1BWP30P140 U124 ( .I(i_data_bus[48]), .ZN(n74) );
  MOAI22D1BWP30P140 U125 ( .A1(n95), .A2(n74), .B1(n93), .B2(i_data_bus[16]), 
        .ZN(N303) );
  INVD1BWP30P140 U126 ( .I(i_data_bus[34]), .ZN(n75) );
  MOAI22D1BWP30P140 U127 ( .A1(n95), .A2(n75), .B1(n93), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140 U128 ( .I(i_data_bus[59]), .ZN(n76) );
  MOAI22D1BWP30P140 U129 ( .A1(n95), .A2(n76), .B1(n93), .B2(i_data_bus[27]), 
        .ZN(N314) );
  INVD1BWP30P140 U130 ( .I(i_data_bus[47]), .ZN(n77) );
  MOAI22D1BWP30P140 U131 ( .A1(n95), .A2(n77), .B1(n93), .B2(i_data_bus[15]), 
        .ZN(N302) );
  INVD1BWP30P140 U132 ( .I(i_data_bus[33]), .ZN(n78) );
  MOAI22D1BWP30P140 U133 ( .A1(n95), .A2(n78), .B1(n93), .B2(i_data_bus[1]), 
        .ZN(N288) );
  INVD1BWP30P140 U134 ( .I(i_data_bus[58]), .ZN(n79) );
  MOAI22D1BWP30P140 U135 ( .A1(n95), .A2(n79), .B1(n93), .B2(i_data_bus[26]), 
        .ZN(N313) );
  INVD1BWP30P140 U136 ( .I(i_data_bus[46]), .ZN(n80) );
  MOAI22D1BWP30P140 U137 ( .A1(n95), .A2(n80), .B1(n93), .B2(i_data_bus[14]), 
        .ZN(N301) );
  INVD1BWP30P140 U138 ( .I(i_data_bus[32]), .ZN(n81) );
  MOAI22D1BWP30P140 U139 ( .A1(n95), .A2(n81), .B1(n93), .B2(i_data_bus[0]), 
        .ZN(N287) );
  INVD1BWP30P140 U140 ( .I(i_data_bus[57]), .ZN(n82) );
  MOAI22D1BWP30P140 U141 ( .A1(n95), .A2(n82), .B1(n93), .B2(i_data_bus[25]), 
        .ZN(N312) );
  INVD1BWP30P140 U142 ( .I(i_data_bus[45]), .ZN(n83) );
  MOAI22D1BWP30P140 U143 ( .A1(n95), .A2(n83), .B1(n93), .B2(i_data_bus[13]), 
        .ZN(N300) );
  INVD1BWP30P140 U144 ( .I(i_data_bus[56]), .ZN(n84) );
  MOAI22D1BWP30P140 U145 ( .A1(n95), .A2(n84), .B1(n93), .B2(i_data_bus[24]), 
        .ZN(N311) );
  INVD1BWP30P140 U146 ( .I(i_data_bus[44]), .ZN(n85) );
  MOAI22D1BWP30P140 U147 ( .A1(n95), .A2(n85), .B1(n93), .B2(i_data_bus[12]), 
        .ZN(N299) );
  INVD1BWP30P140 U148 ( .I(i_data_bus[55]), .ZN(n86) );
  MOAI22D1BWP30P140 U149 ( .A1(n95), .A2(n86), .B1(n93), .B2(i_data_bus[23]), 
        .ZN(N310) );
  INVD1BWP30P140 U150 ( .I(i_data_bus[43]), .ZN(n87) );
  MOAI22D1BWP30P140 U151 ( .A1(n95), .A2(n87), .B1(n93), .B2(i_data_bus[11]), 
        .ZN(N298) );
  INVD1BWP30P140 U152 ( .I(i_data_bus[54]), .ZN(n88) );
  MOAI22D1BWP30P140 U153 ( .A1(n95), .A2(n88), .B1(n93), .B2(i_data_bus[22]), 
        .ZN(N309) );
  INVD1BWP30P140 U154 ( .I(i_data_bus[42]), .ZN(n89) );
  MOAI22D1BWP30P140 U155 ( .A1(n95), .A2(n89), .B1(n93), .B2(i_data_bus[10]), 
        .ZN(N297) );
  INVD1BWP30P140 U156 ( .I(i_data_bus[53]), .ZN(n90) );
  MOAI22D1BWP30P140 U157 ( .A1(n95), .A2(n90), .B1(n93), .B2(i_data_bus[21]), 
        .ZN(N308) );
  INVD1BWP30P140 U158 ( .I(i_data_bus[41]), .ZN(n91) );
  MOAI22D1BWP30P140 U159 ( .A1(n95), .A2(n91), .B1(n93), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140 U160 ( .I(i_data_bus[52]), .ZN(n92) );
  MOAI22D1BWP30P140 U161 ( .A1(n95), .A2(n92), .B1(n93), .B2(i_data_bus[20]), 
        .ZN(N307) );
  INVD1BWP30P140 U162 ( .I(i_data_bus[40]), .ZN(n94) );
  MOAI22D1BWP30P140 U163 ( .A1(n95), .A2(n94), .B1(n93), .B2(i_data_bus[8]), 
        .ZN(N295) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_1 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91;

  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  NR3D0BWP30P140 U3 ( .A1(n52), .A2(n9), .A3(n51), .ZN(n1) );
  INVD1BWP30P140 U4 ( .I(n55), .ZN(n68) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n11), .A2(n10), .ZN(n12) );
  MUX2NUD1BWP30P140 U6 ( .I0(n8), .I1(n52), .S(i_cmd[1]), .ZN(n11) );
  INVD1BWP30P140 U7 ( .I(n3), .ZN(n27) );
  INVD3BWP30P140 U8 ( .I(n14), .ZN(n49) );
  IND2D1BWP30P140 U9 ( .A1(n1), .B1(n26), .ZN(N353) );
  INVD3BWP30P140 U10 ( .I(n14), .ZN(n47) );
  OAI22D1BWP30P140 U11 ( .A1(n26), .A2(n64), .B1(n47), .B2(n21), .ZN(N318) );
  INVD3BWP30P140 U12 ( .I(n68), .ZN(n79) );
  INVD1BWP30P140 U13 ( .I(n89), .ZN(n6) );
  OAI22D1BWP30P140 U14 ( .A1(n50), .A2(n72), .B1(n47), .B2(n44), .ZN(N317) );
  INVD1BWP30P140 U15 ( .I(rst), .ZN(n2) );
  ND2D1BWP30P140 U16 ( .A1(n2), .A2(i_en), .ZN(n51) );
  INVD2BWP30P140 U17 ( .I(i_valid[1]), .ZN(n52) );
  INVD2BWP30P140 U18 ( .I(i_cmd[0]), .ZN(n9) );
  INR2D2BWP30P140 U19 ( .A1(i_valid[0]), .B1(n51), .ZN(n4) );
  CKND2D2BWP30P140 U20 ( .A1(n4), .A2(n9), .ZN(n3) );
  INVD2BWP30P140 U21 ( .I(n27), .ZN(n26) );
  INVD1BWP30P140 U22 ( .I(n4), .ZN(n7) );
  INVD1BWP30P140 U23 ( .I(n51), .ZN(n5) );
  AN3D4BWP30P140 U24 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n5), .Z(n89) );
  OAI21D1BWP30P140 U25 ( .A1(n7), .A2(i_cmd[1]), .B(n6), .ZN(N354) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[19]), .ZN(n81) );
  INVD2BWP30P140 U27 ( .I(i_valid[0]), .ZN(n8) );
  NR2D1BWP30P140 U28 ( .A1(n51), .A2(n9), .ZN(n10) );
  INVD2BWP30P140 U29 ( .I(n12), .ZN(n14) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[51]), .ZN(n13) );
  OAI22D1BWP30P140 U31 ( .A1(n26), .A2(n81), .B1(n49), .B2(n13), .ZN(N306) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[52]), .ZN(n15) );
  OAI22D1BWP30P140 U34 ( .A1(n26), .A2(n80), .B1(n47), .B2(n15), .ZN(N307) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[21]), .ZN(n78) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[53]), .ZN(n16) );
  OAI22D1BWP30P140 U37 ( .A1(n26), .A2(n78), .B1(n47), .B2(n16), .ZN(N308) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[23]), .ZN(n76) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[55]), .ZN(n17) );
  OAI22D1BWP30P140 U40 ( .A1(n26), .A2(n76), .B1(n47), .B2(n17), .ZN(N310) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[25]), .ZN(n67) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[57]), .ZN(n18) );
  OAI22D1BWP30P140 U43 ( .A1(n26), .A2(n67), .B1(n47), .B2(n18), .ZN(N312) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[27]), .ZN(n66) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[59]), .ZN(n19) );
  OAI22D1BWP30P140 U46 ( .A1(n26), .A2(n66), .B1(n47), .B2(n19), .ZN(N314) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[29]), .ZN(n65) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[61]), .ZN(n20) );
  OAI22D1BWP30P140 U49 ( .A1(n26), .A2(n65), .B1(n47), .B2(n20), .ZN(N316) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[31]), .ZN(n64) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[63]), .ZN(n21) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[0]), .ZN(n63) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[32]), .ZN(n22) );
  OAI22D1BWP30P140 U54 ( .A1(n26), .A2(n63), .B1(n49), .B2(n22), .ZN(N287) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[33]), .ZN(n23) );
  OAI22D1BWP30P140 U57 ( .A1(n26), .A2(n59), .B1(n47), .B2(n23), .ZN(N288) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[34]), .ZN(n24) );
  OAI22D1BWP30P140 U60 ( .A1(n26), .A2(n62), .B1(n49), .B2(n24), .ZN(N289) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[3]), .ZN(n58) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[35]), .ZN(n25) );
  OAI22D1BWP30P140 U63 ( .A1(n26), .A2(n58), .B1(n47), .B2(n25), .ZN(N290) );
  INVD2BWP30P140 U64 ( .I(n27), .ZN(n50) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[39]), .ZN(n28) );
  OAI22D1BWP30P140 U67 ( .A1(n50), .A2(n56), .B1(n47), .B2(n28), .ZN(N294) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[8]), .ZN(n91) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[40]), .ZN(n29) );
  OAI22D1BWP30P140 U70 ( .A1(n50), .A2(n91), .B1(n49), .B2(n29), .ZN(N295) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[9]), .ZN(n71) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[41]), .ZN(n30) );
  OAI22D1BWP30P140 U73 ( .A1(n50), .A2(n71), .B1(n49), .B2(n30), .ZN(N296) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[42]), .ZN(n31) );
  OAI22D1BWP30P140 U76 ( .A1(n50), .A2(n88), .B1(n49), .B2(n31), .ZN(N297) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[11]), .ZN(n70) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[43]), .ZN(n32) );
  OAI22D1BWP30P140 U79 ( .A1(n50), .A2(n70), .B1(n49), .B2(n32), .ZN(N298) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[12]), .ZN(n87) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[44]), .ZN(n33) );
  OAI22D1BWP30P140 U82 ( .A1(n50), .A2(n87), .B1(n49), .B2(n33), .ZN(N299) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[13]), .ZN(n69) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[45]), .ZN(n34) );
  OAI22D1BWP30P140 U85 ( .A1(n50), .A2(n69), .B1(n49), .B2(n34), .ZN(N300) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[14]), .ZN(n86) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[46]), .ZN(n35) );
  OAI22D1BWP30P140 U88 ( .A1(n50), .A2(n86), .B1(n49), .B2(n35), .ZN(N301) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[15]), .ZN(n85) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[47]), .ZN(n36) );
  OAI22D1BWP30P140 U91 ( .A1(n50), .A2(n85), .B1(n49), .B2(n36), .ZN(N302) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[16]), .ZN(n84) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[48]), .ZN(n37) );
  OAI22D1BWP30P140 U94 ( .A1(n50), .A2(n84), .B1(n49), .B2(n37), .ZN(N303) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[17]), .ZN(n83) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[49]), .ZN(n38) );
  OAI22D1BWP30P140 U97 ( .A1(n50), .A2(n83), .B1(n49), .B2(n38), .ZN(N304) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[18]), .ZN(n82) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[50]), .ZN(n39) );
  OAI22D1BWP30P140 U100 ( .A1(n50), .A2(n82), .B1(n49), .B2(n39), .ZN(N305) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[22]), .ZN(n77) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[54]), .ZN(n40) );
  OAI22D1BWP30P140 U103 ( .A1(n50), .A2(n77), .B1(n47), .B2(n40), .ZN(N309) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[24]), .ZN(n75) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[56]), .ZN(n41) );
  OAI22D1BWP30P140 U106 ( .A1(n50), .A2(n75), .B1(n47), .B2(n41), .ZN(N311) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[26]), .ZN(n74) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[58]), .ZN(n42) );
  OAI22D1BWP30P140 U109 ( .A1(n50), .A2(n74), .B1(n47), .B2(n42), .ZN(N313) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[28]), .ZN(n73) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[60]), .ZN(n43) );
  OAI22D1BWP30P140 U112 ( .A1(n50), .A2(n73), .B1(n47), .B2(n43), .ZN(N315) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[30]), .ZN(n72) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[62]), .ZN(n44) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[36]), .ZN(n45) );
  OAI22D1BWP30P140 U117 ( .A1(n50), .A2(n61), .B1(n49), .B2(n45), .ZN(N291) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[5]), .ZN(n57) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[37]), .ZN(n46) );
  OAI22D1BWP30P140 U120 ( .A1(n50), .A2(n57), .B1(n47), .B2(n46), .ZN(N292) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[6]), .ZN(n60) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[38]), .ZN(n48) );
  OAI22D1BWP30P140 U123 ( .A1(n50), .A2(n60), .B1(n49), .B2(n48), .ZN(N293) );
  NR2D1BWP30P140 U124 ( .A1(n51), .A2(i_cmd[1]), .ZN(n54) );
  MUX2NUD1BWP30P140 U125 ( .I0(n8), .I1(n52), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U126 ( .A1(n54), .A2(n53), .ZN(n55) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n79), .B1(i_data_bus[39]), .B2(n89), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n79), .B1(i_data_bus[37]), .B2(n89), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n79), .B1(i_data_bus[35]), .B2(n89), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n79), .B1(i_data_bus[33]), .B2(n89), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n79), .B1(i_data_bus[38]), .B2(n89), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n79), .B1(i_data_bus[36]), .B2(n89), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n79), .B1(i_data_bus[34]), .B2(n89), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n79), .B1(i_data_bus[32]), .B2(n89), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n79), .B1(i_data_bus[63]), .B2(n89), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n79), .B1(i_data_bus[61]), .B2(n89), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n79), .B1(i_data_bus[59]), .B2(n89), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n79), .B1(i_data_bus[57]), .B2(n89), 
        .ZN(N344) );
  INVD2BWP30P140 U139 ( .I(n68), .ZN(n90) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n90), .B1(i_data_bus[45]), .B2(n89), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n90), .B1(i_data_bus[43]), .B2(n89), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n90), .B1(i_data_bus[41]), .B2(n89), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n79), .B1(i_data_bus[62]), .B2(n89), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n79), .B1(i_data_bus[60]), .B2(n89), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n79), .B1(i_data_bus[58]), .B2(n89), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n79), .B1(i_data_bus[56]), .B2(n89), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n79), .B1(i_data_bus[55]), .B2(n89), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n79), .B1(i_data_bus[54]), .B2(n89), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n79), .B1(i_data_bus[53]), .B2(n89), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n79), .B1(i_data_bus[52]), .B2(n89), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n90), .B1(i_data_bus[51]), .B2(n89), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n90), .B1(i_data_bus[50]), .B2(n89), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n90), .B1(i_data_bus[49]), .B2(n89), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n90), .B1(i_data_bus[48]), .B2(n89), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n90), .B1(i_data_bus[47]), .B2(n89), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n90), .B1(i_data_bus[46]), .B2(n89), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n90), .B1(i_data_bus[44]), .B2(n89), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n90), .B1(i_data_bus[42]), .B2(n89), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n91), .A2(n90), .B1(i_data_bus[40]), .B2(n89), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_2 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91;

  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  ND2OPTIBD1BWP30P140 U3 ( .A1(n3), .A2(n8), .ZN(n2) );
  INVD3BWP30P140 U4 ( .I(n68), .ZN(n79) );
  INVD1BWP30P140 U5 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U6 ( .I(i_valid[0]), .ZN(n7) );
  INVD1BWP30P140 U7 ( .I(n89), .ZN(n5) );
  INVD1BWP30P140 U8 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U9 ( .A1(n1), .A2(i_en), .ZN(n50) );
  INVD2BWP30P140 U10 ( .I(i_valid[1]), .ZN(n51) );
  INVD2BWP30P140 U11 ( .I(i_cmd[0]), .ZN(n8) );
  INR2D2BWP30P140 U12 ( .A1(i_valid[0]), .B1(n50), .ZN(n3) );
  INVD2BWP30P140 U13 ( .I(n2), .ZN(n26) );
  INVD2BWP30P140 U14 ( .I(n26), .ZN(n25) );
  OAI31D1BWP30P140 U15 ( .A1(n50), .A2(n51), .A3(n8), .B(n25), .ZN(N353) );
  INVD1BWP30P140 U16 ( .I(n3), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n50), .ZN(n4) );
  AN3D4BWP30P140 U18 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n4), .Z(n89) );
  OAI21D1BWP30P140 U19 ( .A1(n6), .A2(i_cmd[1]), .B(n5), .ZN(N354) );
  INVD1BWP30P140 U20 ( .I(i_data_bus[19]), .ZN(n81) );
  MUX2NOPTD2BWP30P140 U21 ( .I0(n7), .I1(n51), .S(i_cmd[1]), .ZN(n10) );
  NR2D1BWP30P140 U22 ( .A1(n50), .A2(n8), .ZN(n9) );
  CKND2D2BWP30P140 U23 ( .A1(n10), .A2(n9), .ZN(n11) );
  INVD2BWP30P140 U24 ( .I(n11), .ZN(n13) );
  INVD2BWP30P140 U25 ( .I(n13), .ZN(n46) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[51]), .ZN(n12) );
  OAI22D1BWP30P140 U27 ( .A1(n25), .A2(n81), .B1(n46), .B2(n12), .ZN(N306) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD2BWP30P140 U29 ( .I(n13), .ZN(n48) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[52]), .ZN(n14) );
  OAI22D1BWP30P140 U31 ( .A1(n25), .A2(n80), .B1(n48), .B2(n14), .ZN(N307) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[21]), .ZN(n78) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[53]), .ZN(n15) );
  OAI22D1BWP30P140 U34 ( .A1(n25), .A2(n78), .B1(n48), .B2(n15), .ZN(N308) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[23]), .ZN(n76) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[55]), .ZN(n16) );
  OAI22D1BWP30P140 U37 ( .A1(n25), .A2(n76), .B1(n48), .B2(n16), .ZN(N310) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[25]), .ZN(n67) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[57]), .ZN(n17) );
  OAI22D1BWP30P140 U40 ( .A1(n25), .A2(n67), .B1(n48), .B2(n17), .ZN(N312) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[27]), .ZN(n66) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[59]), .ZN(n18) );
  OAI22D1BWP30P140 U43 ( .A1(n25), .A2(n66), .B1(n48), .B2(n18), .ZN(N314) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[29]), .ZN(n65) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[61]), .ZN(n19) );
  OAI22D1BWP30P140 U46 ( .A1(n25), .A2(n65), .B1(n48), .B2(n19), .ZN(N316) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[31]), .ZN(n64) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[63]), .ZN(n20) );
  OAI22D1BWP30P140 U49 ( .A1(n25), .A2(n64), .B1(n48), .B2(n20), .ZN(N318) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[0]), .ZN(n63) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[32]), .ZN(n21) );
  OAI22D1BWP30P140 U52 ( .A1(n25), .A2(n63), .B1(n46), .B2(n21), .ZN(N287) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[33]), .ZN(n22) );
  OAI22D1BWP30P140 U55 ( .A1(n25), .A2(n58), .B1(n48), .B2(n22), .ZN(N288) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[34]), .ZN(n23) );
  OAI22D1BWP30P140 U58 ( .A1(n25), .A2(n62), .B1(n46), .B2(n23), .ZN(N289) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[3]), .ZN(n59) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[35]), .ZN(n24) );
  OAI22D1BWP30P140 U61 ( .A1(n25), .A2(n59), .B1(n48), .B2(n24), .ZN(N290) );
  INVD2BWP30P140 U62 ( .I(n26), .ZN(n49) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[8]), .ZN(n91) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[40]), .ZN(n27) );
  OAI22D1BWP30P140 U65 ( .A1(n49), .A2(n91), .B1(n46), .B2(n27), .ZN(N295) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[9]), .ZN(n71) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[41]), .ZN(n28) );
  OAI22D1BWP30P140 U68 ( .A1(n49), .A2(n71), .B1(n46), .B2(n28), .ZN(N296) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[42]), .ZN(n29) );
  OAI22D1BWP30P140 U71 ( .A1(n49), .A2(n88), .B1(n46), .B2(n29), .ZN(N297) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[11]), .ZN(n70) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[43]), .ZN(n30) );
  OAI22D1BWP30P140 U74 ( .A1(n49), .A2(n70), .B1(n46), .B2(n30), .ZN(N298) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[12]), .ZN(n87) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[44]), .ZN(n31) );
  OAI22D1BWP30P140 U77 ( .A1(n49), .A2(n87), .B1(n46), .B2(n31), .ZN(N299) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[13]), .ZN(n69) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[45]), .ZN(n32) );
  OAI22D1BWP30P140 U80 ( .A1(n49), .A2(n69), .B1(n46), .B2(n32), .ZN(N300) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[14]), .ZN(n86) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[46]), .ZN(n33) );
  OAI22D1BWP30P140 U83 ( .A1(n49), .A2(n86), .B1(n46), .B2(n33), .ZN(N301) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[15]), .ZN(n85) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[47]), .ZN(n34) );
  OAI22D1BWP30P140 U86 ( .A1(n49), .A2(n85), .B1(n46), .B2(n34), .ZN(N302) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[16]), .ZN(n84) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[48]), .ZN(n35) );
  OAI22D1BWP30P140 U89 ( .A1(n49), .A2(n84), .B1(n46), .B2(n35), .ZN(N303) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[17]), .ZN(n83) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[49]), .ZN(n36) );
  OAI22D1BWP30P140 U92 ( .A1(n49), .A2(n83), .B1(n46), .B2(n36), .ZN(N304) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[18]), .ZN(n82) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[50]), .ZN(n37) );
  OAI22D1BWP30P140 U95 ( .A1(n49), .A2(n82), .B1(n46), .B2(n37), .ZN(N305) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[22]), .ZN(n77) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[54]), .ZN(n38) );
  OAI22D1BWP30P140 U98 ( .A1(n49), .A2(n77), .B1(n48), .B2(n38), .ZN(N309) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[24]), .ZN(n75) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[56]), .ZN(n39) );
  OAI22D1BWP30P140 U101 ( .A1(n49), .A2(n75), .B1(n48), .B2(n39), .ZN(N311) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[26]), .ZN(n74) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[58]), .ZN(n40) );
  OAI22D1BWP30P140 U104 ( .A1(n49), .A2(n74), .B1(n48), .B2(n40), .ZN(N313) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[28]), .ZN(n73) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[60]), .ZN(n41) );
  OAI22D1BWP30P140 U107 ( .A1(n49), .A2(n73), .B1(n48), .B2(n41), .ZN(N315) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[30]), .ZN(n72) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[62]), .ZN(n42) );
  OAI22D1BWP30P140 U110 ( .A1(n49), .A2(n72), .B1(n48), .B2(n42), .ZN(N317) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[36]), .ZN(n43) );
  OAI22D1BWP30P140 U113 ( .A1(n49), .A2(n61), .B1(n46), .B2(n43), .ZN(N291) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[5]), .ZN(n57) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[37]), .ZN(n44) );
  OAI22D1BWP30P140 U116 ( .A1(n49), .A2(n57), .B1(n48), .B2(n44), .ZN(N292) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[6]), .ZN(n60) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[38]), .ZN(n45) );
  OAI22D1BWP30P140 U119 ( .A1(n49), .A2(n60), .B1(n46), .B2(n45), .ZN(N293) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[39]), .ZN(n47) );
  OAI22D1BWP30P140 U122 ( .A1(n49), .A2(n56), .B1(n48), .B2(n47), .ZN(N294) );
  NR2D1BWP30P140 U123 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n68) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n79), .B1(i_data_bus[39]), .B2(n89), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n79), .B1(i_data_bus[37]), .B2(n89), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n79), .B1(i_data_bus[33]), .B2(n89), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n79), .B1(i_data_bus[35]), .B2(n89), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n79), .B1(i_data_bus[38]), .B2(n89), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n79), .B1(i_data_bus[36]), .B2(n89), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n79), .B1(i_data_bus[34]), .B2(n89), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n79), .B1(i_data_bus[32]), .B2(n89), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n79), .B1(i_data_bus[63]), .B2(n89), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n79), .B1(i_data_bus[61]), .B2(n89), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n79), .B1(i_data_bus[59]), .B2(n89), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n79), .B1(i_data_bus[57]), .B2(n89), 
        .ZN(N344) );
  INVD2BWP30P140 U139 ( .I(n68), .ZN(n90) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n90), .B1(i_data_bus[45]), .B2(n89), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n90), .B1(i_data_bus[43]), .B2(n89), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n90), .B1(i_data_bus[41]), .B2(n89), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n79), .B1(i_data_bus[62]), .B2(n89), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n79), .B1(i_data_bus[60]), .B2(n89), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n79), .B1(i_data_bus[58]), .B2(n89), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n79), .B1(i_data_bus[56]), .B2(n89), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n79), .B1(i_data_bus[55]), .B2(n89), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n79), .B1(i_data_bus[54]), .B2(n89), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n79), .B1(i_data_bus[53]), .B2(n89), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n79), .B1(i_data_bus[52]), .B2(n89), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n90), .B1(i_data_bus[51]), .B2(n89), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n90), .B1(i_data_bus[50]), .B2(n89), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n90), .B1(i_data_bus[49]), .B2(n89), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n90), .B1(i_data_bus[48]), .B2(n89), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n90), .B1(i_data_bus[47]), .B2(n89), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n90), .B1(i_data_bus[46]), .B2(n89), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n90), .B1(i_data_bus[44]), .B2(n89), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n90), .B1(i_data_bus[42]), .B2(n89), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n91), .A2(n90), .B1(i_data_bus[40]), .B2(n89), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_3 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91;

  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  ND2OPTIBD1BWP30P140 U3 ( .A1(n3), .A2(n8), .ZN(n2) );
  INVD3BWP30P140 U4 ( .I(n68), .ZN(n79) );
  INVD1BWP30P140 U5 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U6 ( .I(i_valid[0]), .ZN(n7) );
  INVD1BWP30P140 U7 ( .I(n89), .ZN(n5) );
  INVD1BWP30P140 U8 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U9 ( .A1(n1), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U10 ( .I(i_valid[1]), .ZN(n51) );
  INVD2BWP30P140 U11 ( .I(i_cmd[0]), .ZN(n8) );
  INR2D2BWP30P140 U12 ( .A1(i_valid[0]), .B1(n50), .ZN(n3) );
  INVD2BWP30P140 U13 ( .I(n2), .ZN(n26) );
  INVD2BWP30P140 U14 ( .I(n26), .ZN(n25) );
  OAI31D1BWP30P140 U15 ( .A1(n50), .A2(n51), .A3(n8), .B(n25), .ZN(N353) );
  INVD1BWP30P140 U16 ( .I(n3), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n50), .ZN(n4) );
  AN3D4BWP30P140 U18 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n4), .Z(n89) );
  OAI21D1BWP30P140 U19 ( .A1(n6), .A2(i_cmd[1]), .B(n5), .ZN(N354) );
  INVD1BWP30P140 U20 ( .I(i_data_bus[19]), .ZN(n81) );
  MUX2NOPTD2BWP30P140 U21 ( .I0(n7), .I1(n51), .S(i_cmd[1]), .ZN(n10) );
  NR2D1BWP30P140 U22 ( .A1(n50), .A2(n8), .ZN(n9) );
  CKND2D2BWP30P140 U23 ( .A1(n10), .A2(n9), .ZN(n11) );
  INVD2BWP30P140 U24 ( .I(n11), .ZN(n13) );
  INVD2BWP30P140 U25 ( .I(n13), .ZN(n46) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[51]), .ZN(n12) );
  OAI22D1BWP30P140 U27 ( .A1(n25), .A2(n81), .B1(n46), .B2(n12), .ZN(N306) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD2BWP30P140 U29 ( .I(n13), .ZN(n48) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[52]), .ZN(n14) );
  OAI22D1BWP30P140 U31 ( .A1(n25), .A2(n80), .B1(n48), .B2(n14), .ZN(N307) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[21]), .ZN(n78) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[53]), .ZN(n15) );
  OAI22D1BWP30P140 U34 ( .A1(n25), .A2(n78), .B1(n48), .B2(n15), .ZN(N308) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[23]), .ZN(n76) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[55]), .ZN(n16) );
  OAI22D1BWP30P140 U37 ( .A1(n25), .A2(n76), .B1(n48), .B2(n16), .ZN(N310) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[25]), .ZN(n67) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[57]), .ZN(n17) );
  OAI22D1BWP30P140 U40 ( .A1(n25), .A2(n67), .B1(n48), .B2(n17), .ZN(N312) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[27]), .ZN(n66) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[59]), .ZN(n18) );
  OAI22D1BWP30P140 U43 ( .A1(n25), .A2(n66), .B1(n48), .B2(n18), .ZN(N314) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[29]), .ZN(n65) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[61]), .ZN(n19) );
  OAI22D1BWP30P140 U46 ( .A1(n25), .A2(n65), .B1(n48), .B2(n19), .ZN(N316) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[31]), .ZN(n64) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[63]), .ZN(n20) );
  OAI22D1BWP30P140 U49 ( .A1(n25), .A2(n64), .B1(n48), .B2(n20), .ZN(N318) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[0]), .ZN(n63) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[32]), .ZN(n21) );
  OAI22D1BWP30P140 U52 ( .A1(n25), .A2(n63), .B1(n46), .B2(n21), .ZN(N287) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[33]), .ZN(n22) );
  OAI22D1BWP30P140 U55 ( .A1(n25), .A2(n59), .B1(n48), .B2(n22), .ZN(N288) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[34]), .ZN(n23) );
  OAI22D1BWP30P140 U58 ( .A1(n25), .A2(n62), .B1(n46), .B2(n23), .ZN(N289) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[3]), .ZN(n58) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[35]), .ZN(n24) );
  OAI22D1BWP30P140 U61 ( .A1(n25), .A2(n58), .B1(n48), .B2(n24), .ZN(N290) );
  INVD2BWP30P140 U62 ( .I(n26), .ZN(n49) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[8]), .ZN(n91) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[40]), .ZN(n27) );
  OAI22D1BWP30P140 U65 ( .A1(n49), .A2(n91), .B1(n46), .B2(n27), .ZN(N295) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[9]), .ZN(n71) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[41]), .ZN(n28) );
  OAI22D1BWP30P140 U68 ( .A1(n49), .A2(n71), .B1(n46), .B2(n28), .ZN(N296) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[42]), .ZN(n29) );
  OAI22D1BWP30P140 U71 ( .A1(n49), .A2(n88), .B1(n46), .B2(n29), .ZN(N297) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[11]), .ZN(n70) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[43]), .ZN(n30) );
  OAI22D1BWP30P140 U74 ( .A1(n49), .A2(n70), .B1(n46), .B2(n30), .ZN(N298) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[12]), .ZN(n87) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[44]), .ZN(n31) );
  OAI22D1BWP30P140 U77 ( .A1(n49), .A2(n87), .B1(n46), .B2(n31), .ZN(N299) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[13]), .ZN(n69) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[45]), .ZN(n32) );
  OAI22D1BWP30P140 U80 ( .A1(n49), .A2(n69), .B1(n46), .B2(n32), .ZN(N300) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[14]), .ZN(n86) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[46]), .ZN(n33) );
  OAI22D1BWP30P140 U83 ( .A1(n49), .A2(n86), .B1(n46), .B2(n33), .ZN(N301) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[15]), .ZN(n85) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[47]), .ZN(n34) );
  OAI22D1BWP30P140 U86 ( .A1(n49), .A2(n85), .B1(n46), .B2(n34), .ZN(N302) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[16]), .ZN(n84) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[48]), .ZN(n35) );
  OAI22D1BWP30P140 U89 ( .A1(n49), .A2(n84), .B1(n46), .B2(n35), .ZN(N303) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[17]), .ZN(n83) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[49]), .ZN(n36) );
  OAI22D1BWP30P140 U92 ( .A1(n49), .A2(n83), .B1(n46), .B2(n36), .ZN(N304) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[18]), .ZN(n82) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[50]), .ZN(n37) );
  OAI22D1BWP30P140 U95 ( .A1(n49), .A2(n82), .B1(n46), .B2(n37), .ZN(N305) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[22]), .ZN(n77) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[54]), .ZN(n38) );
  OAI22D1BWP30P140 U98 ( .A1(n49), .A2(n77), .B1(n48), .B2(n38), .ZN(N309) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[24]), .ZN(n75) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[56]), .ZN(n39) );
  OAI22D1BWP30P140 U101 ( .A1(n49), .A2(n75), .B1(n48), .B2(n39), .ZN(N311) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[26]), .ZN(n74) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[58]), .ZN(n40) );
  OAI22D1BWP30P140 U104 ( .A1(n49), .A2(n74), .B1(n48), .B2(n40), .ZN(N313) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[28]), .ZN(n73) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[60]), .ZN(n41) );
  OAI22D1BWP30P140 U107 ( .A1(n49), .A2(n73), .B1(n48), .B2(n41), .ZN(N315) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[30]), .ZN(n72) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[62]), .ZN(n42) );
  OAI22D1BWP30P140 U110 ( .A1(n49), .A2(n72), .B1(n48), .B2(n42), .ZN(N317) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[36]), .ZN(n43) );
  OAI22D1BWP30P140 U113 ( .A1(n49), .A2(n61), .B1(n46), .B2(n43), .ZN(N291) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[5]), .ZN(n57) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[37]), .ZN(n44) );
  OAI22D1BWP30P140 U116 ( .A1(n49), .A2(n57), .B1(n48), .B2(n44), .ZN(N292) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[6]), .ZN(n60) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[38]), .ZN(n45) );
  OAI22D1BWP30P140 U119 ( .A1(n49), .A2(n60), .B1(n46), .B2(n45), .ZN(N293) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[39]), .ZN(n47) );
  OAI22D1BWP30P140 U122 ( .A1(n49), .A2(n56), .B1(n48), .B2(n47), .ZN(N294) );
  NR2D1BWP30P140 U123 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n68) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n79), .B1(i_data_bus[39]), .B2(n89), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n79), .B1(i_data_bus[37]), .B2(n89), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n79), .B1(i_data_bus[35]), .B2(n89), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n79), .B1(i_data_bus[33]), .B2(n89), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n79), .B1(i_data_bus[38]), .B2(n89), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n79), .B1(i_data_bus[36]), .B2(n89), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n79), .B1(i_data_bus[34]), .B2(n89), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n79), .B1(i_data_bus[32]), .B2(n89), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n79), .B1(i_data_bus[63]), .B2(n89), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n79), .B1(i_data_bus[61]), .B2(n89), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n79), .B1(i_data_bus[59]), .B2(n89), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n79), .B1(i_data_bus[57]), .B2(n89), 
        .ZN(N344) );
  INVD2BWP30P140 U139 ( .I(n68), .ZN(n90) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n90), .B1(i_data_bus[45]), .B2(n89), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n90), .B1(i_data_bus[43]), .B2(n89), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n90), .B1(i_data_bus[41]), .B2(n89), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n79), .B1(i_data_bus[62]), .B2(n89), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n79), .B1(i_data_bus[60]), .B2(n89), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n79), .B1(i_data_bus[58]), .B2(n89), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n79), .B1(i_data_bus[56]), .B2(n89), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n79), .B1(i_data_bus[55]), .B2(n89), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n79), .B1(i_data_bus[54]), .B2(n89), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n79), .B1(i_data_bus[53]), .B2(n89), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n79), .B1(i_data_bus[52]), .B2(n89), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n90), .B1(i_data_bus[51]), .B2(n89), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n90), .B1(i_data_bus[50]), .B2(n89), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n90), .B1(i_data_bus[49]), .B2(n89), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n90), .B1(i_data_bus[48]), .B2(n89), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n90), .B1(i_data_bus[47]), .B2(n89), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n90), .B1(i_data_bus[46]), .B2(n89), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n90), .B1(i_data_bus[44]), .B2(n89), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n90), .B1(i_data_bus[42]), .B2(n89), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n91), .A2(n90), .B1(i_data_bus[40]), .B2(n89), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_4 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91;

  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  ND2OPTIBD1BWP30P140 U3 ( .A1(n3), .A2(n8), .ZN(n2) );
  INVD3BWP30P140 U4 ( .I(n69), .ZN(n90) );
  INVD1BWP30P140 U5 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U6 ( .I(i_valid[0]), .ZN(n7) );
  INVD1BWP30P140 U7 ( .I(n89), .ZN(n5) );
  INVD1BWP30P140 U8 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U9 ( .A1(n1), .A2(i_en), .ZN(n50) );
  INVD2BWP30P140 U10 ( .I(i_valid[1]), .ZN(n51) );
  INVD2BWP30P140 U11 ( .I(i_cmd[0]), .ZN(n8) );
  INR2D2BWP30P140 U12 ( .A1(i_valid[0]), .B1(n50), .ZN(n3) );
  INVD2BWP30P140 U13 ( .I(n2), .ZN(n26) );
  INVD2BWP30P140 U14 ( .I(n26), .ZN(n25) );
  OAI31D1BWP30P140 U15 ( .A1(n50), .A2(n51), .A3(n8), .B(n25), .ZN(N353) );
  INVD1BWP30P140 U16 ( .I(n3), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n50), .ZN(n4) );
  AN3D4BWP30P140 U18 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n4), .Z(n89) );
  OAI21D1BWP30P140 U19 ( .A1(n6), .A2(i_cmd[1]), .B(n5), .ZN(N354) );
  INVD1BWP30P140 U20 ( .I(i_data_bus[21]), .ZN(n83) );
  MUX2NOPTD2BWP30P140 U21 ( .I0(n7), .I1(n51), .S(i_cmd[1]), .ZN(n10) );
  NR2D1BWP30P140 U22 ( .A1(n50), .A2(n8), .ZN(n9) );
  CKND2D2BWP30P140 U23 ( .A1(n10), .A2(n9), .ZN(n11) );
  INVD2BWP30P140 U24 ( .I(n11), .ZN(n14) );
  INVD2BWP30P140 U25 ( .I(n14), .ZN(n48) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[53]), .ZN(n12) );
  OAI22D1BWP30P140 U27 ( .A1(n25), .A2(n83), .B1(n48), .B2(n12), .ZN(N308) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[20]), .ZN(n85) );
  INVD1BWP30P140 U29 ( .I(i_data_bus[52]), .ZN(n13) );
  OAI22D1BWP30P140 U30 ( .A1(n25), .A2(n85), .B1(n48), .B2(n13), .ZN(N307) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[19]), .ZN(n86) );
  INVD2BWP30P140 U32 ( .I(n14), .ZN(n46) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[51]), .ZN(n15) );
  OAI22D1BWP30P140 U34 ( .A1(n25), .A2(n86), .B1(n46), .B2(n15), .ZN(N306) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[3]), .ZN(n59) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[35]), .ZN(n16) );
  OAI22D1BWP30P140 U37 ( .A1(n25), .A2(n59), .B1(n48), .B2(n16), .ZN(N290) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[2]), .ZN(n61) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[34]), .ZN(n17) );
  OAI22D1BWP30P140 U40 ( .A1(n25), .A2(n61), .B1(n46), .B2(n17), .ZN(N289) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[1]), .ZN(n56) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[33]), .ZN(n18) );
  OAI22D1BWP30P140 U43 ( .A1(n25), .A2(n56), .B1(n48), .B2(n18), .ZN(N288) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[0]), .ZN(n60) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[32]), .ZN(n19) );
  OAI22D1BWP30P140 U46 ( .A1(n25), .A2(n60), .B1(n46), .B2(n19), .ZN(N287) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[31]), .ZN(n70) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[63]), .ZN(n20) );
  OAI22D1BWP30P140 U49 ( .A1(n25), .A2(n70), .B1(n48), .B2(n20), .ZN(N318) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[29]), .ZN(n71) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[61]), .ZN(n21) );
  OAI22D1BWP30P140 U52 ( .A1(n25), .A2(n71), .B1(n48), .B2(n21), .ZN(N316) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[27]), .ZN(n72) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[59]), .ZN(n22) );
  OAI22D1BWP30P140 U55 ( .A1(n25), .A2(n72), .B1(n48), .B2(n22), .ZN(N314) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[25]), .ZN(n73) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[57]), .ZN(n23) );
  OAI22D1BWP30P140 U58 ( .A1(n25), .A2(n73), .B1(n48), .B2(n23), .ZN(N312) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[23]), .ZN(n81) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[55]), .ZN(n24) );
  OAI22D1BWP30P140 U61 ( .A1(n25), .A2(n81), .B1(n48), .B2(n24), .ZN(N310) );
  INVD2BWP30P140 U62 ( .I(n26), .ZN(n49) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[8]), .ZN(n67) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[40]), .ZN(n27) );
  OAI22D1BWP30P140 U65 ( .A1(n49), .A2(n67), .B1(n46), .B2(n27), .ZN(N295) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[9]), .ZN(n76) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[41]), .ZN(n28) );
  OAI22D1BWP30P140 U68 ( .A1(n49), .A2(n76), .B1(n46), .B2(n28), .ZN(N296) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[10]), .ZN(n66) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[42]), .ZN(n29) );
  OAI22D1BWP30P140 U71 ( .A1(n49), .A2(n66), .B1(n46), .B2(n29), .ZN(N297) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[11]), .ZN(n75) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[43]), .ZN(n30) );
  OAI22D1BWP30P140 U74 ( .A1(n49), .A2(n75), .B1(n46), .B2(n30), .ZN(N298) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[12]), .ZN(n65) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[44]), .ZN(n31) );
  OAI22D1BWP30P140 U77 ( .A1(n49), .A2(n65), .B1(n46), .B2(n31), .ZN(N299) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[13]), .ZN(n74) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[45]), .ZN(n32) );
  OAI22D1BWP30P140 U80 ( .A1(n49), .A2(n74), .B1(n46), .B2(n32), .ZN(N300) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[14]), .ZN(n64) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[46]), .ZN(n33) );
  OAI22D1BWP30P140 U83 ( .A1(n49), .A2(n64), .B1(n46), .B2(n33), .ZN(N301) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[15]), .ZN(n68) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[47]), .ZN(n34) );
  OAI22D1BWP30P140 U86 ( .A1(n49), .A2(n68), .B1(n46), .B2(n34), .ZN(N302) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[16]), .ZN(n91) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[48]), .ZN(n35) );
  OAI22D1BWP30P140 U89 ( .A1(n49), .A2(n91), .B1(n46), .B2(n35), .ZN(N303) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[17]), .ZN(n88) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[49]), .ZN(n36) );
  OAI22D1BWP30P140 U92 ( .A1(n49), .A2(n88), .B1(n46), .B2(n36), .ZN(N304) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[18]), .ZN(n87) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[50]), .ZN(n37) );
  OAI22D1BWP30P140 U95 ( .A1(n49), .A2(n87), .B1(n46), .B2(n37), .ZN(N305) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[22]), .ZN(n82) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[54]), .ZN(n38) );
  OAI22D1BWP30P140 U98 ( .A1(n49), .A2(n82), .B1(n48), .B2(n38), .ZN(N309) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[24]), .ZN(n80) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[56]), .ZN(n39) );
  OAI22D1BWP30P140 U101 ( .A1(n49), .A2(n80), .B1(n48), .B2(n39), .ZN(N311) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[26]), .ZN(n79) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[58]), .ZN(n40) );
  OAI22D1BWP30P140 U104 ( .A1(n49), .A2(n79), .B1(n48), .B2(n40), .ZN(N313) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[28]), .ZN(n78) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[60]), .ZN(n41) );
  OAI22D1BWP30P140 U107 ( .A1(n49), .A2(n78), .B1(n48), .B2(n41), .ZN(N315) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[30]), .ZN(n77) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[62]), .ZN(n42) );
  OAI22D1BWP30P140 U110 ( .A1(n49), .A2(n77), .B1(n48), .B2(n42), .ZN(N317) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[36]), .ZN(n43) );
  OAI22D1BWP30P140 U113 ( .A1(n49), .A2(n62), .B1(n46), .B2(n43), .ZN(N291) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[5]), .ZN(n58) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[37]), .ZN(n44) );
  OAI22D1BWP30P140 U116 ( .A1(n49), .A2(n58), .B1(n48), .B2(n44), .ZN(N292) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[38]), .ZN(n45) );
  OAI22D1BWP30P140 U119 ( .A1(n49), .A2(n63), .B1(n46), .B2(n45), .ZN(N293) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[39]), .ZN(n47) );
  OAI22D1BWP30P140 U122 ( .A1(n49), .A2(n57), .B1(n48), .B2(n47), .ZN(N294) );
  NR2D1BWP30P140 U123 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n69) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n90), .B1(i_data_bus[33]), .B2(n89), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n90), .B1(i_data_bus[39]), .B2(n89), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n90), .B1(i_data_bus[37]), .B2(n89), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n90), .B1(i_data_bus[35]), .B2(n89), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n90), .B1(i_data_bus[32]), .B2(n89), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n90), .B1(i_data_bus[34]), .B2(n89), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n90), .B1(i_data_bus[36]), .B2(n89), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n90), .B1(i_data_bus[38]), .B2(n89), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n90), .B1(i_data_bus[46]), .B2(n89), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n90), .B1(i_data_bus[44]), .B2(n89), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n90), .B1(i_data_bus[42]), .B2(n89), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n90), .B1(i_data_bus[40]), .B2(n89), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n90), .B1(i_data_bus[47]), .B2(n89), 
        .ZN(N334) );
  INVD2BWP30P140 U140 ( .I(n69), .ZN(n84) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n84), .B1(i_data_bus[63]), .B2(n89), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n84), .B1(i_data_bus[61]), .B2(n89), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n84), .B1(i_data_bus[59]), .B2(n89), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n84), .B1(i_data_bus[57]), .B2(n89), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n90), .B1(i_data_bus[45]), .B2(n89), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n90), .B1(i_data_bus[43]), .B2(n89), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n90), .B1(i_data_bus[41]), .B2(n89), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n84), .B1(i_data_bus[62]), .B2(n89), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n84), .B1(i_data_bus[60]), .B2(n89), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n84), .B1(i_data_bus[58]), .B2(n89), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n84), .B1(i_data_bus[56]), .B2(n89), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n84), .B1(i_data_bus[55]), .B2(n89), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n84), .B1(i_data_bus[54]), .B2(n89), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n84), .B1(i_data_bus[53]), .B2(n89), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n84), .B1(i_data_bus[52]), .B2(n89), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n90), .B1(i_data_bus[51]), .B2(n89), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n90), .B1(i_data_bus[50]), .B2(n89), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n90), .B1(i_data_bus[49]), .B2(n89), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U159 ( .A1(n91), .A2(n90), .B1(i_data_bus[48]), .B2(n89), 
        .ZN(N335) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_5 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91;

  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  ND2OPTIBD1BWP30P140 U3 ( .A1(n3), .A2(n8), .ZN(n2) );
  INVD3BWP30P140 U4 ( .I(n68), .ZN(n79) );
  INVD1BWP30P140 U5 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U6 ( .I(i_valid[0]), .ZN(n7) );
  INVD1BWP30P140 U7 ( .I(n89), .ZN(n5) );
  INVD1BWP30P140 U8 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U9 ( .A1(n1), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U10 ( .I(i_valid[1]), .ZN(n51) );
  INVD2BWP30P140 U11 ( .I(i_cmd[0]), .ZN(n8) );
  INR2D2BWP30P140 U12 ( .A1(i_valid[0]), .B1(n50), .ZN(n3) );
  INVD2BWP30P140 U13 ( .I(n2), .ZN(n26) );
  INVD2BWP30P140 U14 ( .I(n26), .ZN(n25) );
  OAI31D1BWP30P140 U15 ( .A1(n50), .A2(n51), .A3(n8), .B(n25), .ZN(N353) );
  INVD1BWP30P140 U16 ( .I(n3), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n50), .ZN(n4) );
  AN3D4BWP30P140 U18 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n4), .Z(n89) );
  OAI21D1BWP30P140 U19 ( .A1(n6), .A2(i_cmd[1]), .B(n5), .ZN(N354) );
  INVD1BWP30P140 U20 ( .I(i_data_bus[0]), .ZN(n56) );
  MUX2NOPTD2BWP30P140 U21 ( .I0(n7), .I1(n51), .S(i_cmd[1]), .ZN(n10) );
  NR2D1BWP30P140 U22 ( .A1(n50), .A2(n8), .ZN(n9) );
  CKND2D2BWP30P140 U23 ( .A1(n10), .A2(n9), .ZN(n11) );
  INVD2BWP30P140 U24 ( .I(n11), .ZN(n13) );
  INVD2BWP30P140 U25 ( .I(n13), .ZN(n46) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[32]), .ZN(n12) );
  OAI22D1BWP30P140 U27 ( .A1(n25), .A2(n56), .B1(n46), .B2(n12), .ZN(N287) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[27]), .ZN(n66) );
  INVD2BWP30P140 U29 ( .I(n13), .ZN(n48) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[59]), .ZN(n14) );
  OAI22D1BWP30P140 U31 ( .A1(n25), .A2(n66), .B1(n48), .B2(n14), .ZN(N314) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[29]), .ZN(n65) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[61]), .ZN(n15) );
  OAI22D1BWP30P140 U34 ( .A1(n25), .A2(n65), .B1(n48), .B2(n15), .ZN(N316) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[1]), .ZN(n60) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[33]), .ZN(n16) );
  OAI22D1BWP30P140 U37 ( .A1(n25), .A2(n60), .B1(n48), .B2(n16), .ZN(N288) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[2]), .ZN(n57) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[34]), .ZN(n17) );
  OAI22D1BWP30P140 U40 ( .A1(n25), .A2(n57), .B1(n46), .B2(n17), .ZN(N289) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[35]), .ZN(n18) );
  OAI22D1BWP30P140 U43 ( .A1(n25), .A2(n61), .B1(n48), .B2(n18), .ZN(N290) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[31]), .ZN(n64) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[63]), .ZN(n19) );
  OAI22D1BWP30P140 U46 ( .A1(n25), .A2(n64), .B1(n48), .B2(n19), .ZN(N318) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[25]), .ZN(n67) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[57]), .ZN(n20) );
  OAI22D1BWP30P140 U49 ( .A1(n25), .A2(n67), .B1(n48), .B2(n20), .ZN(N312) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[19]), .ZN(n81) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[51]), .ZN(n21) );
  OAI22D1BWP30P140 U52 ( .A1(n25), .A2(n81), .B1(n46), .B2(n21), .ZN(N306) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[52]), .ZN(n22) );
  OAI22D1BWP30P140 U55 ( .A1(n25), .A2(n80), .B1(n48), .B2(n22), .ZN(N307) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[21]), .ZN(n78) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[53]), .ZN(n23) );
  OAI22D1BWP30P140 U58 ( .A1(n25), .A2(n78), .B1(n48), .B2(n23), .ZN(N308) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[23]), .ZN(n76) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[55]), .ZN(n24) );
  OAI22D1BWP30P140 U61 ( .A1(n25), .A2(n76), .B1(n48), .B2(n24), .ZN(N310) );
  INVD2BWP30P140 U62 ( .I(n26), .ZN(n49) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[8]), .ZN(n91) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[40]), .ZN(n27) );
  OAI22D1BWP30P140 U65 ( .A1(n49), .A2(n91), .B1(n46), .B2(n27), .ZN(N295) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[9]), .ZN(n71) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[41]), .ZN(n28) );
  OAI22D1BWP30P140 U68 ( .A1(n49), .A2(n71), .B1(n46), .B2(n28), .ZN(N296) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[42]), .ZN(n29) );
  OAI22D1BWP30P140 U71 ( .A1(n49), .A2(n88), .B1(n46), .B2(n29), .ZN(N297) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[11]), .ZN(n70) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[43]), .ZN(n30) );
  OAI22D1BWP30P140 U74 ( .A1(n49), .A2(n70), .B1(n46), .B2(n30), .ZN(N298) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[12]), .ZN(n87) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[44]), .ZN(n31) );
  OAI22D1BWP30P140 U77 ( .A1(n49), .A2(n87), .B1(n46), .B2(n31), .ZN(N299) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[13]), .ZN(n69) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[45]), .ZN(n32) );
  OAI22D1BWP30P140 U80 ( .A1(n49), .A2(n69), .B1(n46), .B2(n32), .ZN(N300) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[14]), .ZN(n86) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[46]), .ZN(n33) );
  OAI22D1BWP30P140 U83 ( .A1(n49), .A2(n86), .B1(n46), .B2(n33), .ZN(N301) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[15]), .ZN(n85) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[47]), .ZN(n34) );
  OAI22D1BWP30P140 U86 ( .A1(n49), .A2(n85), .B1(n46), .B2(n34), .ZN(N302) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[16]), .ZN(n84) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[48]), .ZN(n35) );
  OAI22D1BWP30P140 U89 ( .A1(n49), .A2(n84), .B1(n46), .B2(n35), .ZN(N303) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[17]), .ZN(n83) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[49]), .ZN(n36) );
  OAI22D1BWP30P140 U92 ( .A1(n49), .A2(n83), .B1(n46), .B2(n36), .ZN(N304) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[18]), .ZN(n82) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[50]), .ZN(n37) );
  OAI22D1BWP30P140 U95 ( .A1(n49), .A2(n82), .B1(n46), .B2(n37), .ZN(N305) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[22]), .ZN(n77) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[54]), .ZN(n38) );
  OAI22D1BWP30P140 U98 ( .A1(n49), .A2(n77), .B1(n48), .B2(n38), .ZN(N309) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[24]), .ZN(n75) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[56]), .ZN(n39) );
  OAI22D1BWP30P140 U101 ( .A1(n49), .A2(n75), .B1(n48), .B2(n39), .ZN(N311) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[26]), .ZN(n74) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[58]), .ZN(n40) );
  OAI22D1BWP30P140 U104 ( .A1(n49), .A2(n74), .B1(n48), .B2(n40), .ZN(N313) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[28]), .ZN(n73) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[60]), .ZN(n41) );
  OAI22D1BWP30P140 U107 ( .A1(n49), .A2(n73), .B1(n48), .B2(n41), .ZN(N315) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[30]), .ZN(n72) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[62]), .ZN(n42) );
  OAI22D1BWP30P140 U110 ( .A1(n49), .A2(n72), .B1(n48), .B2(n42), .ZN(N317) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[4]), .ZN(n58) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[36]), .ZN(n43) );
  OAI22D1BWP30P140 U113 ( .A1(n49), .A2(n58), .B1(n46), .B2(n43), .ZN(N291) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[37]), .ZN(n44) );
  OAI22D1BWP30P140 U116 ( .A1(n49), .A2(n62), .B1(n48), .B2(n44), .ZN(N292) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[6]), .ZN(n59) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[38]), .ZN(n45) );
  OAI22D1BWP30P140 U119 ( .A1(n49), .A2(n59), .B1(n46), .B2(n45), .ZN(N293) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[7]), .ZN(n63) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[39]), .ZN(n47) );
  OAI22D1BWP30P140 U122 ( .A1(n49), .A2(n63), .B1(n48), .B2(n47), .ZN(N294) );
  NR2D1BWP30P140 U123 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n68) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n79), .B1(i_data_bus[32]), .B2(n89), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n79), .B1(i_data_bus[34]), .B2(n89), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n79), .B1(i_data_bus[36]), .B2(n89), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n79), .B1(i_data_bus[38]), .B2(n89), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n79), .B1(i_data_bus[33]), .B2(n89), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n79), .B1(i_data_bus[35]), .B2(n89), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n79), .B1(i_data_bus[37]), .B2(n89), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n79), .B1(i_data_bus[39]), .B2(n89), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n79), .B1(i_data_bus[63]), .B2(n89), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n79), .B1(i_data_bus[61]), .B2(n89), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n79), .B1(i_data_bus[59]), .B2(n89), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n79), .B1(i_data_bus[57]), .B2(n89), 
        .ZN(N344) );
  INVD2BWP30P140 U139 ( .I(n68), .ZN(n90) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n90), .B1(i_data_bus[45]), .B2(n89), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n90), .B1(i_data_bus[43]), .B2(n89), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n90), .B1(i_data_bus[41]), .B2(n89), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n79), .B1(i_data_bus[62]), .B2(n89), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n79), .B1(i_data_bus[60]), .B2(n89), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n79), .B1(i_data_bus[58]), .B2(n89), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n79), .B1(i_data_bus[56]), .B2(n89), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n79), .B1(i_data_bus[55]), .B2(n89), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n79), .B1(i_data_bus[54]), .B2(n89), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n79), .B1(i_data_bus[53]), .B2(n89), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n79), .B1(i_data_bus[52]), .B2(n89), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n90), .B1(i_data_bus[51]), .B2(n89), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n90), .B1(i_data_bus[50]), .B2(n89), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n90), .B1(i_data_bus[49]), .B2(n89), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n90), .B1(i_data_bus[48]), .B2(n89), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n90), .B1(i_data_bus[47]), .B2(n89), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n90), .B1(i_data_bus[46]), .B2(n89), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n90), .B1(i_data_bus[44]), .B2(n89), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n90), .B1(i_data_bus[42]), .B2(n89), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n91), .A2(n90), .B1(i_data_bus[40]), .B2(n89), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_6 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91;

  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  ND2OPTIBD1BWP30P140 U3 ( .A1(n3), .A2(n8), .ZN(n2) );
  INVD3BWP30P140 U4 ( .I(n69), .ZN(n90) );
  INVD1BWP30P140 U5 ( .I(i_valid[0]), .ZN(n52) );
  INVD1BWP30P140 U6 ( .I(i_valid[0]), .ZN(n7) );
  INVD1BWP30P140 U7 ( .I(n89), .ZN(n5) );
  INVD1BWP30P140 U8 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U9 ( .A1(n1), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U10 ( .I(i_valid[1]), .ZN(n51) );
  INVD2BWP30P140 U11 ( .I(i_cmd[0]), .ZN(n8) );
  INR2D2BWP30P140 U12 ( .A1(i_valid[0]), .B1(n50), .ZN(n3) );
  INVD2BWP30P140 U13 ( .I(n2), .ZN(n26) );
  INVD2BWP30P140 U14 ( .I(n26), .ZN(n25) );
  OAI31D1BWP30P140 U15 ( .A1(n50), .A2(n51), .A3(n8), .B(n25), .ZN(N353) );
  INVD1BWP30P140 U16 ( .I(n3), .ZN(n6) );
  INVD1BWP30P140 U17 ( .I(n50), .ZN(n4) );
  AN3D4BWP30P140 U18 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n4), .Z(n89) );
  OAI21D1BWP30P140 U19 ( .A1(n6), .A2(i_cmd[1]), .B(n5), .ZN(N354) );
  INVD1BWP30P140 U20 ( .I(i_data_bus[3]), .ZN(n58) );
  MUX2NOPTD2BWP30P140 U21 ( .I0(n7), .I1(n51), .S(i_cmd[1]), .ZN(n10) );
  NR2D1BWP30P140 U22 ( .A1(n50), .A2(n8), .ZN(n9) );
  CKND2D2BWP30P140 U23 ( .A1(n10), .A2(n9), .ZN(n11) );
  INVD2BWP30P140 U24 ( .I(n11), .ZN(n13) );
  INVD2BWP30P140 U25 ( .I(n13), .ZN(n48) );
  INVD1BWP30P140 U26 ( .I(i_data_bus[35]), .ZN(n12) );
  OAI22D1BWP30P140 U27 ( .A1(n25), .A2(n58), .B1(n48), .B2(n12), .ZN(N290) );
  INVD1BWP30P140 U28 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD2BWP30P140 U29 ( .I(n13), .ZN(n46) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[34]), .ZN(n14) );
  OAI22D1BWP30P140 U31 ( .A1(n25), .A2(n62), .B1(n46), .B2(n14), .ZN(N289) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[33]), .ZN(n15) );
  OAI22D1BWP30P140 U34 ( .A1(n25), .A2(n59), .B1(n48), .B2(n15), .ZN(N288) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[0]), .ZN(n63) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[32]), .ZN(n16) );
  OAI22D1BWP30P140 U37 ( .A1(n25), .A2(n63), .B1(n46), .B2(n16), .ZN(N287) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[31]), .ZN(n70) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[63]), .ZN(n17) );
  OAI22D1BWP30P140 U40 ( .A1(n25), .A2(n70), .B1(n48), .B2(n17), .ZN(N318) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[29]), .ZN(n71) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[61]), .ZN(n18) );
  OAI22D1BWP30P140 U43 ( .A1(n25), .A2(n71), .B1(n48), .B2(n18), .ZN(N316) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[27]), .ZN(n72) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[59]), .ZN(n19) );
  OAI22D1BWP30P140 U46 ( .A1(n25), .A2(n72), .B1(n48), .B2(n19), .ZN(N314) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[25]), .ZN(n73) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[57]), .ZN(n20) );
  OAI22D1BWP30P140 U49 ( .A1(n25), .A2(n73), .B1(n48), .B2(n20), .ZN(N312) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[23]), .ZN(n81) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[55]), .ZN(n21) );
  OAI22D1BWP30P140 U52 ( .A1(n25), .A2(n81), .B1(n48), .B2(n21), .ZN(N310) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[21]), .ZN(n83) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[53]), .ZN(n22) );
  OAI22D1BWP30P140 U55 ( .A1(n25), .A2(n83), .B1(n48), .B2(n22), .ZN(N308) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[20]), .ZN(n85) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[52]), .ZN(n23) );
  OAI22D1BWP30P140 U58 ( .A1(n25), .A2(n85), .B1(n48), .B2(n23), .ZN(N307) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[19]), .ZN(n86) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[51]), .ZN(n24) );
  OAI22D1BWP30P140 U61 ( .A1(n25), .A2(n86), .B1(n46), .B2(n24), .ZN(N306) );
  INVD2BWP30P140 U62 ( .I(n26), .ZN(n49) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[40]), .ZN(n27) );
  OAI22D1BWP30P140 U65 ( .A1(n49), .A2(n66), .B1(n46), .B2(n27), .ZN(N295) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[9]), .ZN(n76) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[41]), .ZN(n28) );
  OAI22D1BWP30P140 U68 ( .A1(n49), .A2(n76), .B1(n46), .B2(n28), .ZN(N296) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[10]), .ZN(n65) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[42]), .ZN(n29) );
  OAI22D1BWP30P140 U71 ( .A1(n49), .A2(n65), .B1(n46), .B2(n29), .ZN(N297) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[11]), .ZN(n75) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[43]), .ZN(n30) );
  OAI22D1BWP30P140 U74 ( .A1(n49), .A2(n75), .B1(n46), .B2(n30), .ZN(N298) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[12]), .ZN(n64) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[44]), .ZN(n31) );
  OAI22D1BWP30P140 U77 ( .A1(n49), .A2(n64), .B1(n46), .B2(n31), .ZN(N299) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[13]), .ZN(n74) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[45]), .ZN(n32) );
  OAI22D1BWP30P140 U80 ( .A1(n49), .A2(n74), .B1(n46), .B2(n32), .ZN(N300) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[14]), .ZN(n67) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[46]), .ZN(n33) );
  OAI22D1BWP30P140 U83 ( .A1(n49), .A2(n67), .B1(n46), .B2(n33), .ZN(N301) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[15]), .ZN(n68) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[47]), .ZN(n34) );
  OAI22D1BWP30P140 U86 ( .A1(n49), .A2(n68), .B1(n46), .B2(n34), .ZN(N302) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[16]), .ZN(n91) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[48]), .ZN(n35) );
  OAI22D1BWP30P140 U89 ( .A1(n49), .A2(n91), .B1(n46), .B2(n35), .ZN(N303) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[17]), .ZN(n88) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[49]), .ZN(n36) );
  OAI22D1BWP30P140 U92 ( .A1(n49), .A2(n88), .B1(n46), .B2(n36), .ZN(N304) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[18]), .ZN(n87) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[50]), .ZN(n37) );
  OAI22D1BWP30P140 U95 ( .A1(n49), .A2(n87), .B1(n46), .B2(n37), .ZN(N305) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[22]), .ZN(n82) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[54]), .ZN(n38) );
  OAI22D1BWP30P140 U98 ( .A1(n49), .A2(n82), .B1(n48), .B2(n38), .ZN(N309) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[24]), .ZN(n80) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[56]), .ZN(n39) );
  OAI22D1BWP30P140 U101 ( .A1(n49), .A2(n80), .B1(n48), .B2(n39), .ZN(N311) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[26]), .ZN(n79) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[58]), .ZN(n40) );
  OAI22D1BWP30P140 U104 ( .A1(n49), .A2(n79), .B1(n48), .B2(n40), .ZN(N313) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[28]), .ZN(n78) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[60]), .ZN(n41) );
  OAI22D1BWP30P140 U107 ( .A1(n49), .A2(n78), .B1(n48), .B2(n41), .ZN(N315) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[30]), .ZN(n77) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[62]), .ZN(n42) );
  OAI22D1BWP30P140 U110 ( .A1(n49), .A2(n77), .B1(n48), .B2(n42), .ZN(N317) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[36]), .ZN(n43) );
  OAI22D1BWP30P140 U113 ( .A1(n49), .A2(n61), .B1(n46), .B2(n43), .ZN(N291) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[5]), .ZN(n57) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[37]), .ZN(n44) );
  OAI22D1BWP30P140 U116 ( .A1(n49), .A2(n57), .B1(n48), .B2(n44), .ZN(N292) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[6]), .ZN(n60) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[38]), .ZN(n45) );
  OAI22D1BWP30P140 U119 ( .A1(n49), .A2(n60), .B1(n46), .B2(n45), .ZN(N293) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[39]), .ZN(n47) );
  OAI22D1BWP30P140 U122 ( .A1(n49), .A2(n56), .B1(n48), .B2(n47), .ZN(N294) );
  NR2D1BWP30P140 U123 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  MUX2NUD1BWP30P140 U124 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U126 ( .I(n55), .ZN(n69) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n90), .B1(i_data_bus[39]), .B2(n89), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n90), .B1(i_data_bus[37]), .B2(n89), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n90), .B1(i_data_bus[35]), .B2(n89), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n90), .B1(i_data_bus[33]), .B2(n89), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n90), .B1(i_data_bus[38]), .B2(n89), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n90), .B1(i_data_bus[36]), .B2(n89), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n90), .B1(i_data_bus[34]), .B2(n89), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n90), .B1(i_data_bus[32]), .B2(n89), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n90), .B1(i_data_bus[44]), .B2(n89), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n90), .B1(i_data_bus[42]), .B2(n89), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n90), .B1(i_data_bus[40]), .B2(n89), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n90), .B1(i_data_bus[46]), .B2(n89), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n90), .B1(i_data_bus[47]), .B2(n89), 
        .ZN(N334) );
  INVD2BWP30P140 U140 ( .I(n69), .ZN(n84) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n84), .B1(i_data_bus[63]), .B2(n89), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n84), .B1(i_data_bus[61]), .B2(n89), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n84), .B1(i_data_bus[59]), .B2(n89), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n84), .B1(i_data_bus[57]), .B2(n89), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n90), .B1(i_data_bus[45]), .B2(n89), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n90), .B1(i_data_bus[43]), .B2(n89), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n90), .B1(i_data_bus[41]), .B2(n89), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n84), .B1(i_data_bus[62]), .B2(n89), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n84), .B1(i_data_bus[60]), .B2(n89), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n84), .B1(i_data_bus[58]), .B2(n89), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n84), .B1(i_data_bus[56]), .B2(n89), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n84), .B1(i_data_bus[55]), .B2(n89), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n84), .B1(i_data_bus[54]), .B2(n89), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n84), .B1(i_data_bus[53]), .B2(n89), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n84), .B1(i_data_bus[52]), .B2(n89), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n90), .B1(i_data_bus[51]), .B2(n89), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n90), .B1(i_data_bus[50]), .B2(n89), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n90), .B1(i_data_bus[49]), .B2(n89), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U159 ( .A1(n91), .A2(n90), .B1(i_data_bus[48]), .B2(n89), 
        .ZN(N335) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_7 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90;

  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  ND2OPTIBD1BWP30P140 U3 ( .A1(n9), .A2(n12), .ZN(n7) );
  INR2D1BWP30P140 U4 ( .A1(i_valid[0]), .B1(n13), .ZN(n9) );
  INVD3BWP30P140 U5 ( .I(n67), .ZN(n78) );
  MOAI22D1BWP30P140 U6 ( .A1(n20), .A2(n78), .B1(i_data_bus[34]), .B2(n88), 
        .ZN(N321) );
  INVD1BWP30P140 U7 ( .I(n88), .ZN(n10) );
  INVD1BWP30P140 U8 ( .I(i_data_bus[2]), .ZN(n20) );
  INVD1BWP30P140 U9 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U10 ( .A1(n1), .A2(i_en), .ZN(n13) );
  NR2D1BWP30P140 U11 ( .A1(n13), .A2(i_cmd[1]), .ZN(n4) );
  INVD1BWP30P140 U12 ( .I(i_valid[0]), .ZN(n2) );
  INVD2BWP30P140 U13 ( .I(i_valid[1]), .ZN(n8) );
  MUX2NUD1BWP30P140 U14 ( .I0(n2), .I1(n8), .S(i_cmd[0]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U15 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U16 ( .I(n5), .ZN(n67) );
  INVD1BWP30P140 U17 ( .I(n13), .ZN(n6) );
  AN3D4BWP30P140 U18 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n6), .Z(n88) );
  INVD2BWP30P140 U19 ( .I(i_cmd[0]), .ZN(n12) );
  INVD2BWP30P140 U20 ( .I(n7), .ZN(n32) );
  INVD2BWP30P140 U21 ( .I(n32), .ZN(n31) );
  OAI31D1BWP30P140 U22 ( .A1(n13), .A2(n8), .A3(n12), .B(n31), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n9), .ZN(n11) );
  OAI21D1BWP30P140 U24 ( .A1(n11), .A2(i_cmd[1]), .B(n10), .ZN(N354) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[3]), .ZN(n58) );
  MUX2NOPTD2BWP30P140 U26 ( .I0(n2), .I1(n8), .S(i_cmd[1]), .ZN(n15) );
  NR2D1BWP30P140 U27 ( .A1(n13), .A2(n12), .ZN(n14) );
  CKND2D2BWP30P140 U28 ( .A1(n15), .A2(n14), .ZN(n16) );
  INVD2BWP30P140 U29 ( .I(n16), .ZN(n18) );
  INVD2BWP30P140 U30 ( .I(n18), .ZN(n54) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[35]), .ZN(n17) );
  OAI22D1BWP30P140 U32 ( .A1(n31), .A2(n58), .B1(n54), .B2(n17), .ZN(N290) );
  INVD2BWP30P140 U33 ( .I(n18), .ZN(n52) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[34]), .ZN(n19) );
  OAI22D1BWP30P140 U35 ( .A1(n31), .A2(n20), .B1(n52), .B2(n19), .ZN(N289) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[33]), .ZN(n21) );
  OAI22D1BWP30P140 U38 ( .A1(n31), .A2(n59), .B1(n54), .B2(n21), .ZN(N288) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[0]), .ZN(n61) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[32]), .ZN(n22) );
  OAI22D1BWP30P140 U41 ( .A1(n31), .A2(n61), .B1(n52), .B2(n22), .ZN(N287) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[31]), .ZN(n63) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[63]), .ZN(n23) );
  OAI22D1BWP30P140 U44 ( .A1(n31), .A2(n63), .B1(n54), .B2(n23), .ZN(N318) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[29]), .ZN(n64) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[61]), .ZN(n24) );
  OAI22D1BWP30P140 U47 ( .A1(n31), .A2(n64), .B1(n54), .B2(n24), .ZN(N316) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[27]), .ZN(n65) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[59]), .ZN(n25) );
  OAI22D1BWP30P140 U50 ( .A1(n31), .A2(n65), .B1(n54), .B2(n25), .ZN(N314) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[25]), .ZN(n66) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[57]), .ZN(n26) );
  OAI22D1BWP30P140 U53 ( .A1(n31), .A2(n66), .B1(n54), .B2(n26), .ZN(N312) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[23]), .ZN(n75) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[55]), .ZN(n27) );
  OAI22D1BWP30P140 U56 ( .A1(n31), .A2(n75), .B1(n54), .B2(n27), .ZN(N310) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[21]), .ZN(n77) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[53]), .ZN(n28) );
  OAI22D1BWP30P140 U59 ( .A1(n31), .A2(n77), .B1(n54), .B2(n28), .ZN(N308) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[52]), .ZN(n29) );
  OAI22D1BWP30P140 U62 ( .A1(n31), .A2(n79), .B1(n54), .B2(n29), .ZN(N307) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[19]), .ZN(n80) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[51]), .ZN(n30) );
  OAI22D1BWP30P140 U65 ( .A1(n31), .A2(n80), .B1(n52), .B2(n30), .ZN(N306) );
  INVD2BWP30P140 U66 ( .I(n32), .ZN(n55) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[8]), .ZN(n90) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[40]), .ZN(n33) );
  OAI22D1BWP30P140 U69 ( .A1(n55), .A2(n90), .B1(n52), .B2(n33), .ZN(N295) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[9]), .ZN(n70) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[41]), .ZN(n34) );
  OAI22D1BWP30P140 U72 ( .A1(n55), .A2(n70), .B1(n52), .B2(n34), .ZN(N296) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[10]), .ZN(n87) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[42]), .ZN(n35) );
  OAI22D1BWP30P140 U75 ( .A1(n55), .A2(n87), .B1(n52), .B2(n35), .ZN(N297) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[43]), .ZN(n36) );
  OAI22D1BWP30P140 U78 ( .A1(n55), .A2(n69), .B1(n52), .B2(n36), .ZN(N298) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[44]), .ZN(n37) );
  OAI22D1BWP30P140 U81 ( .A1(n55), .A2(n86), .B1(n52), .B2(n37), .ZN(N299) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[13]), .ZN(n68) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[45]), .ZN(n38) );
  OAI22D1BWP30P140 U84 ( .A1(n55), .A2(n68), .B1(n52), .B2(n38), .ZN(N300) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[14]), .ZN(n85) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[46]), .ZN(n39) );
  OAI22D1BWP30P140 U87 ( .A1(n55), .A2(n85), .B1(n52), .B2(n39), .ZN(N301) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[15]), .ZN(n84) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[47]), .ZN(n40) );
  OAI22D1BWP30P140 U90 ( .A1(n55), .A2(n84), .B1(n52), .B2(n40), .ZN(N302) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[16]), .ZN(n83) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[48]), .ZN(n41) );
  OAI22D1BWP30P140 U93 ( .A1(n55), .A2(n83), .B1(n52), .B2(n41), .ZN(N303) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[17]), .ZN(n82) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[49]), .ZN(n42) );
  OAI22D1BWP30P140 U96 ( .A1(n55), .A2(n82), .B1(n52), .B2(n42), .ZN(N304) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[18]), .ZN(n81) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[50]), .ZN(n43) );
  OAI22D1BWP30P140 U99 ( .A1(n55), .A2(n81), .B1(n52), .B2(n43), .ZN(N305) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[22]), .ZN(n76) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[54]), .ZN(n44) );
  OAI22D1BWP30P140 U102 ( .A1(n55), .A2(n76), .B1(n54), .B2(n44), .ZN(N309) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[24]), .ZN(n74) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[56]), .ZN(n45) );
  OAI22D1BWP30P140 U105 ( .A1(n55), .A2(n74), .B1(n54), .B2(n45), .ZN(N311) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[26]), .ZN(n73) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[58]), .ZN(n46) );
  OAI22D1BWP30P140 U108 ( .A1(n55), .A2(n73), .B1(n54), .B2(n46), .ZN(N313) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[28]), .ZN(n72) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[60]), .ZN(n47) );
  OAI22D1BWP30P140 U111 ( .A1(n55), .A2(n72), .B1(n54), .B2(n47), .ZN(N315) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[30]), .ZN(n71) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[62]), .ZN(n48) );
  OAI22D1BWP30P140 U114 ( .A1(n55), .A2(n71), .B1(n54), .B2(n48), .ZN(N317) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[36]), .ZN(n49) );
  OAI22D1BWP30P140 U117 ( .A1(n55), .A2(n60), .B1(n52), .B2(n49), .ZN(N291) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[5]), .ZN(n57) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[37]), .ZN(n50) );
  OAI22D1BWP30P140 U120 ( .A1(n55), .A2(n57), .B1(n54), .B2(n50), .ZN(N292) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[6]), .ZN(n62) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[38]), .ZN(n51) );
  OAI22D1BWP30P140 U123 ( .A1(n55), .A2(n62), .B1(n52), .B2(n51), .ZN(N293) );
  INVD1BWP30P140 U124 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD1BWP30P140 U125 ( .I(i_data_bus[39]), .ZN(n53) );
  OAI22D1BWP30P140 U126 ( .A1(n55), .A2(n56), .B1(n54), .B2(n53), .ZN(N294) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n78), .B1(i_data_bus[39]), .B2(n88), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n78), .B1(i_data_bus[37]), .B2(n88), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n78), .B1(i_data_bus[35]), .B2(n88), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n78), .B1(i_data_bus[33]), .B2(n88), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n78), .B1(i_data_bus[36]), .B2(n88), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n78), .B1(i_data_bus[32]), .B2(n88), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n78), .B1(i_data_bus[38]), .B2(n88), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n78), .B1(i_data_bus[63]), .B2(n88), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n78), .B1(i_data_bus[61]), .B2(n88), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n78), .B1(i_data_bus[59]), .B2(n88), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n78), .B1(i_data_bus[57]), .B2(n88), 
        .ZN(N344) );
  INVD2BWP30P140 U138 ( .I(n67), .ZN(n89) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n89), .B1(i_data_bus[45]), .B2(n88), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n89), .B1(i_data_bus[43]), .B2(n88), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n89), .B1(i_data_bus[41]), .B2(n88), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n78), .B1(i_data_bus[62]), .B2(n88), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n78), .B1(i_data_bus[60]), .B2(n88), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n78), .B1(i_data_bus[58]), .B2(n88), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n78), .B1(i_data_bus[56]), .B2(n88), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n78), .B1(i_data_bus[55]), .B2(n88), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n78), .B1(i_data_bus[54]), .B2(n88), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n78), .B1(i_data_bus[53]), .B2(n88), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n78), .B1(i_data_bus[52]), .B2(n88), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n89), .B1(i_data_bus[51]), .B2(n88), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n89), .B1(i_data_bus[50]), .B2(n88), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n89), .B1(i_data_bus[49]), .B2(n88), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n89), .B1(i_data_bus[48]), .B2(n88), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n89), .B1(i_data_bus[47]), .B2(n88), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n89), .B1(i_data_bus[46]), .B2(n88), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n89), .B1(i_data_bus[44]), .B2(n88), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n89), .B1(i_data_bus[42]), .B2(n88), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U158 ( .A1(n90), .A2(n89), .B1(i_data_bus[40]), .B2(n88), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_8 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90;

  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  ND2OPTIBD1BWP30P140 U3 ( .A1(n9), .A2(n12), .ZN(n7) );
  INVD3BWP30P140 U4 ( .I(n71), .ZN(n84) );
  MOAI22D1BWP30P140 U5 ( .A1(n54), .A2(n84), .B1(i_data_bus[39]), .B2(n88), 
        .ZN(N326) );
  INVD1BWP30P140 U6 ( .I(n88), .ZN(n10) );
  INVD1BWP30P140 U7 ( .I(i_data_bus[7]), .ZN(n54) );
  INVD1BWP30P140 U8 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U9 ( .A1(n1), .A2(i_en), .ZN(n13) );
  NR2D1BWP30P140 U10 ( .A1(n13), .A2(i_cmd[1]), .ZN(n4) );
  INVD2BWP30P140 U11 ( .I(i_valid[0]), .ZN(n2) );
  INVD1BWP30P140 U12 ( .I(i_valid[1]), .ZN(n8) );
  MUX2NUD1BWP30P140 U13 ( .I0(n2), .I1(n8), .S(i_cmd[0]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U14 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U15 ( .I(n5), .ZN(n71) );
  INVD1BWP30P140 U16 ( .I(n13), .ZN(n6) );
  AN3D4BWP30P140 U17 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n6), .Z(n88) );
  INVD2BWP30P140 U18 ( .I(i_cmd[0]), .ZN(n12) );
  INR2D2BWP30P140 U19 ( .A1(i_valid[0]), .B1(n13), .ZN(n9) );
  INVD2BWP30P140 U20 ( .I(n7), .ZN(n31) );
  INVD2BWP30P140 U21 ( .I(n31), .ZN(n30) );
  OAI31D1BWP30P140 U22 ( .A1(n13), .A2(n8), .A3(n12), .B(n30), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n9), .ZN(n11) );
  OAI21D1BWP30P140 U24 ( .A1(n11), .A2(i_cmd[1]), .B(n10), .ZN(N354) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[21]), .ZN(n69) );
  MUX2NUD1BWP30P140 U26 ( .I0(n2), .I1(n8), .S(i_cmd[1]), .ZN(n15) );
  NR2D1BWP30P140 U27 ( .A1(n13), .A2(n12), .ZN(n14) );
  CKND2D2BWP30P140 U28 ( .A1(n15), .A2(n14), .ZN(n16) );
  INVD2BWP30P140 U29 ( .I(n16), .ZN(n19) );
  INVD2BWP30P140 U30 ( .I(n19), .ZN(n53) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[53]), .ZN(n17) );
  OAI22D1BWP30P140 U32 ( .A1(n30), .A2(n69), .B1(n53), .B2(n17), .ZN(N308) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[23]), .ZN(n67) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[55]), .ZN(n18) );
  OAI22D1BWP30P140 U35 ( .A1(n30), .A2(n67), .B1(n53), .B2(n18), .ZN(N310) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[19]), .ZN(n72) );
  INVD2BWP30P140 U37 ( .I(n19), .ZN(n51) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[51]), .ZN(n20) );
  OAI22D1BWP30P140 U39 ( .A1(n30), .A2(n72), .B1(n51), .B2(n20), .ZN(N306) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[20]), .ZN(n70) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[52]), .ZN(n21) );
  OAI22D1BWP30P140 U42 ( .A1(n30), .A2(n70), .B1(n53), .B2(n21), .ZN(N307) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[25]), .ZN(n85) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[57]), .ZN(n22) );
  OAI22D1BWP30P140 U45 ( .A1(n30), .A2(n85), .B1(n53), .B2(n22), .ZN(N312) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[27]), .ZN(n83) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[59]), .ZN(n23) );
  OAI22D1BWP30P140 U48 ( .A1(n30), .A2(n83), .B1(n53), .B2(n23), .ZN(N314) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[29]), .ZN(n82) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[61]), .ZN(n24) );
  OAI22D1BWP30P140 U51 ( .A1(n30), .A2(n82), .B1(n53), .B2(n24), .ZN(N316) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[31]), .ZN(n81) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[63]), .ZN(n25) );
  OAI22D1BWP30P140 U54 ( .A1(n30), .A2(n81), .B1(n53), .B2(n25), .ZN(N318) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[0]), .ZN(n59) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[32]), .ZN(n26) );
  OAI22D1BWP30P140 U57 ( .A1(n30), .A2(n59), .B1(n51), .B2(n26), .ZN(N287) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[1]), .ZN(n60) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[33]), .ZN(n27) );
  OAI22D1BWP30P140 U60 ( .A1(n30), .A2(n60), .B1(n53), .B2(n27), .ZN(N288) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[2]), .ZN(n58) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[34]), .ZN(n28) );
  OAI22D1BWP30P140 U63 ( .A1(n30), .A2(n58), .B1(n51), .B2(n28), .ZN(N289) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[35]), .ZN(n29) );
  OAI22D1BWP30P140 U66 ( .A1(n30), .A2(n61), .B1(n53), .B2(n29), .ZN(N290) );
  INVD2BWP30P140 U67 ( .I(n31), .ZN(n55) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[8]), .ZN(n80) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[40]), .ZN(n32) );
  OAI22D1BWP30P140 U70 ( .A1(n55), .A2(n80), .B1(n51), .B2(n32), .ZN(N295) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[9]), .ZN(n90) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[41]), .ZN(n33) );
  OAI22D1BWP30P140 U73 ( .A1(n55), .A2(n90), .B1(n51), .B2(n33), .ZN(N296) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[10]), .ZN(n79) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[42]), .ZN(n34) );
  OAI22D1BWP30P140 U76 ( .A1(n55), .A2(n79), .B1(n51), .B2(n34), .ZN(N297) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[11]), .ZN(n87) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[43]), .ZN(n35) );
  OAI22D1BWP30P140 U79 ( .A1(n55), .A2(n87), .B1(n51), .B2(n35), .ZN(N298) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[12]), .ZN(n78) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[44]), .ZN(n36) );
  OAI22D1BWP30P140 U82 ( .A1(n55), .A2(n78), .B1(n51), .B2(n36), .ZN(N299) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[13]), .ZN(n86) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[45]), .ZN(n37) );
  OAI22D1BWP30P140 U85 ( .A1(n55), .A2(n86), .B1(n51), .B2(n37), .ZN(N300) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[14]), .ZN(n77) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[46]), .ZN(n38) );
  OAI22D1BWP30P140 U88 ( .A1(n55), .A2(n77), .B1(n51), .B2(n38), .ZN(N301) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[15]), .ZN(n76) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[47]), .ZN(n39) );
  OAI22D1BWP30P140 U91 ( .A1(n55), .A2(n76), .B1(n51), .B2(n39), .ZN(N302) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[16]), .ZN(n75) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[48]), .ZN(n40) );
  OAI22D1BWP30P140 U94 ( .A1(n55), .A2(n75), .B1(n51), .B2(n40), .ZN(N303) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[49]), .ZN(n41) );
  OAI22D1BWP30P140 U97 ( .A1(n55), .A2(n74), .B1(n51), .B2(n41), .ZN(N304) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[18]), .ZN(n73) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[50]), .ZN(n42) );
  OAI22D1BWP30P140 U100 ( .A1(n55), .A2(n73), .B1(n51), .B2(n42), .ZN(N305) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[22]), .ZN(n68) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[54]), .ZN(n43) );
  OAI22D1BWP30P140 U103 ( .A1(n55), .A2(n68), .B1(n53), .B2(n43), .ZN(N309) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[24]), .ZN(n66) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[56]), .ZN(n44) );
  OAI22D1BWP30P140 U106 ( .A1(n55), .A2(n66), .B1(n53), .B2(n44), .ZN(N311) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[26]), .ZN(n65) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[58]), .ZN(n45) );
  OAI22D1BWP30P140 U109 ( .A1(n55), .A2(n65), .B1(n53), .B2(n45), .ZN(N313) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[28]), .ZN(n64) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[60]), .ZN(n46) );
  OAI22D1BWP30P140 U112 ( .A1(n55), .A2(n64), .B1(n53), .B2(n46), .ZN(N315) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[30]), .ZN(n63) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[62]), .ZN(n47) );
  OAI22D1BWP30P140 U115 ( .A1(n55), .A2(n63), .B1(n53), .B2(n47), .ZN(N317) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[4]), .ZN(n57) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[36]), .ZN(n48) );
  OAI22D1BWP30P140 U118 ( .A1(n55), .A2(n57), .B1(n51), .B2(n48), .ZN(N291) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[37]), .ZN(n49) );
  OAI22D1BWP30P140 U121 ( .A1(n55), .A2(n62), .B1(n53), .B2(n49), .ZN(N292) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[6]), .ZN(n56) );
  INVD1BWP30P140 U123 ( .I(i_data_bus[38]), .ZN(n50) );
  OAI22D1BWP30P140 U124 ( .A1(n55), .A2(n56), .B1(n51), .B2(n50), .ZN(N293) );
  INVD1BWP30P140 U125 ( .I(i_data_bus[39]), .ZN(n52) );
  OAI22D1BWP30P140 U126 ( .A1(n55), .A2(n54), .B1(n53), .B2(n52), .ZN(N294) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n84), .B1(i_data_bus[38]), .B2(n88), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n84), .B1(i_data_bus[36]), .B2(n88), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n84), .B1(i_data_bus[34]), .B2(n88), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n84), .B1(i_data_bus[32]), .B2(n88), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n84), .B1(i_data_bus[33]), .B2(n88), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n84), .B1(i_data_bus[35]), .B2(n88), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n84), .B1(i_data_bus[37]), .B2(n88), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n84), .B1(i_data_bus[62]), .B2(n88), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n84), .B1(i_data_bus[60]), .B2(n88), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n84), .B1(i_data_bus[58]), .B2(n88), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n84), .B1(i_data_bus[56]), .B2(n88), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n84), .B1(i_data_bus[55]), .B2(n88), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n84), .B1(i_data_bus[54]), .B2(n88), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n84), .B1(i_data_bus[53]), .B2(n88), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n84), .B1(i_data_bus[52]), .B2(n88), 
        .ZN(N339) );
  INVD2BWP30P140 U142 ( .I(n71), .ZN(n89) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n89), .B1(i_data_bus[51]), .B2(n88), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n89), .B1(i_data_bus[50]), .B2(n88), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n89), .B1(i_data_bus[49]), .B2(n88), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n89), .B1(i_data_bus[48]), .B2(n88), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n89), .B1(i_data_bus[47]), .B2(n88), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n89), .B1(i_data_bus[46]), .B2(n88), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n89), .B1(i_data_bus[44]), .B2(n88), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n89), .B1(i_data_bus[42]), .B2(n88), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n89), .B1(i_data_bus[40]), .B2(n88), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n84), .B1(i_data_bus[63]), .B2(n88), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n84), .B1(i_data_bus[61]), .B2(n88), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n84), .B1(i_data_bus[59]), .B2(n88), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n84), .B1(i_data_bus[57]), .B2(n88), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n89), .B1(i_data_bus[45]), .B2(n88), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n89), .B1(i_data_bus[43]), .B2(n88), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n90), .A2(n89), .B1(i_data_bus[41]), .B2(n88), 
        .ZN(N328) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_9 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90;

  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  ND2OPTIBD1BWP30P140 U3 ( .A1(n9), .A2(n12), .ZN(n7) );
  INVD3BWP30P140 U4 ( .I(n67), .ZN(n78) );
  MOAI22D1BWP30P140 U5 ( .A1(n27), .A2(n78), .B1(i_data_bus[32]), .B2(n88), 
        .ZN(N319) );
  INVD1BWP30P140 U6 ( .I(n88), .ZN(n10) );
  INVD1BWP30P140 U7 ( .I(i_data_bus[0]), .ZN(n27) );
  INVD1BWP30P140 U8 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U9 ( .A1(n1), .A2(i_en), .ZN(n13) );
  NR2D1BWP30P140 U10 ( .A1(n13), .A2(i_cmd[1]), .ZN(n4) );
  INVD2BWP30P140 U11 ( .I(i_valid[0]), .ZN(n2) );
  INVD1BWP30P140 U12 ( .I(i_valid[1]), .ZN(n8) );
  MUX2NUD1BWP30P140 U13 ( .I0(n2), .I1(n8), .S(i_cmd[0]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U14 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U15 ( .I(n5), .ZN(n67) );
  INVD1BWP30P140 U16 ( .I(n13), .ZN(n6) );
  AN3D4BWP30P140 U17 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n6), .Z(n88) );
  INVD2BWP30P140 U18 ( .I(i_cmd[0]), .ZN(n12) );
  INR2D2BWP30P140 U19 ( .A1(i_valid[0]), .B1(n13), .ZN(n9) );
  INVD2BWP30P140 U20 ( .I(n7), .ZN(n32) );
  INVD2BWP30P140 U21 ( .I(n32), .ZN(n31) );
  OAI31D1BWP30P140 U22 ( .A1(n13), .A2(n8), .A3(n12), .B(n31), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n9), .ZN(n11) );
  OAI21D1BWP30P140 U24 ( .A1(n11), .A2(i_cmd[1]), .B(n10), .ZN(N354) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[19]), .ZN(n80) );
  MUX2NUD1BWP30P140 U26 ( .I0(n2), .I1(n8), .S(i_cmd[1]), .ZN(n15) );
  NR2D1BWP30P140 U27 ( .A1(n13), .A2(n12), .ZN(n14) );
  CKND2D2BWP30P140 U28 ( .A1(n15), .A2(n14), .ZN(n16) );
  INVD2BWP30P140 U29 ( .I(n16), .ZN(n18) );
  INVD2BWP30P140 U30 ( .I(n18), .ZN(n54) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[51]), .ZN(n17) );
  OAI22D1BWP30P140 U32 ( .A1(n31), .A2(n80), .B1(n54), .B2(n17), .ZN(N306) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD2BWP30P140 U34 ( .I(n18), .ZN(n42) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[52]), .ZN(n19) );
  OAI22D1BWP30P140 U36 ( .A1(n31), .A2(n79), .B1(n42), .B2(n19), .ZN(N307) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[21]), .ZN(n77) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[53]), .ZN(n20) );
  OAI22D1BWP30P140 U39 ( .A1(n31), .A2(n77), .B1(n42), .B2(n20), .ZN(N308) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[23]), .ZN(n75) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[55]), .ZN(n21) );
  OAI22D1BWP30P140 U42 ( .A1(n31), .A2(n75), .B1(n42), .B2(n21), .ZN(N310) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[25]), .ZN(n66) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[57]), .ZN(n22) );
  OAI22D1BWP30P140 U45 ( .A1(n31), .A2(n66), .B1(n42), .B2(n22), .ZN(N312) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[27]), .ZN(n65) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[59]), .ZN(n23) );
  OAI22D1BWP30P140 U48 ( .A1(n31), .A2(n65), .B1(n42), .B2(n23), .ZN(N314) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[29]), .ZN(n64) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[61]), .ZN(n24) );
  OAI22D1BWP30P140 U51 ( .A1(n31), .A2(n64), .B1(n42), .B2(n24), .ZN(N316) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[31]), .ZN(n63) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[63]), .ZN(n25) );
  OAI22D1BWP30P140 U54 ( .A1(n31), .A2(n63), .B1(n42), .B2(n25), .ZN(N318) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[32]), .ZN(n26) );
  OAI22D1BWP30P140 U56 ( .A1(n31), .A2(n27), .B1(n54), .B2(n26), .ZN(N287) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[33]), .ZN(n28) );
  OAI22D1BWP30P140 U59 ( .A1(n31), .A2(n59), .B1(n42), .B2(n28), .ZN(N288) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[34]), .ZN(n29) );
  OAI22D1BWP30P140 U62 ( .A1(n31), .A2(n62), .B1(n54), .B2(n29), .ZN(N289) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[3]), .ZN(n58) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[35]), .ZN(n30) );
  OAI22D1BWP30P140 U65 ( .A1(n31), .A2(n58), .B1(n42), .B2(n30), .ZN(N290) );
  INVD2BWP30P140 U66 ( .I(n32), .ZN(n55) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[26]), .ZN(n73) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[58]), .ZN(n33) );
  OAI22D1BWP30P140 U69 ( .A1(n55), .A2(n73), .B1(n42), .B2(n33), .ZN(N313) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[28]), .ZN(n72) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[60]), .ZN(n34) );
  OAI22D1BWP30P140 U72 ( .A1(n55), .A2(n72), .B1(n42), .B2(n34), .ZN(N315) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[30]), .ZN(n71) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[62]), .ZN(n35) );
  OAI22D1BWP30P140 U75 ( .A1(n55), .A2(n71), .B1(n42), .B2(n35), .ZN(N317) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[36]), .ZN(n36) );
  OAI22D1BWP30P140 U78 ( .A1(n55), .A2(n61), .B1(n54), .B2(n36), .ZN(N291) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[5]), .ZN(n57) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[37]), .ZN(n37) );
  OAI22D1BWP30P140 U81 ( .A1(n55), .A2(n57), .B1(n42), .B2(n37), .ZN(N292) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[6]), .ZN(n60) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[38]), .ZN(n38) );
  OAI22D1BWP30P140 U84 ( .A1(n55), .A2(n60), .B1(n54), .B2(n38), .ZN(N293) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[39]), .ZN(n39) );
  OAI22D1BWP30P140 U87 ( .A1(n55), .A2(n56), .B1(n42), .B2(n39), .ZN(N294) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[24]), .ZN(n74) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[56]), .ZN(n40) );
  OAI22D1BWP30P140 U90 ( .A1(n55), .A2(n74), .B1(n42), .B2(n40), .ZN(N311) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[22]), .ZN(n76) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[54]), .ZN(n41) );
  OAI22D1BWP30P140 U93 ( .A1(n55), .A2(n76), .B1(n42), .B2(n41), .ZN(N309) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[18]), .ZN(n81) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[50]), .ZN(n43) );
  OAI22D1BWP30P140 U96 ( .A1(n55), .A2(n81), .B1(n54), .B2(n43), .ZN(N305) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[17]), .ZN(n82) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[49]), .ZN(n44) );
  OAI22D1BWP30P140 U99 ( .A1(n55), .A2(n82), .B1(n54), .B2(n44), .ZN(N304) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[16]), .ZN(n83) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[48]), .ZN(n45) );
  OAI22D1BWP30P140 U102 ( .A1(n55), .A2(n83), .B1(n54), .B2(n45), .ZN(N303) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[15]), .ZN(n84) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[47]), .ZN(n46) );
  OAI22D1BWP30P140 U105 ( .A1(n55), .A2(n84), .B1(n54), .B2(n46), .ZN(N302) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[14]), .ZN(n85) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[46]), .ZN(n47) );
  OAI22D1BWP30P140 U108 ( .A1(n55), .A2(n85), .B1(n54), .B2(n47), .ZN(N301) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[13]), .ZN(n68) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[45]), .ZN(n48) );
  OAI22D1BWP30P140 U111 ( .A1(n55), .A2(n68), .B1(n54), .B2(n48), .ZN(N300) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[44]), .ZN(n49) );
  OAI22D1BWP30P140 U114 ( .A1(n55), .A2(n86), .B1(n54), .B2(n49), .ZN(N299) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[43]), .ZN(n50) );
  OAI22D1BWP30P140 U117 ( .A1(n55), .A2(n69), .B1(n54), .B2(n50), .ZN(N298) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[10]), .ZN(n87) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[42]), .ZN(n51) );
  OAI22D1BWP30P140 U120 ( .A1(n55), .A2(n87), .B1(n54), .B2(n51), .ZN(N297) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[9]), .ZN(n70) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[41]), .ZN(n52) );
  OAI22D1BWP30P140 U123 ( .A1(n55), .A2(n70), .B1(n54), .B2(n52), .ZN(N296) );
  INVD1BWP30P140 U124 ( .I(i_data_bus[8]), .ZN(n90) );
  INVD1BWP30P140 U125 ( .I(i_data_bus[40]), .ZN(n53) );
  OAI22D1BWP30P140 U126 ( .A1(n55), .A2(n90), .B1(n54), .B2(n53), .ZN(N295) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n78), .B1(i_data_bus[39]), .B2(n88), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n78), .B1(i_data_bus[37]), .B2(n88), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n78), .B1(i_data_bus[35]), .B2(n88), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n78), .B1(i_data_bus[33]), .B2(n88), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n78), .B1(i_data_bus[38]), .B2(n88), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n78), .B1(i_data_bus[36]), .B2(n88), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n78), .B1(i_data_bus[34]), .B2(n88), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n78), .B1(i_data_bus[63]), .B2(n88), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n78), .B1(i_data_bus[61]), .B2(n88), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n78), .B1(i_data_bus[59]), .B2(n88), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n78), .B1(i_data_bus[57]), .B2(n88), 
        .ZN(N344) );
  INVD2BWP30P140 U138 ( .I(n67), .ZN(n89) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n89), .B1(i_data_bus[45]), .B2(n88), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n89), .B1(i_data_bus[43]), .B2(n88), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n89), .B1(i_data_bus[41]), .B2(n88), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n78), .B1(i_data_bus[62]), .B2(n88), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n78), .B1(i_data_bus[60]), .B2(n88), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n78), .B1(i_data_bus[58]), .B2(n88), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n78), .B1(i_data_bus[56]), .B2(n88), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n78), .B1(i_data_bus[55]), .B2(n88), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n78), .B1(i_data_bus[54]), .B2(n88), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n78), .B1(i_data_bus[53]), .B2(n88), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n78), .B1(i_data_bus[52]), .B2(n88), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n89), .B1(i_data_bus[51]), .B2(n88), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n89), .B1(i_data_bus[50]), .B2(n88), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n89), .B1(i_data_bus[49]), .B2(n88), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n89), .B1(i_data_bus[48]), .B2(n88), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n89), .B1(i_data_bus[47]), .B2(n88), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n89), .B1(i_data_bus[46]), .B2(n88), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n89), .B1(i_data_bus[44]), .B2(n88), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n89), .B1(i_data_bus[42]), .B2(n88), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U158 ( .A1(n90), .A2(n89), .B1(i_data_bus[40]), .B2(n88), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_10 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90;

  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  ND2OPTIBD1BWP30P140 U3 ( .A1(n9), .A2(n12), .ZN(n7) );
  INVD3BWP30P140 U4 ( .I(n67), .ZN(n78) );
  MOAI22D1BWP30P140 U5 ( .A1(n26), .A2(n78), .B1(i_data_bus[32]), .B2(n88), 
        .ZN(N319) );
  INVD1BWP30P140 U6 ( .I(n88), .ZN(n10) );
  INVD1BWP30P140 U7 ( .I(i_data_bus[0]), .ZN(n26) );
  INVD1BWP30P140 U8 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U9 ( .A1(n1), .A2(i_en), .ZN(n13) );
  NR2D1BWP30P140 U10 ( .A1(n13), .A2(i_cmd[1]), .ZN(n4) );
  INVD2BWP30P140 U11 ( .I(i_valid[0]), .ZN(n2) );
  INVD1BWP30P140 U12 ( .I(i_valid[1]), .ZN(n8) );
  MUX2NUD1BWP30P140 U13 ( .I0(n2), .I1(n8), .S(i_cmd[0]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U14 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U15 ( .I(n5), .ZN(n67) );
  INVD1BWP30P140 U16 ( .I(n13), .ZN(n6) );
  AN3D4BWP30P140 U17 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n6), .Z(n88) );
  INVD2BWP30P140 U18 ( .I(i_cmd[0]), .ZN(n12) );
  INR2D2BWP30P140 U19 ( .A1(i_valid[0]), .B1(n13), .ZN(n9) );
  INVD2BWP30P140 U20 ( .I(n7), .ZN(n32) );
  INVD2BWP30P140 U21 ( .I(n32), .ZN(n31) );
  OAI31D1BWP30P140 U22 ( .A1(n13), .A2(n8), .A3(n12), .B(n31), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n9), .ZN(n11) );
  OAI21D1BWP30P140 U24 ( .A1(n11), .A2(i_cmd[1]), .B(n10), .ZN(N354) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[23]), .ZN(n75) );
  MUX2NUD1BWP30P140 U26 ( .I0(n2), .I1(n8), .S(i_cmd[1]), .ZN(n15) );
  NR2D1BWP30P140 U27 ( .A1(n13), .A2(n12), .ZN(n14) );
  CKND2D2BWP30P140 U28 ( .A1(n15), .A2(n14), .ZN(n16) );
  INVD2BWP30P140 U29 ( .I(n16), .ZN(n21) );
  INVD2BWP30P140 U30 ( .I(n21), .ZN(n42) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[55]), .ZN(n17) );
  OAI22D1BWP30P140 U32 ( .A1(n31), .A2(n75), .B1(n42), .B2(n17), .ZN(N310) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[25]), .ZN(n66) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[57]), .ZN(n18) );
  OAI22D1BWP30P140 U35 ( .A1(n31), .A2(n66), .B1(n42), .B2(n18), .ZN(N312) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[52]), .ZN(n19) );
  OAI22D1BWP30P140 U38 ( .A1(n31), .A2(n79), .B1(n42), .B2(n19), .ZN(N307) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[27]), .ZN(n65) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[59]), .ZN(n20) );
  OAI22D1BWP30P140 U41 ( .A1(n31), .A2(n65), .B1(n42), .B2(n20), .ZN(N314) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[19]), .ZN(n80) );
  INVD2BWP30P140 U43 ( .I(n21), .ZN(n54) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[51]), .ZN(n22) );
  OAI22D1BWP30P140 U45 ( .A1(n31), .A2(n80), .B1(n54), .B2(n22), .ZN(N306) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[29]), .ZN(n64) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[61]), .ZN(n23) );
  OAI22D1BWP30P140 U48 ( .A1(n31), .A2(n64), .B1(n42), .B2(n23), .ZN(N316) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[31]), .ZN(n63) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[63]), .ZN(n24) );
  OAI22D1BWP30P140 U51 ( .A1(n31), .A2(n63), .B1(n42), .B2(n24), .ZN(N318) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[32]), .ZN(n25) );
  OAI22D1BWP30P140 U53 ( .A1(n31), .A2(n26), .B1(n54), .B2(n25), .ZN(N287) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[33]), .ZN(n27) );
  OAI22D1BWP30P140 U56 ( .A1(n31), .A2(n59), .B1(n42), .B2(n27), .ZN(N288) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[34]), .ZN(n28) );
  OAI22D1BWP30P140 U59 ( .A1(n31), .A2(n62), .B1(n54), .B2(n28), .ZN(N289) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[3]), .ZN(n58) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[35]), .ZN(n29) );
  OAI22D1BWP30P140 U62 ( .A1(n31), .A2(n58), .B1(n42), .B2(n29), .ZN(N290) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[21]), .ZN(n77) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[53]), .ZN(n30) );
  OAI22D1BWP30P140 U65 ( .A1(n31), .A2(n77), .B1(n42), .B2(n30), .ZN(N308) );
  INVD2BWP30P140 U66 ( .I(n32), .ZN(n55) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[39]), .ZN(n33) );
  OAI22D1BWP30P140 U69 ( .A1(n55), .A2(n56), .B1(n42), .B2(n33), .ZN(N294) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[6]), .ZN(n60) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[38]), .ZN(n34) );
  OAI22D1BWP30P140 U72 ( .A1(n55), .A2(n60), .B1(n54), .B2(n34), .ZN(N293) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[5]), .ZN(n57) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[37]), .ZN(n35) );
  OAI22D1BWP30P140 U75 ( .A1(n55), .A2(n57), .B1(n42), .B2(n35), .ZN(N292) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[36]), .ZN(n36) );
  OAI22D1BWP30P140 U78 ( .A1(n55), .A2(n61), .B1(n54), .B2(n36), .ZN(N291) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[30]), .ZN(n71) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[62]), .ZN(n37) );
  OAI22D1BWP30P140 U81 ( .A1(n55), .A2(n71), .B1(n42), .B2(n37), .ZN(N317) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[28]), .ZN(n72) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[60]), .ZN(n38) );
  OAI22D1BWP30P140 U84 ( .A1(n55), .A2(n72), .B1(n42), .B2(n38), .ZN(N315) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[26]), .ZN(n73) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[58]), .ZN(n39) );
  OAI22D1BWP30P140 U87 ( .A1(n55), .A2(n73), .B1(n42), .B2(n39), .ZN(N313) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[24]), .ZN(n74) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[56]), .ZN(n40) );
  OAI22D1BWP30P140 U90 ( .A1(n55), .A2(n74), .B1(n42), .B2(n40), .ZN(N311) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[22]), .ZN(n76) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[54]), .ZN(n41) );
  OAI22D1BWP30P140 U93 ( .A1(n55), .A2(n76), .B1(n42), .B2(n41), .ZN(N309) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[18]), .ZN(n81) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[50]), .ZN(n43) );
  OAI22D1BWP30P140 U96 ( .A1(n55), .A2(n81), .B1(n54), .B2(n43), .ZN(N305) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[17]), .ZN(n82) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[49]), .ZN(n44) );
  OAI22D1BWP30P140 U99 ( .A1(n55), .A2(n82), .B1(n54), .B2(n44), .ZN(N304) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[16]), .ZN(n83) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[48]), .ZN(n45) );
  OAI22D1BWP30P140 U102 ( .A1(n55), .A2(n83), .B1(n54), .B2(n45), .ZN(N303) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[15]), .ZN(n84) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[47]), .ZN(n46) );
  OAI22D1BWP30P140 U105 ( .A1(n55), .A2(n84), .B1(n54), .B2(n46), .ZN(N302) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[14]), .ZN(n85) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[46]), .ZN(n47) );
  OAI22D1BWP30P140 U108 ( .A1(n55), .A2(n85), .B1(n54), .B2(n47), .ZN(N301) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[13]), .ZN(n68) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[45]), .ZN(n48) );
  OAI22D1BWP30P140 U111 ( .A1(n55), .A2(n68), .B1(n54), .B2(n48), .ZN(N300) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[44]), .ZN(n49) );
  OAI22D1BWP30P140 U114 ( .A1(n55), .A2(n86), .B1(n54), .B2(n49), .ZN(N299) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[43]), .ZN(n50) );
  OAI22D1BWP30P140 U117 ( .A1(n55), .A2(n69), .B1(n54), .B2(n50), .ZN(N298) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[10]), .ZN(n87) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[42]), .ZN(n51) );
  OAI22D1BWP30P140 U120 ( .A1(n55), .A2(n87), .B1(n54), .B2(n51), .ZN(N297) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[9]), .ZN(n70) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[41]), .ZN(n52) );
  OAI22D1BWP30P140 U123 ( .A1(n55), .A2(n70), .B1(n54), .B2(n52), .ZN(N296) );
  INVD1BWP30P140 U124 ( .I(i_data_bus[8]), .ZN(n90) );
  INVD1BWP30P140 U125 ( .I(i_data_bus[40]), .ZN(n53) );
  OAI22D1BWP30P140 U126 ( .A1(n55), .A2(n90), .B1(n54), .B2(n53), .ZN(N295) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n78), .B1(i_data_bus[39]), .B2(n88), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n78), .B1(i_data_bus[37]), .B2(n88), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n78), .B1(i_data_bus[35]), .B2(n88), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n78), .B1(i_data_bus[33]), .B2(n88), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n78), .B1(i_data_bus[38]), .B2(n88), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n78), .B1(i_data_bus[36]), .B2(n88), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n78), .B1(i_data_bus[34]), .B2(n88), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n78), .B1(i_data_bus[63]), .B2(n88), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n78), .B1(i_data_bus[61]), .B2(n88), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n78), .B1(i_data_bus[59]), .B2(n88), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n78), .B1(i_data_bus[57]), .B2(n88), 
        .ZN(N344) );
  INVD2BWP30P140 U138 ( .I(n67), .ZN(n89) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n89), .B1(i_data_bus[45]), .B2(n88), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n89), .B1(i_data_bus[43]), .B2(n88), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n89), .B1(i_data_bus[41]), .B2(n88), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n78), .B1(i_data_bus[62]), .B2(n88), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n78), .B1(i_data_bus[60]), .B2(n88), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n78), .B1(i_data_bus[58]), .B2(n88), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n78), .B1(i_data_bus[56]), .B2(n88), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n78), .B1(i_data_bus[55]), .B2(n88), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n78), .B1(i_data_bus[54]), .B2(n88), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n78), .B1(i_data_bus[53]), .B2(n88), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n78), .B1(i_data_bus[52]), .B2(n88), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n89), .B1(i_data_bus[51]), .B2(n88), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n89), .B1(i_data_bus[50]), .B2(n88), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n89), .B1(i_data_bus[49]), .B2(n88), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n89), .B1(i_data_bus[48]), .B2(n88), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n89), .B1(i_data_bus[47]), .B2(n88), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n89), .B1(i_data_bus[46]), .B2(n88), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n89), .B1(i_data_bus[44]), .B2(n88), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n89), .B1(i_data_bus[42]), .B2(n88), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U158 ( .A1(n90), .A2(n89), .B1(i_data_bus[40]), .B2(n88), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_11 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90;

  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  ND2OPTIBD1BWP30P140 U3 ( .A1(n9), .A2(n12), .ZN(n7) );
  INVD3BWP30P140 U4 ( .I(n67), .ZN(n78) );
  MOAI22D1BWP30P140 U5 ( .A1(n30), .A2(n78), .B1(i_data_bus[32]), .B2(n88), 
        .ZN(N319) );
  INVD1BWP30P140 U6 ( .I(n88), .ZN(n10) );
  INVD1BWP30P140 U7 ( .I(i_data_bus[0]), .ZN(n30) );
  INVD1BWP30P140 U8 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U9 ( .A1(n1), .A2(i_en), .ZN(n13) );
  NR2D1BWP30P140 U10 ( .A1(n13), .A2(i_cmd[1]), .ZN(n4) );
  INVD2BWP30P140 U11 ( .I(i_valid[0]), .ZN(n2) );
  INVD1BWP30P140 U12 ( .I(i_valid[1]), .ZN(n8) );
  MUX2NUD1BWP30P140 U13 ( .I0(n2), .I1(n8), .S(i_cmd[0]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U14 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U15 ( .I(n5), .ZN(n67) );
  INVD1BWP30P140 U16 ( .I(n13), .ZN(n6) );
  AN3D4BWP30P140 U17 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n6), .Z(n88) );
  INVD2BWP30P140 U18 ( .I(i_cmd[0]), .ZN(n12) );
  INR2D2BWP30P140 U19 ( .A1(i_valid[0]), .B1(n13), .ZN(n9) );
  INVD2BWP30P140 U20 ( .I(n7), .ZN(n32) );
  INVD2BWP30P140 U21 ( .I(n32), .ZN(n31) );
  OAI31D1BWP30P140 U22 ( .A1(n13), .A2(n8), .A3(n12), .B(n31), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n9), .ZN(n11) );
  OAI21D1BWP30P140 U24 ( .A1(n11), .A2(i_cmd[1]), .B(n10), .ZN(N354) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[19]), .ZN(n80) );
  MUX2NUD1BWP30P140 U26 ( .I0(n2), .I1(n8), .S(i_cmd[1]), .ZN(n15) );
  NR2D1BWP30P140 U27 ( .A1(n13), .A2(n12), .ZN(n14) );
  CKND2D2BWP30P140 U28 ( .A1(n15), .A2(n14), .ZN(n16) );
  INVD2BWP30P140 U29 ( .I(n16), .ZN(n18) );
  INVD2BWP30P140 U30 ( .I(n18), .ZN(n54) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[51]), .ZN(n17) );
  OAI22D1BWP30P140 U32 ( .A1(n31), .A2(n80), .B1(n54), .B2(n17), .ZN(N306) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD2BWP30P140 U34 ( .I(n18), .ZN(n42) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[52]), .ZN(n19) );
  OAI22D1BWP30P140 U36 ( .A1(n31), .A2(n79), .B1(n42), .B2(n19), .ZN(N307) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[21]), .ZN(n77) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[53]), .ZN(n20) );
  OAI22D1BWP30P140 U39 ( .A1(n31), .A2(n77), .B1(n42), .B2(n20), .ZN(N308) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[23]), .ZN(n75) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[55]), .ZN(n21) );
  OAI22D1BWP30P140 U42 ( .A1(n31), .A2(n75), .B1(n42), .B2(n21), .ZN(N310) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[25]), .ZN(n66) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[57]), .ZN(n22) );
  OAI22D1BWP30P140 U45 ( .A1(n31), .A2(n66), .B1(n42), .B2(n22), .ZN(N312) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[3]), .ZN(n58) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[35]), .ZN(n23) );
  OAI22D1BWP30P140 U48 ( .A1(n31), .A2(n58), .B1(n42), .B2(n23), .ZN(N290) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[27]), .ZN(n65) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[59]), .ZN(n24) );
  OAI22D1BWP30P140 U51 ( .A1(n31), .A2(n65), .B1(n42), .B2(n24), .ZN(N314) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[34]), .ZN(n25) );
  OAI22D1BWP30P140 U54 ( .A1(n31), .A2(n62), .B1(n54), .B2(n25), .ZN(N289) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[29]), .ZN(n64) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[61]), .ZN(n26) );
  OAI22D1BWP30P140 U57 ( .A1(n31), .A2(n64), .B1(n42), .B2(n26), .ZN(N316) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[33]), .ZN(n27) );
  OAI22D1BWP30P140 U60 ( .A1(n31), .A2(n59), .B1(n42), .B2(n27), .ZN(N288) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[31]), .ZN(n63) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[63]), .ZN(n28) );
  OAI22D1BWP30P140 U63 ( .A1(n31), .A2(n63), .B1(n42), .B2(n28), .ZN(N318) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[32]), .ZN(n29) );
  OAI22D1BWP30P140 U65 ( .A1(n31), .A2(n30), .B1(n54), .B2(n29), .ZN(N287) );
  INVD2BWP30P140 U66 ( .I(n32), .ZN(n55) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[39]), .ZN(n33) );
  OAI22D1BWP30P140 U69 ( .A1(n55), .A2(n56), .B1(n42), .B2(n33), .ZN(N294) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[6]), .ZN(n60) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[38]), .ZN(n34) );
  OAI22D1BWP30P140 U72 ( .A1(n55), .A2(n60), .B1(n54), .B2(n34), .ZN(N293) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[5]), .ZN(n57) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[37]), .ZN(n35) );
  OAI22D1BWP30P140 U75 ( .A1(n55), .A2(n57), .B1(n42), .B2(n35), .ZN(N292) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[36]), .ZN(n36) );
  OAI22D1BWP30P140 U78 ( .A1(n55), .A2(n61), .B1(n54), .B2(n36), .ZN(N291) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[30]), .ZN(n71) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[62]), .ZN(n37) );
  OAI22D1BWP30P140 U81 ( .A1(n55), .A2(n71), .B1(n42), .B2(n37), .ZN(N317) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[28]), .ZN(n72) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[60]), .ZN(n38) );
  OAI22D1BWP30P140 U84 ( .A1(n55), .A2(n72), .B1(n42), .B2(n38), .ZN(N315) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[26]), .ZN(n73) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[58]), .ZN(n39) );
  OAI22D1BWP30P140 U87 ( .A1(n55), .A2(n73), .B1(n42), .B2(n39), .ZN(N313) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[24]), .ZN(n74) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[56]), .ZN(n40) );
  OAI22D1BWP30P140 U90 ( .A1(n55), .A2(n74), .B1(n42), .B2(n40), .ZN(N311) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[22]), .ZN(n76) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[54]), .ZN(n41) );
  OAI22D1BWP30P140 U93 ( .A1(n55), .A2(n76), .B1(n42), .B2(n41), .ZN(N309) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[18]), .ZN(n81) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[50]), .ZN(n43) );
  OAI22D1BWP30P140 U96 ( .A1(n55), .A2(n81), .B1(n54), .B2(n43), .ZN(N305) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[17]), .ZN(n82) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[49]), .ZN(n44) );
  OAI22D1BWP30P140 U99 ( .A1(n55), .A2(n82), .B1(n54), .B2(n44), .ZN(N304) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[16]), .ZN(n83) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[48]), .ZN(n45) );
  OAI22D1BWP30P140 U102 ( .A1(n55), .A2(n83), .B1(n54), .B2(n45), .ZN(N303) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[15]), .ZN(n84) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[47]), .ZN(n46) );
  OAI22D1BWP30P140 U105 ( .A1(n55), .A2(n84), .B1(n54), .B2(n46), .ZN(N302) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[14]), .ZN(n85) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[46]), .ZN(n47) );
  OAI22D1BWP30P140 U108 ( .A1(n55), .A2(n85), .B1(n54), .B2(n47), .ZN(N301) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[13]), .ZN(n68) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[45]), .ZN(n48) );
  OAI22D1BWP30P140 U111 ( .A1(n55), .A2(n68), .B1(n54), .B2(n48), .ZN(N300) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[44]), .ZN(n49) );
  OAI22D1BWP30P140 U114 ( .A1(n55), .A2(n86), .B1(n54), .B2(n49), .ZN(N299) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[43]), .ZN(n50) );
  OAI22D1BWP30P140 U117 ( .A1(n55), .A2(n69), .B1(n54), .B2(n50), .ZN(N298) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[10]), .ZN(n87) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[42]), .ZN(n51) );
  OAI22D1BWP30P140 U120 ( .A1(n55), .A2(n87), .B1(n54), .B2(n51), .ZN(N297) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[9]), .ZN(n70) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[41]), .ZN(n52) );
  OAI22D1BWP30P140 U123 ( .A1(n55), .A2(n70), .B1(n54), .B2(n52), .ZN(N296) );
  INVD1BWP30P140 U124 ( .I(i_data_bus[8]), .ZN(n90) );
  INVD1BWP30P140 U125 ( .I(i_data_bus[40]), .ZN(n53) );
  OAI22D1BWP30P140 U126 ( .A1(n55), .A2(n90), .B1(n54), .B2(n53), .ZN(N295) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n78), .B1(i_data_bus[39]), .B2(n88), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n78), .B1(i_data_bus[37]), .B2(n88), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n78), .B1(i_data_bus[35]), .B2(n88), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n78), .B1(i_data_bus[33]), .B2(n88), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n78), .B1(i_data_bus[38]), .B2(n88), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n78), .B1(i_data_bus[36]), .B2(n88), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n78), .B1(i_data_bus[34]), .B2(n88), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n78), .B1(i_data_bus[63]), .B2(n88), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n78), .B1(i_data_bus[61]), .B2(n88), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n78), .B1(i_data_bus[59]), .B2(n88), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n78), .B1(i_data_bus[57]), .B2(n88), 
        .ZN(N344) );
  INVD2BWP30P140 U138 ( .I(n67), .ZN(n89) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n89), .B1(i_data_bus[45]), .B2(n88), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n89), .B1(i_data_bus[43]), .B2(n88), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n89), .B1(i_data_bus[41]), .B2(n88), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n78), .B1(i_data_bus[62]), .B2(n88), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n78), .B1(i_data_bus[60]), .B2(n88), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n78), .B1(i_data_bus[58]), .B2(n88), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n78), .B1(i_data_bus[56]), .B2(n88), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n78), .B1(i_data_bus[55]), .B2(n88), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n78), .B1(i_data_bus[54]), .B2(n88), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n78), .B1(i_data_bus[53]), .B2(n88), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n78), .B1(i_data_bus[52]), .B2(n88), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n89), .B1(i_data_bus[51]), .B2(n88), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n89), .B1(i_data_bus[50]), .B2(n88), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n89), .B1(i_data_bus[49]), .B2(n88), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n89), .B1(i_data_bus[48]), .B2(n88), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n89), .B1(i_data_bus[47]), .B2(n88), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n89), .B1(i_data_bus[46]), .B2(n88), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n89), .B1(i_data_bus[44]), .B2(n88), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n89), .B1(i_data_bus[42]), .B2(n88), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U158 ( .A1(n90), .A2(n89), .B1(i_data_bus[40]), .B2(n88), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_12 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90;

  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  ND2OPTIBD1BWP30P140 U3 ( .A1(n9), .A2(n12), .ZN(n7) );
  INVD3BWP30P140 U4 ( .I(n65), .ZN(n89) );
  MOAI22D1BWP30P140 U5 ( .A1(n39), .A2(n89), .B1(i_data_bus[39]), .B2(n88), 
        .ZN(N326) );
  INVD1BWP30P140 U6 ( .I(n88), .ZN(n10) );
  INVD1BWP30P140 U7 ( .I(i_data_bus[7]), .ZN(n39) );
  INVD1BWP30P140 U8 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U9 ( .A1(n1), .A2(i_en), .ZN(n13) );
  NR2D1BWP30P140 U10 ( .A1(n13), .A2(i_cmd[1]), .ZN(n4) );
  INVD2BWP30P140 U11 ( .I(i_valid[0]), .ZN(n2) );
  INVD1BWP30P140 U12 ( .I(i_valid[1]), .ZN(n8) );
  MUX2NUD1BWP30P140 U13 ( .I0(n2), .I1(n8), .S(i_cmd[0]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U14 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U15 ( .I(n5), .ZN(n65) );
  INVD1BWP30P140 U16 ( .I(n13), .ZN(n6) );
  AN3D4BWP30P140 U17 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n6), .Z(n88) );
  INVD2BWP30P140 U18 ( .I(i_cmd[0]), .ZN(n12) );
  INR2D2BWP30P140 U19 ( .A1(i_valid[0]), .B1(n13), .ZN(n9) );
  INVD2BWP30P140 U20 ( .I(n7), .ZN(n31) );
  INVD2BWP30P140 U21 ( .I(n31), .ZN(n30) );
  OAI31D1BWP30P140 U22 ( .A1(n13), .A2(n8), .A3(n12), .B(n30), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n9), .ZN(n11) );
  OAI21D1BWP30P140 U24 ( .A1(n11), .A2(i_cmd[1]), .B(n10), .ZN(N354) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[0]), .ZN(n56) );
  MUX2NUD1BWP30P140 U26 ( .I0(n2), .I1(n8), .S(i_cmd[1]), .ZN(n15) );
  NR2D1BWP30P140 U27 ( .A1(n13), .A2(n12), .ZN(n14) );
  CKND2D2BWP30P140 U28 ( .A1(n15), .A2(n14), .ZN(n16) );
  INVD2BWP30P140 U29 ( .I(n16), .ZN(n18) );
  INVD2BWP30P140 U30 ( .I(n18), .ZN(n54) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[32]), .ZN(n17) );
  OAI22D1BWP30P140 U32 ( .A1(n30), .A2(n56), .B1(n54), .B2(n17), .ZN(N287) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[27]), .ZN(n63) );
  INVD2BWP30P140 U34 ( .I(n18), .ZN(n48) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[59]), .ZN(n19) );
  OAI22D1BWP30P140 U36 ( .A1(n30), .A2(n63), .B1(n48), .B2(n19), .ZN(N314) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[29]), .ZN(n87) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[61]), .ZN(n20) );
  OAI22D1BWP30P140 U39 ( .A1(n30), .A2(n87), .B1(n48), .B2(n20), .ZN(N316) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[31]), .ZN(n90) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[63]), .ZN(n21) );
  OAI22D1BWP30P140 U42 ( .A1(n30), .A2(n90), .B1(n48), .B2(n21), .ZN(N318) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[1]), .ZN(n60) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[33]), .ZN(n22) );
  OAI22D1BWP30P140 U45 ( .A1(n30), .A2(n60), .B1(n48), .B2(n22), .ZN(N288) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[2]), .ZN(n57) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[34]), .ZN(n23) );
  OAI22D1BWP30P140 U48 ( .A1(n30), .A2(n57), .B1(n54), .B2(n23), .ZN(N289) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[35]), .ZN(n24) );
  OAI22D1BWP30P140 U51 ( .A1(n30), .A2(n61), .B1(n48), .B2(n24), .ZN(N290) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[19]), .ZN(n77) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[51]), .ZN(n25) );
  OAI22D1BWP30P140 U54 ( .A1(n30), .A2(n77), .B1(n54), .B2(n25), .ZN(N306) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[20]), .ZN(n76) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[52]), .ZN(n26) );
  OAI22D1BWP30P140 U57 ( .A1(n30), .A2(n76), .B1(n48), .B2(n26), .ZN(N307) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[21]), .ZN(n75) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[53]), .ZN(n27) );
  OAI22D1BWP30P140 U60 ( .A1(n30), .A2(n75), .B1(n48), .B2(n27), .ZN(N308) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[23]), .ZN(n73) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[55]), .ZN(n28) );
  OAI22D1BWP30P140 U63 ( .A1(n30), .A2(n73), .B1(n48), .B2(n28), .ZN(N310) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[25]), .ZN(n64) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[57]), .ZN(n29) );
  OAI22D1BWP30P140 U66 ( .A1(n30), .A2(n64), .B1(n48), .B2(n29), .ZN(N312) );
  INVD2BWP30P140 U67 ( .I(n31), .ZN(n55) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[24]), .ZN(n72) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[56]), .ZN(n32) );
  OAI22D1BWP30P140 U70 ( .A1(n55), .A2(n72), .B1(n48), .B2(n32), .ZN(N311) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[54]), .ZN(n33) );
  OAI22D1BWP30P140 U73 ( .A1(n55), .A2(n74), .B1(n48), .B2(n33), .ZN(N309) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[18]), .ZN(n78) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[50]), .ZN(n34) );
  OAI22D1BWP30P140 U76 ( .A1(n55), .A2(n78), .B1(n54), .B2(n34), .ZN(N305) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[9]), .ZN(n68) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[41]), .ZN(n35) );
  OAI22D1BWP30P140 U79 ( .A1(n55), .A2(n68), .B1(n54), .B2(n35), .ZN(N296) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[12]), .ZN(n83) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[44]), .ZN(n36) );
  OAI22D1BWP30P140 U82 ( .A1(n55), .A2(n83), .B1(n54), .B2(n36), .ZN(N299) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[11]), .ZN(n67) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[43]), .ZN(n37) );
  OAI22D1BWP30P140 U85 ( .A1(n55), .A2(n67), .B1(n54), .B2(n37), .ZN(N298) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[39]), .ZN(n38) );
  OAI22D1BWP30P140 U87 ( .A1(n55), .A2(n39), .B1(n48), .B2(n38), .ZN(N294) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[6]), .ZN(n59) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[38]), .ZN(n40) );
  OAI22D1BWP30P140 U90 ( .A1(n55), .A2(n59), .B1(n54), .B2(n40), .ZN(N293) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[4]), .ZN(n58) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[36]), .ZN(n41) );
  OAI22D1BWP30P140 U93 ( .A1(n55), .A2(n58), .B1(n54), .B2(n41), .ZN(N291) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n69) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[62]), .ZN(n42) );
  OAI22D1BWP30P140 U96 ( .A1(n55), .A2(n69), .B1(n48), .B2(n42), .ZN(N317) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[28]), .ZN(n70) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[60]), .ZN(n43) );
  OAI22D1BWP30P140 U99 ( .A1(n55), .A2(n70), .B1(n48), .B2(n43), .ZN(N315) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[8]), .ZN(n86) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[40]), .ZN(n44) );
  OAI22D1BWP30P140 U102 ( .A1(n55), .A2(n86), .B1(n54), .B2(n44), .ZN(N295) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[13]), .ZN(n66) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[45]), .ZN(n45) );
  OAI22D1BWP30P140 U105 ( .A1(n55), .A2(n66), .B1(n54), .B2(n45), .ZN(N300) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[26]), .ZN(n71) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[58]), .ZN(n46) );
  OAI22D1BWP30P140 U108 ( .A1(n55), .A2(n71), .B1(n48), .B2(n46), .ZN(N313) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[37]), .ZN(n47) );
  OAI22D1BWP30P140 U111 ( .A1(n55), .A2(n62), .B1(n48), .B2(n47), .ZN(N292) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[10]), .ZN(n84) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[42]), .ZN(n49) );
  OAI22D1BWP30P140 U114 ( .A1(n55), .A2(n84), .B1(n54), .B2(n49), .ZN(N297) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[15]), .ZN(n81) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[47]), .ZN(n50) );
  OAI22D1BWP30P140 U117 ( .A1(n55), .A2(n81), .B1(n54), .B2(n50), .ZN(N302) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[17]), .ZN(n79) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[49]), .ZN(n51) );
  OAI22D1BWP30P140 U120 ( .A1(n55), .A2(n79), .B1(n54), .B2(n51), .ZN(N304) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[14]), .ZN(n82) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[46]), .ZN(n52) );
  OAI22D1BWP30P140 U123 ( .A1(n55), .A2(n82), .B1(n54), .B2(n52), .ZN(N301) );
  INVD1BWP30P140 U124 ( .I(i_data_bus[16]), .ZN(n80) );
  INVD1BWP30P140 U125 ( .I(i_data_bus[48]), .ZN(n53) );
  OAI22D1BWP30P140 U126 ( .A1(n55), .A2(n80), .B1(n54), .B2(n53), .ZN(N303) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n89), .B1(i_data_bus[32]), .B2(n88), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n89), .B1(i_data_bus[34]), .B2(n88), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n89), .B1(i_data_bus[36]), .B2(n88), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n89), .B1(i_data_bus[38]), .B2(n88), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n89), .B1(i_data_bus[33]), .B2(n88), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n89), .B1(i_data_bus[35]), .B2(n88), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n89), .B1(i_data_bus[37]), .B2(n88), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n89), .B1(i_data_bus[59]), .B2(n88), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n89), .B1(i_data_bus[57]), .B2(n88), 
        .ZN(N344) );
  INVD2BWP30P140 U136 ( .I(n65), .ZN(n85) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n85), .B1(i_data_bus[45]), .B2(n88), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n85), .B1(i_data_bus[43]), .B2(n88), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n85), .B1(i_data_bus[41]), .B2(n88), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n89), .B1(i_data_bus[62]), .B2(n88), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n89), .B1(i_data_bus[60]), .B2(n88), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n89), .B1(i_data_bus[58]), .B2(n88), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n89), .B1(i_data_bus[56]), .B2(n88), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n89), .B1(i_data_bus[55]), .B2(n88), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n89), .B1(i_data_bus[54]), .B2(n88), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n89), .B1(i_data_bus[53]), .B2(n88), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n89), .B1(i_data_bus[52]), .B2(n88), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n85), .B1(i_data_bus[51]), .B2(n88), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n85), .B1(i_data_bus[50]), .B2(n88), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n85), .B1(i_data_bus[49]), .B2(n88), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n85), .B1(i_data_bus[48]), .B2(n88), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n85), .B1(i_data_bus[47]), .B2(n88), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n85), .B1(i_data_bus[46]), .B2(n88), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n85), .B1(i_data_bus[44]), .B2(n88), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n85), .B1(i_data_bus[42]), .B2(n88), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n85), .B1(i_data_bus[40]), .B2(n88), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n89), .B1(i_data_bus[61]), .B2(n88), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U158 ( .A1(n90), .A2(n89), .B1(i_data_bus[63]), .B2(n88), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_13 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90;

  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  ND2OPTIBD1BWP30P140 U3 ( .A1(n9), .A2(n12), .ZN(n7) );
  INVD3BWP30P140 U4 ( .I(n67), .ZN(n78) );
  MOAI22D1BWP30P140 U5 ( .A1(n49), .A2(n78), .B1(i_data_bus[36]), .B2(n88), 
        .ZN(N323) );
  INVD1BWP30P140 U6 ( .I(n88), .ZN(n10) );
  INVD1BWP30P140 U7 ( .I(i_data_bus[4]), .ZN(n49) );
  INVD1BWP30P140 U8 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U9 ( .A1(n1), .A2(i_en), .ZN(n13) );
  NR2D1BWP30P140 U10 ( .A1(n13), .A2(i_cmd[1]), .ZN(n4) );
  INVD2BWP30P140 U11 ( .I(i_valid[0]), .ZN(n2) );
  INVD1BWP30P140 U12 ( .I(i_valid[1]), .ZN(n8) );
  MUX2NUD1BWP30P140 U13 ( .I0(n2), .I1(n8), .S(i_cmd[0]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U14 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U15 ( .I(n5), .ZN(n67) );
  INVD1BWP30P140 U16 ( .I(n13), .ZN(n6) );
  AN3D4BWP30P140 U17 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n6), .Z(n88) );
  INVD2BWP30P140 U18 ( .I(i_cmd[0]), .ZN(n12) );
  INR2D2BWP30P140 U19 ( .A1(i_valid[0]), .B1(n13), .ZN(n9) );
  INVD2BWP30P140 U20 ( .I(n7), .ZN(n31) );
  INVD2BWP30P140 U21 ( .I(n31), .ZN(n30) );
  OAI31D1BWP30P140 U22 ( .A1(n13), .A2(n8), .A3(n12), .B(n30), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n9), .ZN(n11) );
  OAI21D1BWP30P140 U24 ( .A1(n11), .A2(i_cmd[1]), .B(n10), .ZN(N354) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[3]), .ZN(n58) );
  MUX2NUD1BWP30P140 U26 ( .I0(n2), .I1(n8), .S(i_cmd[1]), .ZN(n15) );
  NR2D1BWP30P140 U27 ( .A1(n13), .A2(n12), .ZN(n14) );
  CKND2D2BWP30P140 U28 ( .A1(n15), .A2(n14), .ZN(n16) );
  INVD2BWP30P140 U29 ( .I(n16), .ZN(n18) );
  INVD2BWP30P140 U30 ( .I(n18), .ZN(n54) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[35]), .ZN(n17) );
  OAI22D1BWP30P140 U32 ( .A1(n30), .A2(n58), .B1(n54), .B2(n17), .ZN(N290) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD2BWP30P140 U34 ( .I(n18), .ZN(n52) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[34]), .ZN(n19) );
  OAI22D1BWP30P140 U36 ( .A1(n30), .A2(n62), .B1(n52), .B2(n19), .ZN(N289) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[1]), .ZN(n57) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[33]), .ZN(n20) );
  OAI22D1BWP30P140 U39 ( .A1(n30), .A2(n57), .B1(n54), .B2(n20), .ZN(N288) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[0]), .ZN(n61) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[32]), .ZN(n21) );
  OAI22D1BWP30P140 U42 ( .A1(n30), .A2(n61), .B1(n52), .B2(n21), .ZN(N287) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[31]), .ZN(n63) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[63]), .ZN(n22) );
  OAI22D1BWP30P140 U45 ( .A1(n30), .A2(n63), .B1(n54), .B2(n22), .ZN(N318) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[29]), .ZN(n64) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[61]), .ZN(n23) );
  OAI22D1BWP30P140 U48 ( .A1(n30), .A2(n64), .B1(n54), .B2(n23), .ZN(N316) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[27]), .ZN(n65) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[59]), .ZN(n24) );
  OAI22D1BWP30P140 U51 ( .A1(n30), .A2(n65), .B1(n54), .B2(n24), .ZN(N314) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[25]), .ZN(n66) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[57]), .ZN(n25) );
  OAI22D1BWP30P140 U54 ( .A1(n30), .A2(n66), .B1(n54), .B2(n25), .ZN(N312) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[23]), .ZN(n75) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[55]), .ZN(n26) );
  OAI22D1BWP30P140 U57 ( .A1(n30), .A2(n75), .B1(n54), .B2(n26), .ZN(N310) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[21]), .ZN(n77) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[53]), .ZN(n27) );
  OAI22D1BWP30P140 U60 ( .A1(n30), .A2(n77), .B1(n54), .B2(n27), .ZN(N308) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[52]), .ZN(n28) );
  OAI22D1BWP30P140 U63 ( .A1(n30), .A2(n79), .B1(n54), .B2(n28), .ZN(N307) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[19]), .ZN(n80) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[51]), .ZN(n29) );
  OAI22D1BWP30P140 U66 ( .A1(n30), .A2(n80), .B1(n52), .B2(n29), .ZN(N306) );
  INVD2BWP30P140 U67 ( .I(n31), .ZN(n55) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[8]), .ZN(n90) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[40]), .ZN(n32) );
  OAI22D1BWP30P140 U70 ( .A1(n55), .A2(n90), .B1(n52), .B2(n32), .ZN(N295) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[9]), .ZN(n70) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[41]), .ZN(n33) );
  OAI22D1BWP30P140 U73 ( .A1(n55), .A2(n70), .B1(n52), .B2(n33), .ZN(N296) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[10]), .ZN(n87) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[42]), .ZN(n34) );
  OAI22D1BWP30P140 U76 ( .A1(n55), .A2(n87), .B1(n52), .B2(n34), .ZN(N297) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[43]), .ZN(n35) );
  OAI22D1BWP30P140 U79 ( .A1(n55), .A2(n69), .B1(n52), .B2(n35), .ZN(N298) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[44]), .ZN(n36) );
  OAI22D1BWP30P140 U82 ( .A1(n55), .A2(n86), .B1(n52), .B2(n36), .ZN(N299) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[13]), .ZN(n68) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[45]), .ZN(n37) );
  OAI22D1BWP30P140 U85 ( .A1(n55), .A2(n68), .B1(n52), .B2(n37), .ZN(N300) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[14]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[46]), .ZN(n38) );
  OAI22D1BWP30P140 U88 ( .A1(n55), .A2(n85), .B1(n52), .B2(n38), .ZN(N301) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[15]), .ZN(n84) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[47]), .ZN(n39) );
  OAI22D1BWP30P140 U91 ( .A1(n55), .A2(n84), .B1(n52), .B2(n39), .ZN(N302) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[16]), .ZN(n83) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[48]), .ZN(n40) );
  OAI22D1BWP30P140 U94 ( .A1(n55), .A2(n83), .B1(n52), .B2(n40), .ZN(N303) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[17]), .ZN(n82) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[49]), .ZN(n41) );
  OAI22D1BWP30P140 U97 ( .A1(n55), .A2(n82), .B1(n52), .B2(n41), .ZN(N304) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[18]), .ZN(n81) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[50]), .ZN(n42) );
  OAI22D1BWP30P140 U100 ( .A1(n55), .A2(n81), .B1(n52), .B2(n42), .ZN(N305) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[22]), .ZN(n76) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[54]), .ZN(n43) );
  OAI22D1BWP30P140 U103 ( .A1(n55), .A2(n76), .B1(n54), .B2(n43), .ZN(N309) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[24]), .ZN(n74) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[56]), .ZN(n44) );
  OAI22D1BWP30P140 U106 ( .A1(n55), .A2(n74), .B1(n54), .B2(n44), .ZN(N311) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[26]), .ZN(n73) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[58]), .ZN(n45) );
  OAI22D1BWP30P140 U109 ( .A1(n55), .A2(n73), .B1(n54), .B2(n45), .ZN(N313) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[28]), .ZN(n72) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[60]), .ZN(n46) );
  OAI22D1BWP30P140 U112 ( .A1(n55), .A2(n72), .B1(n54), .B2(n46), .ZN(N315) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[30]), .ZN(n71) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[62]), .ZN(n47) );
  OAI22D1BWP30P140 U115 ( .A1(n55), .A2(n71), .B1(n54), .B2(n47), .ZN(N317) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[36]), .ZN(n48) );
  OAI22D1BWP30P140 U117 ( .A1(n55), .A2(n49), .B1(n52), .B2(n48), .ZN(N291) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[37]), .ZN(n50) );
  OAI22D1BWP30P140 U120 ( .A1(n55), .A2(n59), .B1(n54), .B2(n50), .ZN(N292) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[6]), .ZN(n56) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[38]), .ZN(n51) );
  OAI22D1BWP30P140 U123 ( .A1(n55), .A2(n56), .B1(n52), .B2(n51), .ZN(N293) );
  INVD1BWP30P140 U124 ( .I(i_data_bus[7]), .ZN(n60) );
  INVD1BWP30P140 U125 ( .I(i_data_bus[39]), .ZN(n53) );
  OAI22D1BWP30P140 U126 ( .A1(n55), .A2(n60), .B1(n54), .B2(n53), .ZN(N294) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n78), .B1(i_data_bus[38]), .B2(n88), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n78), .B1(i_data_bus[33]), .B2(n88), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n78), .B1(i_data_bus[35]), .B2(n88), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n78), .B1(i_data_bus[37]), .B2(n88), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n78), .B1(i_data_bus[39]), .B2(n88), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n78), .B1(i_data_bus[32]), .B2(n88), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n78), .B1(i_data_bus[34]), .B2(n88), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n78), .B1(i_data_bus[63]), .B2(n88), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n78), .B1(i_data_bus[61]), .B2(n88), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n78), .B1(i_data_bus[59]), .B2(n88), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n78), .B1(i_data_bus[57]), .B2(n88), 
        .ZN(N344) );
  INVD2BWP30P140 U138 ( .I(n67), .ZN(n89) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n89), .B1(i_data_bus[45]), .B2(n88), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n89), .B1(i_data_bus[43]), .B2(n88), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n89), .B1(i_data_bus[41]), .B2(n88), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n78), .B1(i_data_bus[62]), .B2(n88), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n78), .B1(i_data_bus[60]), .B2(n88), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n78), .B1(i_data_bus[58]), .B2(n88), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n78), .B1(i_data_bus[56]), .B2(n88), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n78), .B1(i_data_bus[55]), .B2(n88), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n78), .B1(i_data_bus[54]), .B2(n88), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n78), .B1(i_data_bus[53]), .B2(n88), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n78), .B1(i_data_bus[52]), .B2(n88), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n89), .B1(i_data_bus[51]), .B2(n88), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n89), .B1(i_data_bus[50]), .B2(n88), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n89), .B1(i_data_bus[49]), .B2(n88), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n89), .B1(i_data_bus[48]), .B2(n88), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n89), .B1(i_data_bus[47]), .B2(n88), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n89), .B1(i_data_bus[46]), .B2(n88), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n89), .B1(i_data_bus[44]), .B2(n88), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n89), .B1(i_data_bus[42]), .B2(n88), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U158 ( .A1(n90), .A2(n89), .B1(i_data_bus[40]), .B2(n88), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_14 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90;

  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  ND2OPTIBD1BWP30P140 U3 ( .A1(n9), .A2(n12), .ZN(n7) );
  INVD3BWP30P140 U4 ( .I(n72), .ZN(n83) );
  MOAI22D1BWP30P140 U5 ( .A1(n21), .A2(n83), .B1(i_data_bus[33]), .B2(n88), 
        .ZN(N320) );
  INVD1BWP30P140 U6 ( .I(n88), .ZN(n10) );
  INVD1BWP30P140 U7 ( .I(i_data_bus[1]), .ZN(n21) );
  INVD1BWP30P140 U8 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U9 ( .A1(n1), .A2(i_en), .ZN(n13) );
  NR2D1BWP30P140 U10 ( .A1(n13), .A2(i_cmd[1]), .ZN(n4) );
  INVD2BWP30P140 U11 ( .I(i_valid[0]), .ZN(n2) );
  INVD1BWP30P140 U12 ( .I(i_valid[1]), .ZN(n8) );
  MUX2NUD1BWP30P140 U13 ( .I0(n2), .I1(n8), .S(i_cmd[0]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U14 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U15 ( .I(n5), .ZN(n72) );
  INVD1BWP30P140 U16 ( .I(n13), .ZN(n6) );
  AN3D4BWP30P140 U17 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n6), .Z(n88) );
  INVD2BWP30P140 U18 ( .I(i_cmd[0]), .ZN(n12) );
  INR2D2BWP30P140 U19 ( .A1(i_valid[0]), .B1(n13), .ZN(n9) );
  INVD2BWP30P140 U20 ( .I(n7), .ZN(n32) );
  INVD2BWP30P140 U21 ( .I(n32), .ZN(n31) );
  OAI31D1BWP30P140 U22 ( .A1(n13), .A2(n8), .A3(n12), .B(n31), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n9), .ZN(n11) );
  OAI21D1BWP30P140 U24 ( .A1(n11), .A2(i_cmd[1]), .B(n10), .ZN(N354) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[3]), .ZN(n62) );
  MUX2NUD1BWP30P140 U26 ( .I0(n2), .I1(n8), .S(i_cmd[1]), .ZN(n15) );
  NR2D1BWP30P140 U27 ( .A1(n13), .A2(n12), .ZN(n14) );
  CKND2D2BWP30P140 U28 ( .A1(n15), .A2(n14), .ZN(n16) );
  INVD2BWP30P140 U29 ( .I(n16), .ZN(n18) );
  INVD2BWP30P140 U30 ( .I(n18), .ZN(n54) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[35]), .ZN(n17) );
  OAI22D1BWP30P140 U32 ( .A1(n31), .A2(n62), .B1(n54), .B2(n17), .ZN(N290) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[2]), .ZN(n58) );
  INVD2BWP30P140 U34 ( .I(n18), .ZN(n52) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[34]), .ZN(n19) );
  OAI22D1BWP30P140 U36 ( .A1(n31), .A2(n58), .B1(n52), .B2(n19), .ZN(N289) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[33]), .ZN(n20) );
  OAI22D1BWP30P140 U38 ( .A1(n31), .A2(n21), .B1(n54), .B2(n20), .ZN(N288) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[0]), .ZN(n59) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[32]), .ZN(n22) );
  OAI22D1BWP30P140 U41 ( .A1(n31), .A2(n59), .B1(n52), .B2(n22), .ZN(N287) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[31]), .ZN(n90) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[63]), .ZN(n23) );
  OAI22D1BWP30P140 U44 ( .A1(n31), .A2(n90), .B1(n54), .B2(n23), .ZN(N318) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[29]), .ZN(n87) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[61]), .ZN(n24) );
  OAI22D1BWP30P140 U47 ( .A1(n31), .A2(n87), .B1(n54), .B2(n24), .ZN(N316) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[59]), .ZN(n25) );
  OAI22D1BWP30P140 U50 ( .A1(n31), .A2(n86), .B1(n54), .B2(n25), .ZN(N314) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[25]), .ZN(n85) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[57]), .ZN(n26) );
  OAI22D1BWP30P140 U53 ( .A1(n31), .A2(n85), .B1(n54), .B2(n26), .ZN(N312) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[23]), .ZN(n76) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[55]), .ZN(n27) );
  OAI22D1BWP30P140 U56 ( .A1(n31), .A2(n76), .B1(n54), .B2(n27), .ZN(N310) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[21]), .ZN(n74) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[53]), .ZN(n28) );
  OAI22D1BWP30P140 U59 ( .A1(n31), .A2(n74), .B1(n54), .B2(n28), .ZN(N308) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[20]), .ZN(n73) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[52]), .ZN(n29) );
  OAI22D1BWP30P140 U62 ( .A1(n31), .A2(n73), .B1(n54), .B2(n29), .ZN(N307) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[19]), .ZN(n71) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[51]), .ZN(n30) );
  OAI22D1BWP30P140 U65 ( .A1(n31), .A2(n71), .B1(n52), .B2(n30), .ZN(N306) );
  INVD2BWP30P140 U66 ( .I(n32), .ZN(n55) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[8]), .ZN(n63) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[40]), .ZN(n33) );
  OAI22D1BWP30P140 U69 ( .A1(n55), .A2(n63), .B1(n52), .B2(n33), .ZN(N295) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[9]), .ZN(n81) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[41]), .ZN(n34) );
  OAI22D1BWP30P140 U72 ( .A1(n55), .A2(n81), .B1(n52), .B2(n34), .ZN(N296) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[10]), .ZN(n64) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[42]), .ZN(n35) );
  OAI22D1BWP30P140 U75 ( .A1(n55), .A2(n64), .B1(n52), .B2(n35), .ZN(N297) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[11]), .ZN(n82) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[43]), .ZN(n36) );
  OAI22D1BWP30P140 U78 ( .A1(n55), .A2(n82), .B1(n52), .B2(n36), .ZN(N298) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[12]), .ZN(n65) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[44]), .ZN(n37) );
  OAI22D1BWP30P140 U81 ( .A1(n55), .A2(n65), .B1(n52), .B2(n37), .ZN(N299) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[13]), .ZN(n84) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[45]), .ZN(n38) );
  OAI22D1BWP30P140 U84 ( .A1(n55), .A2(n84), .B1(n52), .B2(n38), .ZN(N300) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[14]), .ZN(n66) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[46]), .ZN(n39) );
  OAI22D1BWP30P140 U87 ( .A1(n55), .A2(n66), .B1(n52), .B2(n39), .ZN(N301) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[15]), .ZN(n67) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[47]), .ZN(n40) );
  OAI22D1BWP30P140 U90 ( .A1(n55), .A2(n67), .B1(n52), .B2(n40), .ZN(N302) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[16]), .ZN(n68) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[48]), .ZN(n41) );
  OAI22D1BWP30P140 U93 ( .A1(n55), .A2(n68), .B1(n52), .B2(n41), .ZN(N303) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[17]), .ZN(n69) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[49]), .ZN(n42) );
  OAI22D1BWP30P140 U96 ( .A1(n55), .A2(n69), .B1(n52), .B2(n42), .ZN(N304) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[18]), .ZN(n70) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[50]), .ZN(n43) );
  OAI22D1BWP30P140 U99 ( .A1(n55), .A2(n70), .B1(n52), .B2(n43), .ZN(N305) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[22]), .ZN(n75) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[54]), .ZN(n44) );
  OAI22D1BWP30P140 U102 ( .A1(n55), .A2(n75), .B1(n54), .B2(n44), .ZN(N309) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[24]), .ZN(n77) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[56]), .ZN(n45) );
  OAI22D1BWP30P140 U105 ( .A1(n55), .A2(n77), .B1(n54), .B2(n45), .ZN(N311) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[26]), .ZN(n78) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[58]), .ZN(n46) );
  OAI22D1BWP30P140 U108 ( .A1(n55), .A2(n78), .B1(n54), .B2(n46), .ZN(N313) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[28]), .ZN(n79) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[60]), .ZN(n47) );
  OAI22D1BWP30P140 U111 ( .A1(n55), .A2(n79), .B1(n54), .B2(n47), .ZN(N315) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[30]), .ZN(n80) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[62]), .ZN(n48) );
  OAI22D1BWP30P140 U114 ( .A1(n55), .A2(n80), .B1(n54), .B2(n48), .ZN(N317) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[4]), .ZN(n57) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[36]), .ZN(n49) );
  OAI22D1BWP30P140 U117 ( .A1(n55), .A2(n57), .B1(n52), .B2(n49), .ZN(N291) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[5]), .ZN(n61) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[37]), .ZN(n50) );
  OAI22D1BWP30P140 U120 ( .A1(n55), .A2(n61), .B1(n54), .B2(n50), .ZN(N292) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[6]), .ZN(n56) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[38]), .ZN(n51) );
  OAI22D1BWP30P140 U123 ( .A1(n55), .A2(n56), .B1(n52), .B2(n51), .ZN(N293) );
  INVD1BWP30P140 U124 ( .I(i_data_bus[7]), .ZN(n60) );
  INVD1BWP30P140 U125 ( .I(i_data_bus[39]), .ZN(n53) );
  OAI22D1BWP30P140 U126 ( .A1(n55), .A2(n60), .B1(n54), .B2(n53), .ZN(N294) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n83), .B1(i_data_bus[38]), .B2(n88), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n83), .B1(i_data_bus[36]), .B2(n88), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n83), .B1(i_data_bus[34]), .B2(n88), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n83), .B1(i_data_bus[32]), .B2(n88), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n83), .B1(i_data_bus[39]), .B2(n88), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n83), .B1(i_data_bus[37]), .B2(n88), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n83), .B1(i_data_bus[35]), .B2(n88), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n83), .B1(i_data_bus[40]), .B2(n88), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n83), .B1(i_data_bus[42]), .B2(n88), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n83), .B1(i_data_bus[44]), .B2(n88), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n83), .B1(i_data_bus[46]), .B2(n88), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n83), .B1(i_data_bus[47]), .B2(n88), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n83), .B1(i_data_bus[48]), .B2(n88), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n83), .B1(i_data_bus[49]), .B2(n88), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n83), .B1(i_data_bus[50]), .B2(n88), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n83), .B1(i_data_bus[51]), .B2(n88), 
        .ZN(N338) );
  INVD2BWP30P140 U143 ( .I(n72), .ZN(n89) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n89), .B1(i_data_bus[52]), .B2(n88), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n89), .B1(i_data_bus[53]), .B2(n88), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n89), .B1(i_data_bus[54]), .B2(n88), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n89), .B1(i_data_bus[55]), .B2(n88), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n89), .B1(i_data_bus[56]), .B2(n88), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n89), .B1(i_data_bus[58]), .B2(n88), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n89), .B1(i_data_bus[60]), .B2(n88), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n89), .B1(i_data_bus[62]), .B2(n88), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n83), .B1(i_data_bus[41]), .B2(n88), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n83), .B1(i_data_bus[43]), .B2(n88), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n83), .B1(i_data_bus[45]), .B2(n88), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n89), .B1(i_data_bus[57]), .B2(n88), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n89), .B1(i_data_bus[59]), .B2(n88), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n89), .B1(i_data_bus[61]), .B2(n88), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U158 ( .A1(n90), .A2(n89), .B1(i_data_bus[63]), .B2(n88), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_15 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90;

  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  ND2OPTIBD1BWP30P140 U3 ( .A1(n9), .A2(n12), .ZN(n7) );
  INVD3BWP30P140 U4 ( .I(n72), .ZN(n83) );
  MOAI22D1BWP30P140 U5 ( .A1(n54), .A2(n83), .B1(i_data_bus[39]), .B2(n88), 
        .ZN(N326) );
  INVD1BWP30P140 U6 ( .I(n88), .ZN(n10) );
  INVD1BWP30P140 U7 ( .I(i_data_bus[7]), .ZN(n54) );
  INVD1BWP30P140 U8 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U9 ( .A1(n1), .A2(i_en), .ZN(n13) );
  NR2D1BWP30P140 U10 ( .A1(n13), .A2(i_cmd[1]), .ZN(n4) );
  INVD2BWP30P140 U11 ( .I(i_valid[0]), .ZN(n2) );
  INVD1BWP30P140 U12 ( .I(i_valid[1]), .ZN(n8) );
  MUX2NUD1BWP30P140 U13 ( .I0(n2), .I1(n8), .S(i_cmd[0]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U14 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U15 ( .I(n5), .ZN(n72) );
  INVD1BWP30P140 U16 ( .I(n13), .ZN(n6) );
  AN3D4BWP30P140 U17 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n6), .Z(n88) );
  INVD2BWP30P140 U18 ( .I(i_cmd[0]), .ZN(n12) );
  INR2D2BWP30P140 U19 ( .A1(i_valid[0]), .B1(n13), .ZN(n9) );
  INVD2BWP30P140 U20 ( .I(n7), .ZN(n31) );
  INVD2BWP30P140 U21 ( .I(n31), .ZN(n30) );
  OAI31D1BWP30P140 U22 ( .A1(n13), .A2(n8), .A3(n12), .B(n30), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n9), .ZN(n11) );
  OAI21D1BWP30P140 U24 ( .A1(n11), .A2(i_cmd[1]), .B(n10), .ZN(N354) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[20]), .ZN(n73) );
  MUX2NUD1BWP30P140 U26 ( .I0(n2), .I1(n8), .S(i_cmd[1]), .ZN(n15) );
  NR2D1BWP30P140 U27 ( .A1(n13), .A2(n12), .ZN(n14) );
  CKND2D2BWP30P140 U28 ( .A1(n15), .A2(n14), .ZN(n16) );
  INVD2BWP30P140 U29 ( .I(n16), .ZN(n18) );
  INVD2BWP30P140 U30 ( .I(n18), .ZN(n53) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[52]), .ZN(n17) );
  OAI22D1BWP30P140 U32 ( .A1(n30), .A2(n73), .B1(n53), .B2(n17), .ZN(N307) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[19]), .ZN(n71) );
  INVD2BWP30P140 U34 ( .I(n18), .ZN(n51) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[51]), .ZN(n19) );
  OAI22D1BWP30P140 U36 ( .A1(n30), .A2(n71), .B1(n51), .B2(n19), .ZN(N306) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[1]), .ZN(n60) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[33]), .ZN(n20) );
  OAI22D1BWP30P140 U39 ( .A1(n30), .A2(n60), .B1(n53), .B2(n20), .ZN(N288) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[23]), .ZN(n76) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[55]), .ZN(n21) );
  OAI22D1BWP30P140 U42 ( .A1(n30), .A2(n76), .B1(n53), .B2(n21), .ZN(N310) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[35]), .ZN(n22) );
  OAI22D1BWP30P140 U45 ( .A1(n30), .A2(n61), .B1(n53), .B2(n22), .ZN(N290) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[2]), .ZN(n57) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[34]), .ZN(n23) );
  OAI22D1BWP30P140 U48 ( .A1(n30), .A2(n57), .B1(n51), .B2(n23), .ZN(N289) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[29]), .ZN(n87) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[61]), .ZN(n24) );
  OAI22D1BWP30P140 U51 ( .A1(n30), .A2(n87), .B1(n53), .B2(n24), .ZN(N316) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[31]), .ZN(n90) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[63]), .ZN(n25) );
  OAI22D1BWP30P140 U54 ( .A1(n30), .A2(n90), .B1(n53), .B2(n25), .ZN(N318) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[59]), .ZN(n26) );
  OAI22D1BWP30P140 U57 ( .A1(n30), .A2(n86), .B1(n53), .B2(n26), .ZN(N314) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[25]), .ZN(n85) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[57]), .ZN(n27) );
  OAI22D1BWP30P140 U60 ( .A1(n30), .A2(n85), .B1(n53), .B2(n27), .ZN(N312) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[21]), .ZN(n74) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[53]), .ZN(n28) );
  OAI22D1BWP30P140 U63 ( .A1(n30), .A2(n74), .B1(n53), .B2(n28), .ZN(N308) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[0]), .ZN(n56) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[32]), .ZN(n29) );
  OAI22D1BWP30P140 U66 ( .A1(n30), .A2(n56), .B1(n51), .B2(n29), .ZN(N287) );
  INVD2BWP30P140 U67 ( .I(n31), .ZN(n55) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[8]), .ZN(n63) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[40]), .ZN(n32) );
  OAI22D1BWP30P140 U70 ( .A1(n55), .A2(n63), .B1(n51), .B2(n32), .ZN(N295) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[9]), .ZN(n81) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[41]), .ZN(n33) );
  OAI22D1BWP30P140 U73 ( .A1(n55), .A2(n81), .B1(n51), .B2(n33), .ZN(N296) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[10]), .ZN(n64) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[42]), .ZN(n34) );
  OAI22D1BWP30P140 U76 ( .A1(n55), .A2(n64), .B1(n51), .B2(n34), .ZN(N297) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[11]), .ZN(n82) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[43]), .ZN(n35) );
  OAI22D1BWP30P140 U79 ( .A1(n55), .A2(n82), .B1(n51), .B2(n35), .ZN(N298) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[12]), .ZN(n65) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[44]), .ZN(n36) );
  OAI22D1BWP30P140 U82 ( .A1(n55), .A2(n65), .B1(n51), .B2(n36), .ZN(N299) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[13]), .ZN(n84) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[45]), .ZN(n37) );
  OAI22D1BWP30P140 U85 ( .A1(n55), .A2(n84), .B1(n51), .B2(n37), .ZN(N300) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[14]), .ZN(n66) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[46]), .ZN(n38) );
  OAI22D1BWP30P140 U88 ( .A1(n55), .A2(n66), .B1(n51), .B2(n38), .ZN(N301) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[15]), .ZN(n67) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[47]), .ZN(n39) );
  OAI22D1BWP30P140 U91 ( .A1(n55), .A2(n67), .B1(n51), .B2(n39), .ZN(N302) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[16]), .ZN(n68) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[48]), .ZN(n40) );
  OAI22D1BWP30P140 U94 ( .A1(n55), .A2(n68), .B1(n51), .B2(n40), .ZN(N303) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[17]), .ZN(n69) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[49]), .ZN(n41) );
  OAI22D1BWP30P140 U97 ( .A1(n55), .A2(n69), .B1(n51), .B2(n41), .ZN(N304) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[18]), .ZN(n70) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[50]), .ZN(n42) );
  OAI22D1BWP30P140 U100 ( .A1(n55), .A2(n70), .B1(n51), .B2(n42), .ZN(N305) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[22]), .ZN(n75) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[54]), .ZN(n43) );
  OAI22D1BWP30P140 U103 ( .A1(n55), .A2(n75), .B1(n53), .B2(n43), .ZN(N309) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[24]), .ZN(n77) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[56]), .ZN(n44) );
  OAI22D1BWP30P140 U106 ( .A1(n55), .A2(n77), .B1(n53), .B2(n44), .ZN(N311) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[26]), .ZN(n78) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[58]), .ZN(n45) );
  OAI22D1BWP30P140 U109 ( .A1(n55), .A2(n78), .B1(n53), .B2(n45), .ZN(N313) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[28]), .ZN(n79) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[60]), .ZN(n46) );
  OAI22D1BWP30P140 U112 ( .A1(n55), .A2(n79), .B1(n53), .B2(n46), .ZN(N315) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[30]), .ZN(n80) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[62]), .ZN(n47) );
  OAI22D1BWP30P140 U115 ( .A1(n55), .A2(n80), .B1(n53), .B2(n47), .ZN(N317) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[4]), .ZN(n58) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[36]), .ZN(n48) );
  OAI22D1BWP30P140 U118 ( .A1(n55), .A2(n58), .B1(n51), .B2(n48), .ZN(N291) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[37]), .ZN(n49) );
  OAI22D1BWP30P140 U121 ( .A1(n55), .A2(n62), .B1(n53), .B2(n49), .ZN(N292) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[6]), .ZN(n59) );
  INVD1BWP30P140 U123 ( .I(i_data_bus[38]), .ZN(n50) );
  OAI22D1BWP30P140 U124 ( .A1(n55), .A2(n59), .B1(n51), .B2(n50), .ZN(N293) );
  INVD1BWP30P140 U125 ( .I(i_data_bus[39]), .ZN(n52) );
  OAI22D1BWP30P140 U126 ( .A1(n55), .A2(n54), .B1(n53), .B2(n52), .ZN(N294) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n83), .B1(i_data_bus[32]), .B2(n88), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n83), .B1(i_data_bus[34]), .B2(n88), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n83), .B1(i_data_bus[36]), .B2(n88), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n83), .B1(i_data_bus[38]), .B2(n88), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n83), .B1(i_data_bus[33]), .B2(n88), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n83), .B1(i_data_bus[35]), .B2(n88), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n83), .B1(i_data_bus[37]), .B2(n88), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n83), .B1(i_data_bus[40]), .B2(n88), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n83), .B1(i_data_bus[42]), .B2(n88), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n83), .B1(i_data_bus[44]), .B2(n88), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n83), .B1(i_data_bus[46]), .B2(n88), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n83), .B1(i_data_bus[47]), .B2(n88), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n83), .B1(i_data_bus[48]), .B2(n88), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n83), .B1(i_data_bus[49]), .B2(n88), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n83), .B1(i_data_bus[50]), .B2(n88), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n83), .B1(i_data_bus[51]), .B2(n88), 
        .ZN(N338) );
  INVD2BWP30P140 U143 ( .I(n72), .ZN(n89) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n89), .B1(i_data_bus[52]), .B2(n88), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n89), .B1(i_data_bus[53]), .B2(n88), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n89), .B1(i_data_bus[54]), .B2(n88), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n89), .B1(i_data_bus[55]), .B2(n88), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n89), .B1(i_data_bus[56]), .B2(n88), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n89), .B1(i_data_bus[58]), .B2(n88), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n89), .B1(i_data_bus[60]), .B2(n88), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n89), .B1(i_data_bus[62]), .B2(n88), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n83), .B1(i_data_bus[41]), .B2(n88), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n83), .B1(i_data_bus[43]), .B2(n88), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n83), .B1(i_data_bus[45]), .B2(n88), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n89), .B1(i_data_bus[57]), .B2(n88), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n89), .B1(i_data_bus[59]), .B2(n88), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n89), .B1(i_data_bus[61]), .B2(n88), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U158 ( .A1(n90), .A2(n89), .B1(i_data_bus[63]), .B2(n88), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_16 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90;

  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD2BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  ND2OPTIBD1BWP30P140 U3 ( .A1(n9), .A2(n12), .ZN(n7) );
  INVD3BWP30P140 U4 ( .I(n72), .ZN(n83) );
  MOAI22D1BWP30P140 U5 ( .A1(n54), .A2(n83), .B1(i_data_bus[39]), .B2(n88), 
        .ZN(N326) );
  INVD1BWP30P140 U6 ( .I(n88), .ZN(n10) );
  INVD1BWP30P140 U7 ( .I(i_data_bus[7]), .ZN(n54) );
  INVD1BWP30P140 U8 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U9 ( .A1(n1), .A2(i_en), .ZN(n13) );
  NR2D1BWP30P140 U10 ( .A1(n13), .A2(i_cmd[1]), .ZN(n4) );
  INVD2BWP30P140 U11 ( .I(i_valid[0]), .ZN(n2) );
  INVD1BWP30P140 U12 ( .I(i_valid[1]), .ZN(n8) );
  MUX2NUD1BWP30P140 U13 ( .I0(n2), .I1(n8), .S(i_cmd[0]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U14 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U15 ( .I(n5), .ZN(n72) );
  INVD1BWP30P140 U16 ( .I(n13), .ZN(n6) );
  AN3D4BWP30P140 U17 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n6), .Z(n88) );
  INVD2BWP30P140 U18 ( .I(i_cmd[0]), .ZN(n12) );
  INR2D2BWP30P140 U19 ( .A1(i_valid[0]), .B1(n13), .ZN(n9) );
  INVD2BWP30P140 U20 ( .I(n7), .ZN(n31) );
  INVD2BWP30P140 U21 ( .I(n31), .ZN(n30) );
  OAI31D1BWP30P140 U22 ( .A1(n13), .A2(n8), .A3(n12), .B(n30), .ZN(N353) );
  INVD1BWP30P140 U23 ( .I(n9), .ZN(n11) );
  OAI21D1BWP30P140 U24 ( .A1(n11), .A2(i_cmd[1]), .B(n10), .ZN(N354) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[3]), .ZN(n61) );
  MUX2NUD1BWP30P140 U26 ( .I0(n2), .I1(n8), .S(i_cmd[1]), .ZN(n15) );
  NR2D1BWP30P140 U27 ( .A1(n13), .A2(n12), .ZN(n14) );
  CKND2D2BWP30P140 U28 ( .A1(n15), .A2(n14), .ZN(n16) );
  INVD2BWP30P140 U29 ( .I(n16), .ZN(n18) );
  INVD2BWP30P140 U30 ( .I(n18), .ZN(n53) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[35]), .ZN(n17) );
  OAI22D1BWP30P140 U32 ( .A1(n30), .A2(n61), .B1(n53), .B2(n17), .ZN(N290) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[2]), .ZN(n57) );
  INVD2BWP30P140 U34 ( .I(n18), .ZN(n51) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[34]), .ZN(n19) );
  OAI22D1BWP30P140 U36 ( .A1(n30), .A2(n57), .B1(n51), .B2(n19), .ZN(N289) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[1]), .ZN(n60) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[33]), .ZN(n20) );
  OAI22D1BWP30P140 U39 ( .A1(n30), .A2(n60), .B1(n53), .B2(n20), .ZN(N288) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[0]), .ZN(n56) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[32]), .ZN(n21) );
  OAI22D1BWP30P140 U42 ( .A1(n30), .A2(n56), .B1(n51), .B2(n21), .ZN(N287) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[31]), .ZN(n90) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[63]), .ZN(n22) );
  OAI22D1BWP30P140 U45 ( .A1(n30), .A2(n90), .B1(n53), .B2(n22), .ZN(N318) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[29]), .ZN(n87) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[61]), .ZN(n23) );
  OAI22D1BWP30P140 U48 ( .A1(n30), .A2(n87), .B1(n53), .B2(n23), .ZN(N316) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[59]), .ZN(n24) );
  OAI22D1BWP30P140 U51 ( .A1(n30), .A2(n86), .B1(n53), .B2(n24), .ZN(N314) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[25]), .ZN(n85) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[57]), .ZN(n25) );
  OAI22D1BWP30P140 U54 ( .A1(n30), .A2(n85), .B1(n53), .B2(n25), .ZN(N312) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[23]), .ZN(n76) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[55]), .ZN(n26) );
  OAI22D1BWP30P140 U57 ( .A1(n30), .A2(n76), .B1(n53), .B2(n26), .ZN(N310) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[21]), .ZN(n74) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[53]), .ZN(n27) );
  OAI22D1BWP30P140 U60 ( .A1(n30), .A2(n74), .B1(n53), .B2(n27), .ZN(N308) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[20]), .ZN(n73) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[52]), .ZN(n28) );
  OAI22D1BWP30P140 U63 ( .A1(n30), .A2(n73), .B1(n53), .B2(n28), .ZN(N307) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[19]), .ZN(n71) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[51]), .ZN(n29) );
  OAI22D1BWP30P140 U66 ( .A1(n30), .A2(n71), .B1(n51), .B2(n29), .ZN(N306) );
  INVD2BWP30P140 U67 ( .I(n31), .ZN(n55) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[8]), .ZN(n63) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[40]), .ZN(n32) );
  OAI22D1BWP30P140 U70 ( .A1(n55), .A2(n63), .B1(n51), .B2(n32), .ZN(N295) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[9]), .ZN(n81) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[41]), .ZN(n33) );
  OAI22D1BWP30P140 U73 ( .A1(n55), .A2(n81), .B1(n51), .B2(n33), .ZN(N296) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[10]), .ZN(n64) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[42]), .ZN(n34) );
  OAI22D1BWP30P140 U76 ( .A1(n55), .A2(n64), .B1(n51), .B2(n34), .ZN(N297) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[11]), .ZN(n82) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[43]), .ZN(n35) );
  OAI22D1BWP30P140 U79 ( .A1(n55), .A2(n82), .B1(n51), .B2(n35), .ZN(N298) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[12]), .ZN(n65) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[44]), .ZN(n36) );
  OAI22D1BWP30P140 U82 ( .A1(n55), .A2(n65), .B1(n51), .B2(n36), .ZN(N299) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[13]), .ZN(n84) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[45]), .ZN(n37) );
  OAI22D1BWP30P140 U85 ( .A1(n55), .A2(n84), .B1(n51), .B2(n37), .ZN(N300) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[14]), .ZN(n66) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[46]), .ZN(n38) );
  OAI22D1BWP30P140 U88 ( .A1(n55), .A2(n66), .B1(n51), .B2(n38), .ZN(N301) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[15]), .ZN(n67) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[47]), .ZN(n39) );
  OAI22D1BWP30P140 U91 ( .A1(n55), .A2(n67), .B1(n51), .B2(n39), .ZN(N302) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[16]), .ZN(n68) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[48]), .ZN(n40) );
  OAI22D1BWP30P140 U94 ( .A1(n55), .A2(n68), .B1(n51), .B2(n40), .ZN(N303) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[17]), .ZN(n69) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[49]), .ZN(n41) );
  OAI22D1BWP30P140 U97 ( .A1(n55), .A2(n69), .B1(n51), .B2(n41), .ZN(N304) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[18]), .ZN(n70) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[50]), .ZN(n42) );
  OAI22D1BWP30P140 U100 ( .A1(n55), .A2(n70), .B1(n51), .B2(n42), .ZN(N305) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[22]), .ZN(n75) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[54]), .ZN(n43) );
  OAI22D1BWP30P140 U103 ( .A1(n55), .A2(n75), .B1(n53), .B2(n43), .ZN(N309) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[24]), .ZN(n77) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[56]), .ZN(n44) );
  OAI22D1BWP30P140 U106 ( .A1(n55), .A2(n77), .B1(n53), .B2(n44), .ZN(N311) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[26]), .ZN(n78) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[58]), .ZN(n45) );
  OAI22D1BWP30P140 U109 ( .A1(n55), .A2(n78), .B1(n53), .B2(n45), .ZN(N313) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[28]), .ZN(n79) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[60]), .ZN(n46) );
  OAI22D1BWP30P140 U112 ( .A1(n55), .A2(n79), .B1(n53), .B2(n46), .ZN(N315) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[30]), .ZN(n80) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[62]), .ZN(n47) );
  OAI22D1BWP30P140 U115 ( .A1(n55), .A2(n80), .B1(n53), .B2(n47), .ZN(N317) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[4]), .ZN(n58) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[36]), .ZN(n48) );
  OAI22D1BWP30P140 U118 ( .A1(n55), .A2(n58), .B1(n51), .B2(n48), .ZN(N291) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[37]), .ZN(n49) );
  OAI22D1BWP30P140 U121 ( .A1(n55), .A2(n62), .B1(n53), .B2(n49), .ZN(N292) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[6]), .ZN(n59) );
  INVD1BWP30P140 U123 ( .I(i_data_bus[38]), .ZN(n50) );
  OAI22D1BWP30P140 U124 ( .A1(n55), .A2(n59), .B1(n51), .B2(n50), .ZN(N293) );
  INVD1BWP30P140 U125 ( .I(i_data_bus[39]), .ZN(n52) );
  OAI22D1BWP30P140 U126 ( .A1(n55), .A2(n54), .B1(n53), .B2(n52), .ZN(N294) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n83), .B1(i_data_bus[32]), .B2(n88), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n83), .B1(i_data_bus[34]), .B2(n88), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n83), .B1(i_data_bus[36]), .B2(n88), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n83), .B1(i_data_bus[38]), .B2(n88), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n83), .B1(i_data_bus[33]), .B2(n88), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n83), .B1(i_data_bus[35]), .B2(n88), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n83), .B1(i_data_bus[37]), .B2(n88), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n83), .B1(i_data_bus[40]), .B2(n88), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n83), .B1(i_data_bus[42]), .B2(n88), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n83), .B1(i_data_bus[44]), .B2(n88), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n83), .B1(i_data_bus[46]), .B2(n88), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n83), .B1(i_data_bus[47]), .B2(n88), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n83), .B1(i_data_bus[48]), .B2(n88), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n83), .B1(i_data_bus[49]), .B2(n88), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n83), .B1(i_data_bus[50]), .B2(n88), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n83), .B1(i_data_bus[51]), .B2(n88), 
        .ZN(N338) );
  INVD2BWP30P140 U143 ( .I(n72), .ZN(n89) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n89), .B1(i_data_bus[52]), .B2(n88), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n89), .B1(i_data_bus[53]), .B2(n88), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n89), .B1(i_data_bus[54]), .B2(n88), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n89), .B1(i_data_bus[55]), .B2(n88), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n89), .B1(i_data_bus[56]), .B2(n88), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n89), .B1(i_data_bus[58]), .B2(n88), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n89), .B1(i_data_bus[60]), .B2(n88), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n89), .B1(i_data_bus[62]), .B2(n88), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n83), .B1(i_data_bus[41]), .B2(n88), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n83), .B1(i_data_bus[43]), .B2(n88), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n83), .B1(i_data_bus[45]), .B2(n88), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n89), .B1(i_data_bus[57]), .B2(n88), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n89), .B1(i_data_bus[59]), .B2(n88), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n89), .B1(i_data_bus[61]), .B2(n88), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U158 ( .A1(n90), .A2(n89), .B1(i_data_bus[63]), .B2(n88), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_17 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n32), .A2(n6), .B1(n40), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n32), .A2(n7), .B1(n40), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n32), .A2(n8), .B1(n40), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n32), .A2(n9), .B1(n40), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n32), .A2(n10), .B1(n40), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n32), .A2(n11), .B1(n40), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n32), .A2(n12), .B1(n40), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n32), .A2(n13), .B1(n40), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n32), .A2(n14), .B1(n40), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n32), .A2(n16), .B1(n40), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n32), .A2(n15), .B1(n40), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n29), .A2(n28), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n29), .A2(n27), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n29), .A2(n26), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n29), .A2(n25), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n29), .A2(n24), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n29), .A2(n23), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n29), .A2(n22), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n29), .A2(n21), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n29), .A2(n20), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n29), .A2(n19), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n29), .A2(n18), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n29), .A2(n17), .B1(n30), .B2(n92), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[50]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[49]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD2BWP30P140 U68 ( .I(n35), .ZN(n29) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[63]), .ZN(n17) );
  INVD2BWP30P140 U70 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[62]), .ZN(n18) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[61]), .ZN(n19) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[60]), .ZN(n20) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[59]), .ZN(n21) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[58]), .ZN(n22) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[57]), .ZN(n23) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[56]), .ZN(n24) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[55]), .ZN(n25) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[54]), .ZN(n26) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[53]), .ZN(n27) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[52]), .ZN(n28) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[51]), .ZN(n31) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[19]), .ZN(n77) );
  OAI22D1BWP30P140 U96 ( .A1(n32), .A2(n31), .B1(n30), .B2(n77), .ZN(N306) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n64), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n63), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n62), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n61), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n60), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n59), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n58), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n57), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_18 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n6), .B1(n40), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n7), .B1(n40), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n8), .B1(n40), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n9), .B1(n40), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n10), .B1(n40), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n11), .B1(n40), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n12), .B1(n40), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n13), .B1(n40), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n14), .B1(n40), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n15), .B1(n40), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n16), .B1(n40), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n19), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n20), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n21), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n22), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n23), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n24), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n25), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n26), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n27), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n28), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n29), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n31), .B1(n30), .B2(n92), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n77) );
  OAI22D1BWP30P140 U71 ( .A1(n18), .A2(n17), .B1(n30), .B2(n77), .ZN(N306) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n57), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n58), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n59), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n60), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n61), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n62), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n63), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_19 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n25), .A2(n6), .B1(n46), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n25), .A2(n7), .B1(n46), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n25), .A2(n8), .B1(n46), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n25), .A2(n9), .B1(n46), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n25), .A2(n10), .B1(n46), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n25), .A2(n11), .B1(n46), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n25), .A2(n12), .B1(n46), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n25), .A2(n13), .B1(n46), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n25), .A2(n14), .B1(n46), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n25), .A2(n15), .B1(n46), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n25), .A2(n16), .B1(n46), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n26), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n27), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n28), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n29), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n31), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n17), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n18), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n19), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n20), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n21), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n22), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n23), .B1(n30), .B2(n92), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n25) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n46) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD2BWP30P140 U68 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[57]), .ZN(n17) );
  INVD2BWP30P140 U70 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[58]), .ZN(n18) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[59]), .ZN(n19) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[60]), .ZN(n20) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[61]), .ZN(n21) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[62]), .ZN(n22) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[63]), .ZN(n23) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[51]), .ZN(n24) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[19]), .ZN(n77) );
  OAI22D1BWP30P140 U86 ( .A1(n25), .A2(n24), .B1(n30), .B2(n77), .ZN(N306) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[52]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[53]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[54]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[55]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[56]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n40) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n40), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[35]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n60), .B1(n45), .B2(n36), .ZN(N290) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[32]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n57), .B1(n45), .B2(n37), .ZN(N287) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[33]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n58), .B1(n45), .B2(n38), .ZN(N288) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[34]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n59), .B1(n45), .B2(n39), .ZN(N289) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[39]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n64), .B1(n45), .B2(n41), .ZN(N294) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[38]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n63), .B1(n45), .B2(n42), .ZN(N293) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[37]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n62), .B1(n45), .B2(n43), .ZN(N292) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[36]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n61), .B1(n45), .B2(n44), .ZN(N291) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_20 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n74), .ZN(n91) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n74) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n6), .B1(n46), .B2(n92), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n7), .B1(n46), .B2(n89), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n8), .B1(n46), .B2(n88), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n9), .B1(n46), .B2(n65), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n10), .B1(n46), .B2(n66), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n11), .B1(n46), .B2(n67), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n12), .B1(n46), .B2(n68), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n13), .B1(n46), .B2(n69), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n14), .B1(n46), .B2(n70), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n15), .B1(n46), .B2(n71), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n16), .B1(n46), .B2(n72), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n19), .B1(n30), .B2(n75), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n20), .B1(n30), .B2(n76), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n21), .B1(n30), .B2(n77), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n22), .B1(n30), .B2(n78), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n23), .B1(n30), .B2(n79), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n24), .B1(n30), .B2(n80), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n25), .B1(n30), .B2(n81), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n26), .B1(n30), .B2(n82), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n27), .B1(n30), .B2(n83), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n28), .B1(n30), .B2(n84), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n29), .B1(n30), .B2(n85), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n31), .B1(n30), .B2(n87), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n46) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[8]), .ZN(n92) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[9]), .ZN(n89) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[11]), .ZN(n65) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n66) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n67) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[14]), .ZN(n68) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n69) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[16]), .ZN(n70) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[17]), .ZN(n71) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[18]), .ZN(n72) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n73) );
  OAI22D1BWP30P140 U71 ( .A1(n18), .A2(n17), .B1(n30), .B2(n73), .ZN(N306) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n75) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n76) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n77) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n78) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n79) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n80) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n81) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n82) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n83) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n84) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n85) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n87) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n40) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n40), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[32]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n57), .B1(n45), .B2(n36), .ZN(N287) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[33]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n58), .B1(n45), .B2(n37), .ZN(N288) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[34]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n59), .B1(n45), .B2(n38), .ZN(N289) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[35]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n60), .B1(n45), .B2(n39), .ZN(N290) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[36]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n61), .B1(n45), .B2(n41), .ZN(N291) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[37]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n62), .B1(n45), .B2(n42), .ZN(N292) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[38]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n63), .B1(n45), .B2(n43), .ZN(N293) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[39]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N294) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n91), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n91), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n91), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n91), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n91), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n91), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n91), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U145 ( .I(n74), .ZN(n86) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n86), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n86), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n86), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n86), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n86), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n86), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n86), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n86), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n86), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n86), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U156 ( .A1(n85), .A2(n86), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n86), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_21 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n6), .B1(n46), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n7), .B1(n46), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n8), .B1(n46), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n9), .B1(n46), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n10), .B1(n46), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n11), .B1(n46), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n12), .B1(n46), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n16), .B1(n46), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n13), .B1(n46), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n14), .B1(n46), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n15), .B1(n46), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n19), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n20), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n21), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n22), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n23), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n24), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n25), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n26), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n27), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n28), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n29), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n31), .B1(n30), .B2(n92), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n46) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[48]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[49]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[50]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[47]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n77) );
  OAI22D1BWP30P140 U71 ( .A1(n18), .A2(n17), .B1(n30), .B2(n77), .ZN(N306) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n40) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n40), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[32]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n57), .B1(n45), .B2(n36), .ZN(N287) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[33]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n58), .B1(n45), .B2(n37), .ZN(N288) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[34]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n59), .B1(n45), .B2(n38), .ZN(N289) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[35]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n60), .B1(n45), .B2(n39), .ZN(N290) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[36]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n61), .B1(n45), .B2(n41), .ZN(N291) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[37]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n62), .B1(n45), .B2(n42), .ZN(N292) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[38]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n63), .B1(n45), .B2(n43), .ZN(N293) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[39]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N294) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_22 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n6), .B1(n46), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n7), .B1(n46), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n8), .B1(n46), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n9), .B1(n46), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n10), .B1(n46), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n11), .B1(n46), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n12), .B1(n46), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n13), .B1(n46), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n14), .B1(n46), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n15), .B1(n46), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n16), .B1(n46), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n19), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n20), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n21), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n22), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n23), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n24), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n25), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n26), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n27), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n28), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n29), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n31), .B1(n30), .B2(n92), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n46) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n77) );
  OAI22D1BWP30P140 U71 ( .A1(n18), .A2(n17), .B1(n30), .B2(n77), .ZN(N306) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n40) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n40), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[32]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n57), .B1(n45), .B2(n36), .ZN(N287) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[33]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n58), .B1(n45), .B2(n37), .ZN(N288) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[34]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n59), .B1(n45), .B2(n38), .ZN(N289) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[35]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n60), .B1(n45), .B2(n39), .ZN(N290) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[36]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n61), .B1(n45), .B2(n41), .ZN(N291) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[37]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n62), .B1(n45), .B2(n42), .ZN(N292) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[38]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n63), .B1(n45), .B2(n43), .ZN(N293) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[39]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N294) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_23 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n76), .ZN(n91) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n76) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n6), .B1(n43), .B2(n89), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n7), .B1(n43), .B2(n87), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n8), .B1(n43), .B2(n86), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n9), .B1(n43), .B2(n85), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n10), .B1(n43), .B2(n84), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n11), .B1(n43), .B2(n83), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n12), .B1(n43), .B2(n82), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n13), .B1(n43), .B2(n81), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n14), .B1(n43), .B2(n80), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n15), .B1(n43), .B2(n79), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n16), .B1(n43), .B2(n78), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n19), .B1(n30), .B2(n75), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n20), .B1(n30), .B2(n74), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n21), .B1(n30), .B2(n73), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n22), .B1(n30), .B2(n72), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n23), .B1(n30), .B2(n71), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n24), .B1(n30), .B2(n70), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n25), .B1(n30), .B2(n69), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n26), .B1(n30), .B2(n68), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n27), .B1(n30), .B2(n67), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n28), .B1(n30), .B2(n66), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n29), .B1(n30), .B2(n65), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n31), .B1(n30), .B2(n92), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n43) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[8]), .ZN(n89) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[9]), .ZN(n87) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[10]), .ZN(n86) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[11]), .ZN(n85) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n84) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n83) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[14]), .ZN(n82) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n81) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[16]), .ZN(n80) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[17]), .ZN(n79) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[18]), .ZN(n78) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n77) );
  OAI22D1BWP30P140 U71 ( .A1(n18), .A2(n17), .B1(n30), .B2(n77), .ZN(N306) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n75) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n74) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n73) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n72) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n71) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n70) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n69) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n68) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n67) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n66) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n65) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[2]), .ZN(n58) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[34]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n46), .A2(n58), .B1(n45), .B2(n36), .ZN(N289) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[3]), .ZN(n59) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[35]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n46), .A2(n59), .B1(n45), .B2(n37), .ZN(N290) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[36]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n43), .A2(n60), .B1(n45), .B2(n38), .ZN(N291) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[32]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n46), .A2(n57), .B1(n45), .B2(n39), .ZN(N287) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[5]), .ZN(n61) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[37]), .ZN(n40) );
  OAI22D1BWP30P140 U114 ( .A1(n43), .A2(n61), .B1(n45), .B2(n40), .ZN(N292) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[6]), .ZN(n62) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[38]), .ZN(n41) );
  OAI22D1BWP30P140 U117 ( .A1(n43), .A2(n62), .B1(n45), .B2(n41), .ZN(N293) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[7]), .ZN(n63) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[39]), .ZN(n42) );
  OAI22D1BWP30P140 U120 ( .A1(n43), .A2(n63), .B1(n45), .B2(n42), .ZN(N294) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[1]), .ZN(n64) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[33]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N288) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n91), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n91), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n91), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n91), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n91), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n91), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n91), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  INVD2BWP30P140 U147 ( .I(n76), .ZN(n88) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n88), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n88), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n88), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n88), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n88), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n88), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n88), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n88), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U156 ( .A1(n85), .A2(n88), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U157 ( .A1(n86), .A2(n88), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U158 ( .A1(n87), .A2(n88), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n88), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_24 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n6), .B1(n40), .B2(n89), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n7), .B1(n40), .B2(n92), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n8), .B1(n40), .B2(n88), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n9), .B1(n40), .B2(n87), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n10), .B1(n40), .B2(n86), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n11), .B1(n40), .B2(n85), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n12), .B1(n40), .B2(n84), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n13), .B1(n40), .B2(n83), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n14), .B1(n40), .B2(n82), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n15), .B1(n40), .B2(n81), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n16), .B1(n40), .B2(n80), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n19), .B1(n30), .B2(n77), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n20), .B1(n30), .B2(n75), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n21), .B1(n30), .B2(n74), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n22), .B1(n30), .B2(n73), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n23), .B1(n30), .B2(n72), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n24), .B1(n30), .B2(n71), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n25), .B1(n30), .B2(n70), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n26), .B1(n30), .B2(n69), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n27), .B1(n30), .B2(n68), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n28), .B1(n30), .B2(n67), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n29), .B1(n30), .B2(n66), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n31), .B1(n30), .B2(n65), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[8]), .ZN(n89) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[9]), .ZN(n92) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[11]), .ZN(n87) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n85) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[14]), .ZN(n84) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n83) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[16]), .ZN(n82) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[17]), .ZN(n81) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[18]), .ZN(n80) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n79) );
  OAI22D1BWP30P140 U71 ( .A1(n18), .A2(n17), .B1(n30), .B2(n79), .ZN(N306) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n75) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n73) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n72) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n71) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n70) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n68) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n67) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n66) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n65) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n57), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n58), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n59), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n60), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n61), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n62), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n63), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_25 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n8), .B1(n40), .B2(n92), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n9), .B1(n40), .B2(n89), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n10), .B1(n40), .B2(n88), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n11), .B1(n40), .B2(n87), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n12), .B1(n40), .B2(n86), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n13), .B1(n40), .B2(n85), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n14), .B1(n40), .B2(n84), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n15), .B1(n40), .B2(n83), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n16), .B1(n40), .B2(n82), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n6), .B1(n40), .B2(n81), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n7), .B1(n40), .B2(n80), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n19), .B1(n30), .B2(n77), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n20), .B1(n30), .B2(n75), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n21), .B1(n30), .B2(n74), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n22), .B1(n30), .B2(n73), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n23), .B1(n30), .B2(n72), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n24), .B1(n30), .B2(n71), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n25), .B1(n30), .B2(n70), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n26), .B1(n30), .B2(n69), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n27), .B1(n30), .B2(n68), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n28), .B1(n30), .B2(n67), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n29), .B1(n30), .B2(n66), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n31), .B1(n30), .B2(n65), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[49]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[17]), .ZN(n81) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[50]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[18]), .ZN(n80) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[40]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[8]), .ZN(n92) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[41]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[9]), .ZN(n89) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[42]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[43]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[11]), .ZN(n87) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[44]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[45]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[13]), .ZN(n85) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[46]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[14]), .ZN(n84) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[47]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[15]), .ZN(n83) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[48]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[16]), .ZN(n82) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n79) );
  OAI22D1BWP30P140 U71 ( .A1(n18), .A2(n17), .B1(n30), .B2(n79), .ZN(N306) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n75) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n73) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n72) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n71) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n70) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n68) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n67) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n66) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n65) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n57), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n58), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n59), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n60), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n61), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n62), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n63), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_26 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n6), .B1(n40), .B2(n92), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n7), .B1(n40), .B2(n89), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n8), .B1(n40), .B2(n88), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n9), .B1(n40), .B2(n87), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n10), .B1(n40), .B2(n86), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n11), .B1(n40), .B2(n85), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n12), .B1(n40), .B2(n84), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n13), .B1(n40), .B2(n83), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n14), .B1(n40), .B2(n82), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n15), .B1(n40), .B2(n81), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n16), .B1(n40), .B2(n80), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n19), .B1(n30), .B2(n77), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n20), .B1(n30), .B2(n75), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n21), .B1(n30), .B2(n74), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n22), .B1(n30), .B2(n73), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n23), .B1(n30), .B2(n72), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n24), .B1(n30), .B2(n71), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n25), .B1(n30), .B2(n70), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n26), .B1(n30), .B2(n69), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n27), .B1(n30), .B2(n68), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n28), .B1(n30), .B2(n67), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n29), .B1(n30), .B2(n66), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n31), .B1(n30), .B2(n65), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[8]), .ZN(n92) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[9]), .ZN(n89) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[11]), .ZN(n87) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n85) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[14]), .ZN(n84) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n83) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[16]), .ZN(n82) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[17]), .ZN(n81) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[18]), .ZN(n80) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n79) );
  OAI22D1BWP30P140 U71 ( .A1(n18), .A2(n17), .B1(n30), .B2(n79), .ZN(N306) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n75) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n73) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n72) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n71) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n70) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n68) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n67) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n66) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n65) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n57), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n58), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n59), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n60), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n61), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n62), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n63), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_27 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n66), .ZN(n91) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n66) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n6), .B1(n40), .B2(n81), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n7), .B1(n40), .B2(n80), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n8), .B1(n40), .B2(n79), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n9), .B1(n40), .B2(n78), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n10), .B1(n40), .B2(n82), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n11), .B1(n40), .B2(n72), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n12), .B1(n40), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n13), .B1(n40), .B2(n70), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n14), .B1(n40), .B2(n77), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n15), .B1(n40), .B2(n67), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n16), .B1(n40), .B2(n68), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n19), .B1(n30), .B2(n85), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n20), .B1(n30), .B2(n84), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n21), .B1(n30), .B2(n69), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n22), .B1(n30), .B2(n76), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n23), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n24), .B1(n30), .B2(n65), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n25), .B1(n30), .B2(n74), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n26), .B1(n30), .B2(n73), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n27), .B1(n30), .B2(n75), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n28), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n29), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n31), .B1(n30), .B2(n92), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[8]), .ZN(n81) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[9]), .ZN(n80) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[10]), .ZN(n79) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[11]), .ZN(n78) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n82) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n72) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n70) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[16]), .ZN(n77) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[17]), .ZN(n67) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[18]), .ZN(n68) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n87) );
  OAI22D1BWP30P140 U71 ( .A1(n18), .A2(n17), .B1(n30), .B2(n87), .ZN(N306) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n85) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n84) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n69) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n76) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n65) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n74) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n73) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n75) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n57), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n58), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n59), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n60), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n61), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n62), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n63), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n91), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n91), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n91), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n91), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n91), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n91), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n91), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  INVD2BWP30P140 U137 ( .I(n66), .ZN(n86) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n86), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n86), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n86), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n86), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n86), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n86), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n86), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n86), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n86), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n86), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n86), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U156 ( .A1(n85), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n86), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_28 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n12), .B1(n40), .B2(n66), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n15), .B1(n40), .B2(n67), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n13), .B1(n40), .B2(n65), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n14), .B1(n40), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n16), .B1(n40), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n6), .B1(n40), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n7), .B1(n40), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n8), .B1(n40), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n9), .B1(n40), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n10), .B1(n40), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n11), .B1(n40), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n19), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n20), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n21), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n22), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n23), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n24), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n25), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n26), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n27), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n28), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n29), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n31), .B1(n30), .B2(n92), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[45]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[46]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[47]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[48]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[49]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[50]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[40]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[42]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[10]), .ZN(n65) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[43]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[41]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[9]), .ZN(n67) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[44]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n77) );
  OAI22D1BWP30P140 U71 ( .A1(n18), .A2(n17), .B1(n30), .B2(n77), .ZN(N306) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n57), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n58), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n59), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n60), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n61), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n62), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n63), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_29 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n6), .B1(n40), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n7), .B1(n40), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n8), .B1(n40), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n9), .B1(n40), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n10), .B1(n40), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n11), .B1(n40), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n12), .B1(n40), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n13), .B1(n40), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n14), .B1(n40), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n15), .B1(n40), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n16), .B1(n40), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n19), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n20), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n21), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n22), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n23), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n24), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n25), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n26), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n27), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n29), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n28), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n31), .B1(n30), .B2(n92), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n77) );
  OAI22D1BWP30P140 U71 ( .A1(n18), .A2(n17), .B1(n30), .B2(n77), .ZN(N306) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[62]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[61]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n61) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n61), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n57) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n57), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n64) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n64), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n59), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n60), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n62), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n58), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n63) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n63), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_30 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n6), .B1(n46), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n7), .B1(n46), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n8), .B1(n46), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n9), .B1(n46), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n10), .B1(n46), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n11), .B1(n46), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n12), .B1(n46), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n13), .B1(n46), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n14), .B1(n46), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n15), .B1(n46), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n16), .B1(n46), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n19), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n20), .B1(n30), .B2(n92), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n21), .B1(n30), .B2(n80), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n22), .B1(n30), .B2(n81), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n23), .B1(n30), .B2(n82), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n24), .B1(n30), .B2(n83), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n25), .B1(n30), .B2(n84), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n26), .B1(n30), .B2(n85), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n27), .B1(n30), .B2(n86), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n28), .B1(n30), .B2(n87), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n29), .B1(n30), .B2(n88), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n31), .B1(n30), .B2(n89), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n46) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n77) );
  OAI22D1BWP30P140 U71 ( .A1(n18), .A2(n17), .B1(n30), .B2(n77), .ZN(N306) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n92) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n80) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n81) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n82) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n83) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n84) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n85) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n86) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n87) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n88) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n89) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n40) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n40), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[0]), .ZN(n63) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[32]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n63), .B1(n45), .B2(n36), .ZN(N287) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[1]), .ZN(n62) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[33]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n62), .B1(n45), .B2(n37), .ZN(N288) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[2]), .ZN(n61) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[34]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n61), .B1(n45), .B2(n38), .ZN(N289) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[35]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n60), .B1(n45), .B2(n39), .ZN(N290) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[36]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n59), .B1(n45), .B2(n41), .ZN(N291) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[5]), .ZN(n64) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[37]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n64), .B1(n45), .B2(n42), .ZN(N292) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[38]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n58), .B1(n45), .B2(n43), .ZN(N293) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[39]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n57), .B1(n45), .B2(n44), .ZN(N294) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_31 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n6), .B1(n46), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n7), .B1(n46), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n8), .B1(n46), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n9), .B1(n46), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n10), .B1(n46), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n11), .B1(n46), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n12), .B1(n46), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n13), .B1(n46), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n14), .B1(n46), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n15), .B1(n46), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n16), .B1(n46), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n19), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n20), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n21), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n22), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n23), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n24), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n25), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n26), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n27), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n28), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n29), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n31), .B1(n30), .B2(n92), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n46) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n77) );
  OAI22D1BWP30P140 U71 ( .A1(n18), .A2(n17), .B1(n30), .B2(n77), .ZN(N306) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n40) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n40), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[32]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n57), .B1(n45), .B2(n36), .ZN(N287) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[33]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n58), .B1(n45), .B2(n37), .ZN(N288) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[34]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n59), .B1(n45), .B2(n38), .ZN(N289) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[35]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n60), .B1(n45), .B2(n39), .ZN(N290) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[36]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n61), .B1(n45), .B2(n41), .ZN(N291) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[37]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n62), .B1(n45), .B2(n42), .ZN(N292) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[38]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n63), .B1(n45), .B2(n43), .ZN(N293) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[39]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N294) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_32 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n76), .ZN(n91) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n76) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n6), .B1(n46), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n7), .B1(n46), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n8), .B1(n46), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n9), .B1(n46), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n10), .B1(n46), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n11), .B1(n46), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n12), .B1(n46), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n13), .B1(n46), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n14), .B1(n46), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n15), .B1(n46), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n16), .B1(n46), .B2(n92), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n19), .B1(n30), .B2(n77), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n20), .B1(n30), .B2(n78), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n21), .B1(n30), .B2(n79), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n22), .B1(n30), .B2(n80), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n23), .B1(n30), .B2(n81), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n24), .B1(n30), .B2(n82), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n25), .B1(n30), .B2(n83), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n26), .B1(n30), .B2(n84), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n27), .B1(n30), .B2(n85), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n28), .B1(n30), .B2(n86), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n29), .B1(n30), .B2(n87), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n31), .B1(n30), .B2(n89), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n46) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[18]), .ZN(n92) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n75) );
  OAI22D1BWP30P140 U71 ( .A1(n18), .A2(n17), .B1(n30), .B2(n75), .ZN(N306) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n78) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n79) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n80) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n81) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n82) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n83) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n84) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n85) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n86) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n87) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n89) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n40) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n40), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[32]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n57), .B1(n45), .B2(n36), .ZN(N287) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[33]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n58), .B1(n45), .B2(n37), .ZN(N288) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[34]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n59), .B1(n45), .B2(n38), .ZN(N289) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[35]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n60), .B1(n45), .B2(n39), .ZN(N290) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[36]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n61), .B1(n45), .B2(n41), .ZN(N291) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[37]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n62), .B1(n45), .B2(n42), .ZN(N292) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[38]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n63), .B1(n45), .B2(n43), .ZN(N293) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[39]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N294) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n91), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n91), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n91), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n91), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n91), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n91), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n91), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U147 ( .I(n76), .ZN(n88) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n88), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n88), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n88), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n88), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n88), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n88), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n88), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n88), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U156 ( .A1(n85), .A2(n88), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U157 ( .A1(n86), .A2(n88), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U158 ( .A1(n87), .A2(n88), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n88), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_33 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  OAI22D1BWP30P140 U5 ( .A1(n18), .A2(n8), .B1(n46), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U6 ( .A1(n18), .A2(n9), .B1(n46), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U7 ( .A1(n18), .A2(n10), .B1(n46), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U8 ( .A1(n18), .A2(n11), .B1(n46), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U9 ( .A1(n18), .A2(n12), .B1(n46), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n13), .B1(n46), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n14), .B1(n46), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n15), .B1(n46), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n16), .B1(n46), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n6), .B1(n46), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n7), .B1(n46), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U16 ( .A1(n32), .A2(n19), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U17 ( .A1(n32), .A2(n20), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U18 ( .A1(n32), .A2(n21), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U19 ( .A1(n32), .A2(n22), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U20 ( .A1(n32), .A2(n23), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n24), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n25), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n26), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n27), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n28), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n29), .B1(n30), .B2(n92), .ZN(N317) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n31), .B1(n30), .B2(n89), .ZN(N318) );
  ND2OPTIBD1BWP30P140 U28 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U29 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U30 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U31 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U32 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U33 ( .A1(n18), .A2(n17), .B1(n30), .B2(n77), .ZN(N306) );
  INVD1BWP30P140 U34 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U35 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U36 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U38 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U39 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U41 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U42 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[49]), .ZN(n6) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U45 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U46 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U47 ( .I(n33), .ZN(n46) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[50]), .ZN(n7) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[40]), .ZN(n8) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[41]), .ZN(n9) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[42]), .ZN(n10) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[43]), .ZN(n11) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[44]), .ZN(n12) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[45]), .ZN(n13) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[46]), .ZN(n14) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[47]), .ZN(n15) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[48]), .ZN(n16) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U70 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n77) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n92) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n89) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n40) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n40), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[32]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n64), .B1(n45), .B2(n36), .ZN(N287) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[33]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n63), .B1(n45), .B2(n37), .ZN(N288) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[34]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n62), .B1(n45), .B2(n38), .ZN(N289) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[35]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n61), .B1(n45), .B2(n39), .ZN(N290) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[36]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n60), .B1(n45), .B2(n41), .ZN(N291) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[37]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n59), .B1(n45), .B2(n42), .ZN(N292) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[38]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n58), .B1(n45), .B2(n43), .ZN(N293) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[39]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n57), .B1(n45), .B2(n44), .ZN(N294) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_34 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  OAI22D1BWP30P140 U5 ( .A1(n18), .A2(n6), .B1(n46), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U6 ( .A1(n18), .A2(n7), .B1(n46), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U7 ( .A1(n18), .A2(n8), .B1(n46), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U8 ( .A1(n18), .A2(n9), .B1(n46), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U9 ( .A1(n18), .A2(n10), .B1(n46), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n11), .B1(n46), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n12), .B1(n46), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n13), .B1(n46), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n14), .B1(n46), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n15), .B1(n46), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n16), .B1(n46), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U16 ( .A1(n32), .A2(n19), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U17 ( .A1(n32), .A2(n20), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U18 ( .A1(n32), .A2(n21), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U19 ( .A1(n32), .A2(n22), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U20 ( .A1(n32), .A2(n23), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n24), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n25), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n26), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n27), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n28), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n29), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n31), .B1(n30), .B2(n92), .ZN(N318) );
  ND2OPTIBD1BWP30P140 U28 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U29 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U30 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U31 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U32 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U33 ( .A1(n18), .A2(n17), .B1(n30), .B2(n77), .ZN(N306) );
  INVD1BWP30P140 U34 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U35 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U36 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U38 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U39 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U41 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U42 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U45 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U46 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U47 ( .I(n33), .ZN(n46) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U70 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n77) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n40) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n40), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[0]), .ZN(n63) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[32]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n63), .B1(n45), .B2(n36), .ZN(N287) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[1]), .ZN(n62) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[33]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n62), .B1(n45), .B2(n37), .ZN(N288) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[2]), .ZN(n61) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[34]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n61), .B1(n45), .B2(n38), .ZN(N289) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[35]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n60), .B1(n45), .B2(n39), .ZN(N290) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[36]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n59), .B1(n45), .B2(n41), .ZN(N291) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[5]), .ZN(n58) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[37]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n58), .B1(n45), .B2(n42), .ZN(N292) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[6]), .ZN(n57) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[38]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n57), .B1(n45), .B2(n43), .ZN(N293) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[39]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N294) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_35 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  INVD3BWP30P140 U3 ( .I(n73), .ZN(n91) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n73) );
  OAI22D1BWP30P140 U5 ( .A1(n18), .A2(n6), .B1(n46), .B2(n74), .ZN(N295) );
  OAI22D1BWP30P140 U6 ( .A1(n18), .A2(n7), .B1(n46), .B2(n75), .ZN(N296) );
  OAI22D1BWP30P140 U7 ( .A1(n18), .A2(n8), .B1(n46), .B2(n76), .ZN(N297) );
  OAI22D1BWP30P140 U8 ( .A1(n18), .A2(n9), .B1(n46), .B2(n77), .ZN(N298) );
  OAI22D1BWP30P140 U9 ( .A1(n18), .A2(n10), .B1(n46), .B2(n78), .ZN(N299) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n11), .B1(n46), .B2(n79), .ZN(N300) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n12), .B1(n46), .B2(n80), .ZN(N301) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n13), .B1(n46), .B2(n81), .ZN(N302) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n14), .B1(n46), .B2(n82), .ZN(N303) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n15), .B1(n46), .B2(n83), .ZN(N304) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n16), .B1(n46), .B2(n84), .ZN(N305) );
  OAI22D1BWP30P140 U16 ( .A1(n32), .A2(n31), .B1(n30), .B2(n87), .ZN(N307) );
  OAI22D1BWP30P140 U17 ( .A1(n32), .A2(n19), .B1(n30), .B2(n88), .ZN(N308) );
  OAI22D1BWP30P140 U18 ( .A1(n32), .A2(n20), .B1(n30), .B2(n89), .ZN(N309) );
  OAI22D1BWP30P140 U19 ( .A1(n32), .A2(n21), .B1(n30), .B2(n92), .ZN(N310) );
  OAI22D1BWP30P140 U20 ( .A1(n32), .A2(n22), .B1(n30), .B2(n72), .ZN(N311) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n23), .B1(n30), .B2(n71), .ZN(N312) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n24), .B1(n30), .B2(n65), .ZN(N313) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n25), .B1(n30), .B2(n66), .ZN(N314) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n26), .B1(n30), .B2(n67), .ZN(N315) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n27), .B1(n30), .B2(n68), .ZN(N316) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n28), .B1(n30), .B2(n69), .ZN(N317) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n29), .B1(n30), .B2(n70), .ZN(N318) );
  ND2OPTIBD1BWP30P140 U28 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U29 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U30 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U31 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U32 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U33 ( .A1(n18), .A2(n17), .B1(n30), .B2(n86), .ZN(N306) );
  INVD1BWP30P140 U34 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U35 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U36 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U38 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U39 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U41 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U42 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U45 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U46 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U47 ( .I(n33), .ZN(n46) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n74) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n75) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n76) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n77) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n78) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n79) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[14]), .ZN(n80) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[15]), .ZN(n81) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n82) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n83) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n84) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U70 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n86) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[53]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[21]), .ZN(n88) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[54]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[22]), .ZN(n89) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[55]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[23]), .ZN(n92) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[56]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[24]), .ZN(n72) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[57]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[25]), .ZN(n71) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[58]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[26]), .ZN(n65) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[59]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[27]), .ZN(n66) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[60]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[28]), .ZN(n67) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[61]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[29]), .ZN(n68) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[62]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[30]), .ZN(n69) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[63]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[31]), .ZN(n70) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[52]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[20]), .ZN(n87) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n40) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n40), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[32]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n64), .B1(n45), .B2(n36), .ZN(N287) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[33]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n63), .B1(n45), .B2(n37), .ZN(N288) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[34]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n62), .B1(n45), .B2(n38), .ZN(N289) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[35]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n61), .B1(n45), .B2(n39), .ZN(N290) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[36]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n60), .B1(n45), .B2(n41), .ZN(N291) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[37]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n59), .B1(n45), .B2(n42), .ZN(N292) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[38]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n58), .B1(n45), .B2(n43), .ZN(N293) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[39]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n57), .B1(n45), .B2(n44), .ZN(N294) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n91), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n91), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n91), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n91), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n91), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n91), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n91), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  INVD2BWP30P140 U144 ( .I(n73), .ZN(n85) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n85), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n85), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n85), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n85), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n85), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n85), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n85), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n85), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n85), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n85), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n85), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n85), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_36 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  OAI22D1BWP30P140 U5 ( .A1(n18), .A2(n6), .B1(n41), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U6 ( .A1(n18), .A2(n7), .B1(n41), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U7 ( .A1(n18), .A2(n8), .B1(n41), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U8 ( .A1(n18), .A2(n9), .B1(n41), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U9 ( .A1(n18), .A2(n10), .B1(n41), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n11), .B1(n41), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n12), .B1(n41), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n13), .B1(n41), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n14), .B1(n41), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n15), .B1(n41), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n16), .B1(n41), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U16 ( .A1(n32), .A2(n19), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U17 ( .A1(n32), .A2(n20), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U18 ( .A1(n32), .A2(n21), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U19 ( .A1(n32), .A2(n22), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U20 ( .A1(n32), .A2(n23), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n24), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n25), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n26), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n27), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n28), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n29), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n31), .B1(n30), .B2(n92), .ZN(N318) );
  ND2OPTIBD1BWP30P140 U28 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U29 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U30 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U31 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U32 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U33 ( .A1(n18), .A2(n17), .B1(n30), .B2(n77), .ZN(N306) );
  INVD1BWP30P140 U34 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U35 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U36 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U38 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U39 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U41 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U42 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U45 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U46 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U47 ( .I(n33), .ZN(n41) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U70 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n77) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[35]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n46), .A2(n61), .B1(n45), .B2(n36), .ZN(N290) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[37]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n41), .A2(n59), .B1(n45), .B2(n37), .ZN(N292) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[36]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n41), .A2(n60), .B1(n45), .B2(n38), .ZN(N291) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[39]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n41), .A2(n57), .B1(n45), .B2(n39), .ZN(N294) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[38]), .ZN(n40) );
  OAI22D1BWP30P140 U114 ( .A1(n41), .A2(n58), .B1(n45), .B2(n40), .ZN(N293) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n62), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n63), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_37 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n7), .B1(n46), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n6), .B1(n46), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n15), .B1(n46), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n16), .B1(n46), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n8), .B1(n46), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n9), .B1(n46), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n10), .B1(n46), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n11), .B1(n46), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n12), .B1(n46), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n13), .B1(n46), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n14), .B1(n46), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n19), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n20), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n21), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n22), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n23), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n24), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n25), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n26), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n27), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n28), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n29), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n31), .B1(n30), .B2(n92), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[41]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n46) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[40]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[44]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[45]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[46]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[47]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[48]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[49]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[50]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[42]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[43]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n77) );
  OAI22D1BWP30P140 U71 ( .A1(n18), .A2(n17), .B1(n30), .B2(n77), .ZN(N306) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n40) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n40), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[32]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n57), .B1(n45), .B2(n36), .ZN(N287) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[33]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n58), .B1(n45), .B2(n37), .ZN(N288) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[34]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n59), .B1(n45), .B2(n38), .ZN(N289) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[35]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n60), .B1(n45), .B2(n39), .ZN(N290) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[36]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n61), .B1(n45), .B2(n41), .ZN(N291) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[37]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n62), .B1(n45), .B2(n42), .ZN(N292) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[39]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n64), .B1(n45), .B2(n43), .ZN(N294) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[38]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n63), .B1(n45), .B2(n44), .ZN(N293) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_38 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n75), .ZN(n91) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n75) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n32), .A2(n16), .B1(n46), .B2(n88), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n32), .A2(n15), .B1(n46), .B2(n86), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n32), .A2(n14), .B1(n46), .B2(n85), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n32), .A2(n13), .B1(n46), .B2(n84), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n32), .A2(n12), .B1(n46), .B2(n83), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n32), .A2(n11), .B1(n46), .B2(n82), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n32), .A2(n10), .B1(n46), .B2(n81), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n32), .A2(n9), .B1(n46), .B2(n80), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n32), .A2(n8), .B1(n46), .B2(n79), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n32), .A2(n7), .B1(n46), .B2(n78), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n32), .A2(n6), .B1(n46), .B2(n77), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n29), .A2(n28), .B1(n30), .B2(n74), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n29), .A2(n27), .B1(n30), .B2(n73), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n29), .A2(n26), .B1(n30), .B2(n72), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n29), .A2(n25), .B1(n30), .B2(n71), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n29), .A2(n24), .B1(n30), .B2(n70), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n29), .A2(n23), .B1(n30), .B2(n69), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n29), .A2(n22), .B1(n30), .B2(n68), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n29), .A2(n21), .B1(n30), .B2(n67), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n29), .A2(n20), .B1(n30), .B2(n66), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n29), .A2(n19), .B1(n30), .B2(n65), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n29), .A2(n18), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n29), .A2(n17), .B1(n30), .B2(n92), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[50]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n46) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[18]), .ZN(n77) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[49]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[17]), .ZN(n78) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[48]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[16]), .ZN(n79) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[47]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[15]), .ZN(n80) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[46]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[14]), .ZN(n81) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n82) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[44]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[12]), .ZN(n83) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[43]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[11]), .ZN(n84) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[42]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[10]), .ZN(n85) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[41]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[9]), .ZN(n86) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[40]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[8]), .ZN(n88) );
  INVD2BWP30P140 U68 ( .I(n35), .ZN(n29) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[63]), .ZN(n17) );
  INVD2BWP30P140 U70 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[62]), .ZN(n18) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[61]), .ZN(n19) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[29]), .ZN(n65) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[60]), .ZN(n20) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[28]), .ZN(n66) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[59]), .ZN(n21) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[27]), .ZN(n67) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[58]), .ZN(n22) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[26]), .ZN(n68) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[57]), .ZN(n23) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[25]), .ZN(n69) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[56]), .ZN(n24) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[24]), .ZN(n70) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[55]), .ZN(n25) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[23]), .ZN(n71) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[54]), .ZN(n26) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[22]), .ZN(n72) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[53]), .ZN(n27) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[21]), .ZN(n73) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[52]), .ZN(n28) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[20]), .ZN(n74) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[51]), .ZN(n31) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[19]), .ZN(n76) );
  OAI22D1BWP30P140 U96 ( .A1(n32), .A2(n31), .B1(n30), .B2(n76), .ZN(N306) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n40) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n40), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[32]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n64), .B1(n45), .B2(n36), .ZN(N287) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[33]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n63), .B1(n45), .B2(n37), .ZN(N288) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[34]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n62), .B1(n45), .B2(n38), .ZN(N289) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[35]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n61), .B1(n45), .B2(n39), .ZN(N290) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[36]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n60), .B1(n45), .B2(n41), .ZN(N291) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[37]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n59), .B1(n45), .B2(n42), .ZN(N292) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[38]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n58), .B1(n45), .B2(n43), .ZN(N293) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[39]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n57), .B1(n45), .B2(n44), .ZN(N294) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n91), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n91), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n91), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n91), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n91), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n91), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n91), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  INVD2BWP30P140 U146 ( .I(n75), .ZN(n87) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n87), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n87), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n87), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n87), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n87), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n87), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n87), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n87), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n87), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U156 ( .A1(n85), .A2(n87), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U157 ( .A1(n86), .A2(n87), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n87), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_39 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n32), .A2(n16), .B1(n46), .B2(n92), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n32), .A2(n15), .B1(n46), .B2(n89), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n32), .A2(n14), .B1(n46), .B2(n88), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n32), .A2(n13), .B1(n46), .B2(n87), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n32), .A2(n12), .B1(n46), .B2(n86), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n32), .A2(n11), .B1(n46), .B2(n85), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n32), .A2(n10), .B1(n46), .B2(n84), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n32), .A2(n9), .B1(n46), .B2(n83), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n32), .A2(n8), .B1(n46), .B2(n82), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n32), .A2(n7), .B1(n46), .B2(n81), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n32), .A2(n6), .B1(n46), .B2(n80), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n29), .A2(n28), .B1(n30), .B2(n77), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n29), .A2(n27), .B1(n30), .B2(n75), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n29), .A2(n26), .B1(n30), .B2(n74), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n29), .A2(n25), .B1(n30), .B2(n73), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n29), .A2(n24), .B1(n30), .B2(n72), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n29), .A2(n23), .B1(n30), .B2(n71), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n29), .A2(n22), .B1(n30), .B2(n70), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n29), .A2(n21), .B1(n30), .B2(n69), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n29), .A2(n20), .B1(n30), .B2(n68), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n29), .A2(n19), .B1(n30), .B2(n67), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n29), .A2(n18), .B1(n30), .B2(n66), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n29), .A2(n17), .B1(n30), .B2(n65), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[50]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n46) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[18]), .ZN(n80) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[49]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[17]), .ZN(n81) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[48]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[16]), .ZN(n82) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[47]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[15]), .ZN(n83) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[46]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[14]), .ZN(n84) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n85) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[44]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[43]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[11]), .ZN(n87) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[42]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[41]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[9]), .ZN(n89) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[40]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[8]), .ZN(n92) );
  INVD2BWP30P140 U68 ( .I(n35), .ZN(n29) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[63]), .ZN(n17) );
  INVD2BWP30P140 U70 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[31]), .ZN(n65) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[62]), .ZN(n18) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[30]), .ZN(n66) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[61]), .ZN(n19) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[29]), .ZN(n67) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[60]), .ZN(n20) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[28]), .ZN(n68) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[59]), .ZN(n21) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[58]), .ZN(n22) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[26]), .ZN(n70) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[57]), .ZN(n23) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[25]), .ZN(n71) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[56]), .ZN(n24) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[24]), .ZN(n72) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[55]), .ZN(n25) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[23]), .ZN(n73) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[54]), .ZN(n26) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[53]), .ZN(n27) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[21]), .ZN(n75) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[52]), .ZN(n28) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[51]), .ZN(n31) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[19]), .ZN(n79) );
  OAI22D1BWP30P140 U96 ( .A1(n32), .A2(n31), .B1(n30), .B2(n79), .ZN(N306) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n43) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n43), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[37]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n46), .A2(n62), .B1(n45), .B2(n36), .ZN(N292) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[39]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n46), .A2(n64), .B1(n45), .B2(n37), .ZN(N294) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[36]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n46), .A2(n61), .B1(n45), .B2(n38), .ZN(N291) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[35]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n43), .A2(n60), .B1(n45), .B2(n39), .ZN(N290) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[34]), .ZN(n40) );
  OAI22D1BWP30P140 U114 ( .A1(n43), .A2(n59), .B1(n45), .B2(n40), .ZN(N289) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[33]), .ZN(n41) );
  OAI22D1BWP30P140 U117 ( .A1(n43), .A2(n58), .B1(n45), .B2(n41), .ZN(N288) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[32]), .ZN(n42) );
  OAI22D1BWP30P140 U120 ( .A1(n43), .A2(n57), .B1(n45), .B2(n42), .ZN(N287) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[38]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n63), .B1(n45), .B2(n44), .ZN(N293) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_40 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n16), .B1(n40), .B2(n92), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n15), .B1(n40), .B2(n89), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n14), .B1(n40), .B2(n88), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n13), .B1(n40), .B2(n87), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n12), .B1(n40), .B2(n86), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n11), .B1(n40), .B2(n85), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n10), .B1(n40), .B2(n84), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n9), .B1(n40), .B2(n83), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n8), .B1(n40), .B2(n82), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n7), .B1(n40), .B2(n81), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n6), .B1(n40), .B2(n80), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n19), .B1(n30), .B2(n77), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n31), .B1(n30), .B2(n75), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n29), .B1(n30), .B2(n74), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n28), .B1(n30), .B2(n73), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n27), .B1(n30), .B2(n72), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n26), .B1(n30), .B2(n71), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n25), .B1(n30), .B2(n70), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n24), .B1(n30), .B2(n69), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n23), .B1(n30), .B2(n68), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n22), .B1(n30), .B2(n67), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n21), .B1(n30), .B2(n66), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n20), .B1(n30), .B2(n65), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[50]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[18]), .ZN(n80) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[49]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[17]), .ZN(n81) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[48]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[16]), .ZN(n82) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[47]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[15]), .ZN(n83) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[46]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[14]), .ZN(n84) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n85) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[44]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[43]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[11]), .ZN(n87) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[42]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[41]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[9]), .ZN(n89) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[40]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[8]), .ZN(n92) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n79) );
  OAI22D1BWP30P140 U71 ( .A1(n18), .A2(n17), .B1(n30), .B2(n79), .ZN(N306) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[63]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[31]), .ZN(n65) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[62]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[30]), .ZN(n66) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[61]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[29]), .ZN(n67) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[60]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[28]), .ZN(n68) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[59]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n70) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[57]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[25]), .ZN(n71) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[56]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[24]), .ZN(n72) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[55]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[23]), .ZN(n73) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[54]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[53]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[21]), .ZN(n75) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n64), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n57) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n57), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n63) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n63), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n62), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n61), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n60), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n59), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n58) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n58), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_41 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  OAI22D1BWP30P140 U5 ( .A1(n32), .A2(n16), .B1(n40), .B2(n92), .ZN(N295) );
  OAI22D1BWP30P140 U6 ( .A1(n32), .A2(n15), .B1(n40), .B2(n89), .ZN(N296) );
  OAI22D1BWP30P140 U7 ( .A1(n32), .A2(n14), .B1(n40), .B2(n88), .ZN(N297) );
  OAI22D1BWP30P140 U8 ( .A1(n32), .A2(n13), .B1(n40), .B2(n87), .ZN(N298) );
  OAI22D1BWP30P140 U9 ( .A1(n32), .A2(n12), .B1(n40), .B2(n86), .ZN(N299) );
  OAI22D1BWP30P140 U10 ( .A1(n32), .A2(n11), .B1(n40), .B2(n85), .ZN(N300) );
  OAI22D1BWP30P140 U11 ( .A1(n32), .A2(n10), .B1(n40), .B2(n84), .ZN(N301) );
  OAI22D1BWP30P140 U12 ( .A1(n32), .A2(n9), .B1(n40), .B2(n83), .ZN(N302) );
  OAI22D1BWP30P140 U13 ( .A1(n32), .A2(n8), .B1(n40), .B2(n82), .ZN(N303) );
  OAI22D1BWP30P140 U14 ( .A1(n32), .A2(n7), .B1(n40), .B2(n81), .ZN(N304) );
  OAI22D1BWP30P140 U15 ( .A1(n32), .A2(n6), .B1(n40), .B2(n80), .ZN(N305) );
  OAI22D1BWP30P140 U16 ( .A1(n29), .A2(n28), .B1(n30), .B2(n77), .ZN(N307) );
  OAI22D1BWP30P140 U17 ( .A1(n29), .A2(n27), .B1(n30), .B2(n75), .ZN(N308) );
  OAI22D1BWP30P140 U18 ( .A1(n29), .A2(n26), .B1(n30), .B2(n74), .ZN(N309) );
  OAI22D1BWP30P140 U19 ( .A1(n29), .A2(n25), .B1(n30), .B2(n73), .ZN(N310) );
  OAI22D1BWP30P140 U20 ( .A1(n29), .A2(n24), .B1(n30), .B2(n72), .ZN(N311) );
  OAI22D1BWP30P140 U21 ( .A1(n29), .A2(n23), .B1(n30), .B2(n71), .ZN(N312) );
  OAI22D1BWP30P140 U22 ( .A1(n29), .A2(n22), .B1(n30), .B2(n70), .ZN(N313) );
  OAI22D1BWP30P140 U23 ( .A1(n29), .A2(n21), .B1(n30), .B2(n69), .ZN(N314) );
  OAI22D1BWP30P140 U24 ( .A1(n29), .A2(n20), .B1(n30), .B2(n68), .ZN(N315) );
  OAI22D1BWP30P140 U25 ( .A1(n29), .A2(n19), .B1(n30), .B2(n67), .ZN(N316) );
  OAI22D1BWP30P140 U26 ( .A1(n29), .A2(n18), .B1(n30), .B2(n66), .ZN(N317) );
  OAI22D1BWP30P140 U27 ( .A1(n29), .A2(n17), .B1(n30), .B2(n65), .ZN(N318) );
  ND2OPTIBD1BWP30P140 U28 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U29 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U30 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U31 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U32 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U33 ( .A1(n32), .A2(n31), .B1(n30), .B2(n79), .ZN(N306) );
  INVD1BWP30P140 U34 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U35 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U36 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U38 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U39 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U41 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U42 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[50]), .ZN(n6) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U45 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U46 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U47 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[18]), .ZN(n80) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[49]), .ZN(n7) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[17]), .ZN(n81) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[48]), .ZN(n8) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[16]), .ZN(n82) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[47]), .ZN(n9) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[15]), .ZN(n83) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[46]), .ZN(n10) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[14]), .ZN(n84) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n85) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[44]), .ZN(n12) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[43]), .ZN(n13) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[11]), .ZN(n87) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[42]), .ZN(n14) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[41]), .ZN(n15) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[9]), .ZN(n89) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[40]), .ZN(n16) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[8]), .ZN(n92) );
  INVD2BWP30P140 U69 ( .I(n35), .ZN(n29) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[63]), .ZN(n17) );
  INVD2BWP30P140 U71 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[31]), .ZN(n65) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[62]), .ZN(n18) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[30]), .ZN(n66) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[61]), .ZN(n19) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[29]), .ZN(n67) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[60]), .ZN(n20) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[28]), .ZN(n68) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[59]), .ZN(n21) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[58]), .ZN(n22) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[26]), .ZN(n70) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n23) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n71) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[56]), .ZN(n24) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[24]), .ZN(n72) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[55]), .ZN(n25) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[23]), .ZN(n73) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[54]), .ZN(n26) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[53]), .ZN(n27) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[21]), .ZN(n75) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[52]), .ZN(n28) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[51]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[19]), .ZN(n79) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n62) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n62), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n61) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n61), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n60) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n60), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n59), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n58) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n58), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n57) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n57), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n63), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_42 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  OAI22D1BWP30P140 U5 ( .A1(n29), .A2(n16), .B1(n40), .B2(n77), .ZN(N295) );
  OAI22D1BWP30P140 U6 ( .A1(n29), .A2(n15), .B1(n40), .B2(n75), .ZN(N296) );
  OAI22D1BWP30P140 U7 ( .A1(n29), .A2(n14), .B1(n40), .B2(n74), .ZN(N297) );
  OAI22D1BWP30P140 U8 ( .A1(n29), .A2(n13), .B1(n40), .B2(n73), .ZN(N298) );
  OAI22D1BWP30P140 U9 ( .A1(n29), .A2(n12), .B1(n40), .B2(n72), .ZN(N299) );
  OAI22D1BWP30P140 U10 ( .A1(n29), .A2(n11), .B1(n40), .B2(n71), .ZN(N300) );
  OAI22D1BWP30P140 U11 ( .A1(n29), .A2(n10), .B1(n40), .B2(n70), .ZN(N301) );
  OAI22D1BWP30P140 U12 ( .A1(n29), .A2(n9), .B1(n40), .B2(n69), .ZN(N302) );
  OAI22D1BWP30P140 U13 ( .A1(n29), .A2(n8), .B1(n40), .B2(n68), .ZN(N303) );
  OAI22D1BWP30P140 U14 ( .A1(n29), .A2(n7), .B1(n40), .B2(n67), .ZN(N304) );
  OAI22D1BWP30P140 U15 ( .A1(n29), .A2(n6), .B1(n40), .B2(n66), .ZN(N305) );
  OAI22D1BWP30P140 U16 ( .A1(n32), .A2(n27), .B1(n30), .B2(n92), .ZN(N307) );
  OAI22D1BWP30P140 U17 ( .A1(n32), .A2(n31), .B1(n30), .B2(n89), .ZN(N308) );
  OAI22D1BWP30P140 U18 ( .A1(n32), .A2(n26), .B1(n30), .B2(n88), .ZN(N309) );
  OAI22D1BWP30P140 U19 ( .A1(n32), .A2(n25), .B1(n30), .B2(n87), .ZN(N310) );
  OAI22D1BWP30P140 U20 ( .A1(n32), .A2(n24), .B1(n30), .B2(n86), .ZN(N311) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n23), .B1(n30), .B2(n85), .ZN(N312) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n22), .B1(n30), .B2(n84), .ZN(N313) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n21), .B1(n30), .B2(n83), .ZN(N314) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n20), .B1(n30), .B2(n82), .ZN(N315) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n19), .B1(n30), .B2(n81), .ZN(N316) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n18), .B1(n30), .B2(n80), .ZN(N317) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n17), .B1(n30), .B2(n79), .ZN(N318) );
  ND2OPTIBD1BWP30P140 U28 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U29 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U30 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U31 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U32 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U33 ( .A1(n29), .A2(n28), .B1(n30), .B2(n65), .ZN(N306) );
  INVD1BWP30P140 U34 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U35 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U36 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U38 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U39 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U41 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U42 ( .I(n35), .ZN(n29) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[50]), .ZN(n6) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U45 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U46 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U47 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[18]), .ZN(n66) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[49]), .ZN(n7) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[17]), .ZN(n67) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[48]), .ZN(n8) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[16]), .ZN(n68) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[47]), .ZN(n9) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[15]), .ZN(n69) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[46]), .ZN(n10) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[14]), .ZN(n70) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n71) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[44]), .ZN(n12) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[12]), .ZN(n72) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[43]), .ZN(n13) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[11]), .ZN(n73) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[42]), .ZN(n14) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[10]), .ZN(n74) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[41]), .ZN(n15) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[9]), .ZN(n75) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[40]), .ZN(n16) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[8]), .ZN(n77) );
  INVD2BWP30P140 U69 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[63]), .ZN(n17) );
  INVD2BWP30P140 U71 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[31]), .ZN(n79) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[62]), .ZN(n18) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[30]), .ZN(n80) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[61]), .ZN(n19) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[29]), .ZN(n81) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[60]), .ZN(n20) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[28]), .ZN(n82) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[59]), .ZN(n21) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[27]), .ZN(n83) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[58]), .ZN(n22) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[26]), .ZN(n84) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n23) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n85) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[56]), .ZN(n24) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[24]), .ZN(n86) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[55]), .ZN(n25) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[23]), .ZN(n87) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[54]), .ZN(n26) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[22]), .ZN(n88) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[52]), .ZN(n27) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[20]), .ZN(n92) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[51]), .ZN(n28) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[19]), .ZN(n65) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[53]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[21]), .ZN(n89) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n64), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n63), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n62), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n61), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n60), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n59), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n58), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n57), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_43 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n71), .ZN(n91) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n71) );
  OAI22D1BWP30P140 U5 ( .A1(n32), .A2(n16), .B1(n40), .B2(n68), .ZN(N295) );
  OAI22D1BWP30P140 U6 ( .A1(n32), .A2(n15), .B1(n40), .B2(n67), .ZN(N296) );
  OAI22D1BWP30P140 U7 ( .A1(n32), .A2(n14), .B1(n40), .B2(n66), .ZN(N297) );
  OAI22D1BWP30P140 U8 ( .A1(n32), .A2(n13), .B1(n40), .B2(n65), .ZN(N298) );
  OAI22D1BWP30P140 U9 ( .A1(n32), .A2(n12), .B1(n40), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U10 ( .A1(n32), .A2(n11), .B1(n40), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U11 ( .A1(n32), .A2(n10), .B1(n40), .B2(n92), .ZN(N301) );
  OAI22D1BWP30P140 U12 ( .A1(n32), .A2(n9), .B1(n40), .B2(n89), .ZN(N302) );
  OAI22D1BWP30P140 U13 ( .A1(n32), .A2(n8), .B1(n40), .B2(n88), .ZN(N303) );
  OAI22D1BWP30P140 U14 ( .A1(n32), .A2(n7), .B1(n40), .B2(n87), .ZN(N304) );
  OAI22D1BWP30P140 U15 ( .A1(n32), .A2(n6), .B1(n40), .B2(n86), .ZN(N305) );
  OAI22D1BWP30P140 U16 ( .A1(n29), .A2(n28), .B1(n30), .B2(n84), .ZN(N307) );
  OAI22D1BWP30P140 U17 ( .A1(n29), .A2(n27), .B1(n30), .B2(n82), .ZN(N308) );
  OAI22D1BWP30P140 U18 ( .A1(n29), .A2(n26), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U19 ( .A1(n29), .A2(n25), .B1(n30), .B2(n80), .ZN(N310) );
  OAI22D1BWP30P140 U20 ( .A1(n29), .A2(n24), .B1(n30), .B2(n79), .ZN(N311) );
  OAI22D1BWP30P140 U21 ( .A1(n29), .A2(n23), .B1(n30), .B2(n78), .ZN(N312) );
  OAI22D1BWP30P140 U22 ( .A1(n29), .A2(n22), .B1(n30), .B2(n77), .ZN(N313) );
  OAI22D1BWP30P140 U23 ( .A1(n29), .A2(n21), .B1(n30), .B2(n76), .ZN(N314) );
  OAI22D1BWP30P140 U24 ( .A1(n29), .A2(n20), .B1(n30), .B2(n75), .ZN(N315) );
  OAI22D1BWP30P140 U25 ( .A1(n29), .A2(n19), .B1(n30), .B2(n74), .ZN(N316) );
  OAI22D1BWP30P140 U26 ( .A1(n29), .A2(n18), .B1(n30), .B2(n73), .ZN(N317) );
  OAI22D1BWP30P140 U27 ( .A1(n29), .A2(n17), .B1(n30), .B2(n72), .ZN(N318) );
  ND2OPTIBD1BWP30P140 U28 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U29 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U30 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U31 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U32 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U33 ( .A1(n32), .A2(n31), .B1(n30), .B2(n85), .ZN(N306) );
  INVD1BWP30P140 U34 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U35 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U36 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U38 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U39 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U41 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U42 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[50]), .ZN(n6) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U45 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U46 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U47 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[18]), .ZN(n86) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[49]), .ZN(n7) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[17]), .ZN(n87) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[48]), .ZN(n8) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[16]), .ZN(n88) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[47]), .ZN(n9) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[15]), .ZN(n89) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[46]), .ZN(n10) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[14]), .ZN(n92) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[44]), .ZN(n12) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[43]), .ZN(n13) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[11]), .ZN(n65) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[42]), .ZN(n14) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[10]), .ZN(n66) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[41]), .ZN(n15) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[9]), .ZN(n67) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[40]), .ZN(n16) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[8]), .ZN(n68) );
  INVD2BWP30P140 U69 ( .I(n35), .ZN(n29) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[63]), .ZN(n17) );
  INVD2BWP30P140 U71 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[31]), .ZN(n72) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[62]), .ZN(n18) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[30]), .ZN(n73) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[61]), .ZN(n19) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[29]), .ZN(n74) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[60]), .ZN(n20) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[28]), .ZN(n75) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[59]), .ZN(n21) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[27]), .ZN(n76) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[58]), .ZN(n22) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[26]), .ZN(n77) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n23) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n78) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[56]), .ZN(n24) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[24]), .ZN(n79) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[55]), .ZN(n25) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[23]), .ZN(n80) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[54]), .ZN(n26) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[53]), .ZN(n27) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[21]), .ZN(n82) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[52]), .ZN(n28) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[20]), .ZN(n84) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[51]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[19]), .ZN(n85) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n57), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n58), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n64) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n64), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n63) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n63), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n62) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n62), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n61) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n61), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n60) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n60), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n59) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n59), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n91), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n91), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n91), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n91), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n91), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n91), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n91), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  INVD2BWP30P140 U142 ( .I(n71), .ZN(n83) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n83), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n83), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n83), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n83), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n83), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n83), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n83), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n83), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n83), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n83), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n83), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n83), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_44 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n68), .ZN(n91) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n68) );
  OAI22D1BWP30P140 U5 ( .A1(n32), .A2(n15), .B1(n40), .B2(n69), .ZN(N295) );
  OAI22D1BWP30P140 U6 ( .A1(n32), .A2(n16), .B1(n40), .B2(n70), .ZN(N296) );
  OAI22D1BWP30P140 U7 ( .A1(n32), .A2(n14), .B1(n40), .B2(n76), .ZN(N297) );
  OAI22D1BWP30P140 U8 ( .A1(n32), .A2(n13), .B1(n40), .B2(n77), .ZN(N298) );
  OAI22D1BWP30P140 U9 ( .A1(n32), .A2(n12), .B1(n40), .B2(n78), .ZN(N299) );
  OAI22D1BWP30P140 U10 ( .A1(n32), .A2(n11), .B1(n40), .B2(n79), .ZN(N300) );
  OAI22D1BWP30P140 U11 ( .A1(n32), .A2(n10), .B1(n40), .B2(n80), .ZN(N301) );
  OAI22D1BWP30P140 U12 ( .A1(n32), .A2(n9), .B1(n40), .B2(n81), .ZN(N302) );
  OAI22D1BWP30P140 U13 ( .A1(n32), .A2(n8), .B1(n40), .B2(n82), .ZN(N303) );
  OAI22D1BWP30P140 U14 ( .A1(n32), .A2(n7), .B1(n40), .B2(n83), .ZN(N304) );
  OAI22D1BWP30P140 U15 ( .A1(n32), .A2(n6), .B1(n40), .B2(n84), .ZN(N305) );
  OAI22D1BWP30P140 U16 ( .A1(n29), .A2(n28), .B1(n30), .B2(n87), .ZN(N307) );
  OAI22D1BWP30P140 U17 ( .A1(n29), .A2(n27), .B1(n30), .B2(n88), .ZN(N308) );
  OAI22D1BWP30P140 U18 ( .A1(n29), .A2(n26), .B1(n30), .B2(n89), .ZN(N309) );
  OAI22D1BWP30P140 U19 ( .A1(n29), .A2(n25), .B1(n30), .B2(n92), .ZN(N310) );
  OAI22D1BWP30P140 U20 ( .A1(n29), .A2(n24), .B1(n30), .B2(n65), .ZN(N311) );
  OAI22D1BWP30P140 U21 ( .A1(n29), .A2(n23), .B1(n30), .B2(n66), .ZN(N312) );
  OAI22D1BWP30P140 U22 ( .A1(n29), .A2(n22), .B1(n30), .B2(n67), .ZN(N313) );
  OAI22D1BWP30P140 U23 ( .A1(n29), .A2(n21), .B1(n30), .B2(n71), .ZN(N314) );
  OAI22D1BWP30P140 U24 ( .A1(n29), .A2(n20), .B1(n30), .B2(n72), .ZN(N315) );
  OAI22D1BWP30P140 U25 ( .A1(n29), .A2(n19), .B1(n30), .B2(n73), .ZN(N316) );
  OAI22D1BWP30P140 U26 ( .A1(n29), .A2(n18), .B1(n30), .B2(n74), .ZN(N317) );
  OAI22D1BWP30P140 U27 ( .A1(n29), .A2(n17), .B1(n30), .B2(n75), .ZN(N318) );
  ND2OPTIBD1BWP30P140 U28 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U29 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U30 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U31 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U32 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U33 ( .A1(n32), .A2(n31), .B1(n30), .B2(n86), .ZN(N306) );
  INVD1BWP30P140 U34 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U35 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U36 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U38 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U39 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U41 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U42 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[50]), .ZN(n6) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U45 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U46 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U47 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[18]), .ZN(n84) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[49]), .ZN(n7) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[17]), .ZN(n83) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[48]), .ZN(n8) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[16]), .ZN(n82) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[47]), .ZN(n9) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[15]), .ZN(n81) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[46]), .ZN(n10) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[14]), .ZN(n80) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n79) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[44]), .ZN(n12) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[12]), .ZN(n78) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[43]), .ZN(n13) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[11]), .ZN(n77) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[42]), .ZN(n14) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[10]), .ZN(n76) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[40]), .ZN(n15) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[8]), .ZN(n69) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[41]), .ZN(n16) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[9]), .ZN(n70) );
  INVD2BWP30P140 U69 ( .I(n35), .ZN(n29) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[63]), .ZN(n17) );
  INVD2BWP30P140 U71 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[31]), .ZN(n75) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[62]), .ZN(n18) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[30]), .ZN(n74) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[61]), .ZN(n19) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[29]), .ZN(n73) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[60]), .ZN(n20) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[28]), .ZN(n72) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[59]), .ZN(n21) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[27]), .ZN(n71) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[58]), .ZN(n22) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[26]), .ZN(n67) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n23) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n66) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[56]), .ZN(n24) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[24]), .ZN(n65) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[55]), .ZN(n25) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[23]), .ZN(n92) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[54]), .ZN(n26) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[22]), .ZN(n89) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[53]), .ZN(n27) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[21]), .ZN(n88) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[52]), .ZN(n28) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[20]), .ZN(n87) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[51]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[19]), .ZN(n86) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n64), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n63), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n62), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n61), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n60), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n59), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n58), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n57), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n91), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n91), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n91), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n91), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n91), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n91), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n91), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  INVD2BWP30P140 U139 ( .I(n68), .ZN(n85) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n85), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n85), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n85), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n85), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n85), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n85), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n85), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n85), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n85), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n85), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n85), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n85), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_45 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n28), .A2(n16), .B1(n42), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n28), .A2(n15), .B1(n42), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n28), .A2(n14), .B1(n42), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n28), .A2(n13), .B1(n42), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n28), .A2(n12), .B1(n42), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n28), .A2(n11), .B1(n42), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n28), .A2(n10), .B1(n42), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n28), .A2(n9), .B1(n42), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n28), .A2(n8), .B1(n42), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n28), .A2(n7), .B1(n42), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n28), .A2(n6), .B1(n42), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n26), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n25), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n24), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n23), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n22), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n21), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n20), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n19), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n18), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n17), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n31), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n29), .B1(n30), .B2(n92), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n28) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[50]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n42) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[49]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[48]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[47]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[46]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[44]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[43]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[42]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[41]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[40]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD2BWP30P140 U68 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[61]), .ZN(n17) );
  INVD2BWP30P140 U70 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[60]), .ZN(n18) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[59]), .ZN(n19) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[58]), .ZN(n20) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[57]), .ZN(n21) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[56]), .ZN(n22) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[55]), .ZN(n23) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[54]), .ZN(n24) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[53]), .ZN(n25) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[52]), .ZN(n26) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[51]), .ZN(n27) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[19]), .ZN(n77) );
  OAI22D1BWP30P140 U92 ( .A1(n28), .A2(n27), .B1(n30), .B2(n77), .ZN(N306) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[63]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[62]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n42), .A2(n64), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n42), .A2(n63), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n42), .A2(n62), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[34]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n46), .A2(n59), .B1(n45), .B2(n39), .ZN(N289) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[33]), .ZN(n40) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n58), .B1(n45), .B2(n40), .ZN(N288) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[36]), .ZN(n41) );
  OAI22D1BWP30P140 U117 ( .A1(n42), .A2(n61), .B1(n45), .B2(n41), .ZN(N291) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[35]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n60), .B1(n45), .B2(n43), .ZN(N290) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n57), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_46 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n32), .A2(n9), .B1(n46), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n32), .A2(n8), .B1(n46), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n32), .A2(n7), .B1(n46), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n32), .A2(n6), .B1(n46), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n32), .A2(n16), .B1(n46), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n32), .A2(n15), .B1(n46), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n32), .A2(n14), .B1(n46), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n32), .A2(n13), .B1(n46), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n32), .A2(n12), .B1(n46), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n32), .A2(n11), .B1(n46), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n32), .A2(n10), .B1(n46), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n29), .A2(n28), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n29), .A2(n27), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n29), .A2(n26), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n29), .A2(n25), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n29), .A2(n24), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n29), .A2(n23), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n29), .A2(n22), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n29), .A2(n21), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n29), .A2(n20), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n29), .A2(n19), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n29), .A2(n18), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n29), .A2(n17), .B1(n30), .B2(n92), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[43]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n46) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[42]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[41]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[40]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[50]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[49]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[48]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[46]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[45]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[44]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD2BWP30P140 U68 ( .I(n35), .ZN(n29) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[63]), .ZN(n17) );
  INVD2BWP30P140 U70 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[62]), .ZN(n18) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[61]), .ZN(n19) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[60]), .ZN(n20) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[59]), .ZN(n21) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[58]), .ZN(n22) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[57]), .ZN(n23) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[56]), .ZN(n24) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[55]), .ZN(n25) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[54]), .ZN(n26) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[53]), .ZN(n27) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[52]), .ZN(n28) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[51]), .ZN(n31) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[19]), .ZN(n77) );
  OAI22D1BWP30P140 U96 ( .A1(n32), .A2(n31), .B1(n30), .B2(n77), .ZN(N306) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n43) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n43), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[37]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n46), .A2(n62), .B1(n45), .B2(n36), .ZN(N292) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[34]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n43), .A2(n59), .B1(n45), .B2(n37), .ZN(N289) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[33]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n43), .A2(n58), .B1(n45), .B2(n38), .ZN(N288) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[35]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n43), .A2(n60), .B1(n45), .B2(n39), .ZN(N290) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[36]), .ZN(n40) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n61), .B1(n45), .B2(n40), .ZN(N291) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[38]), .ZN(n41) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n63), .B1(n45), .B2(n41), .ZN(N293) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[32]), .ZN(n42) );
  OAI22D1BWP30P140 U120 ( .A1(n43), .A2(n57), .B1(n45), .B2(n42), .ZN(N287) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[39]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N294) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_47 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n71), .ZN(n91) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n71) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n32), .A2(n16), .B1(n46), .B2(n88), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n32), .A2(n15), .B1(n46), .B2(n87), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n32), .A2(n14), .B1(n46), .B2(n86), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n32), .A2(n13), .B1(n46), .B2(n85), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n32), .A2(n12), .B1(n46), .B2(n89), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n32), .A2(n11), .B1(n46), .B2(n92), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n32), .A2(n10), .B1(n46), .B2(n65), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n32), .A2(n9), .B1(n46), .B2(n66), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n32), .A2(n8), .B1(n46), .B2(n67), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n32), .A2(n7), .B1(n46), .B2(n68), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n32), .A2(n6), .B1(n46), .B2(n69), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n29), .A2(n28), .B1(n30), .B2(n72), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n29), .A2(n27), .B1(n30), .B2(n73), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n29), .A2(n26), .B1(n30), .B2(n74), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n29), .A2(n25), .B1(n30), .B2(n75), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n29), .A2(n24), .B1(n30), .B2(n76), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n29), .A2(n23), .B1(n30), .B2(n77), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n29), .A2(n22), .B1(n30), .B2(n78), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n29), .A2(n21), .B1(n30), .B2(n79), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n29), .A2(n20), .B1(n30), .B2(n80), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n29), .A2(n19), .B1(n30), .B2(n81), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n29), .A2(n18), .B1(n30), .B2(n82), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n29), .A2(n17), .B1(n30), .B2(n84), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[50]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n46) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[18]), .ZN(n69) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[49]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[17]), .ZN(n68) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[48]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[16]), .ZN(n67) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[47]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[15]), .ZN(n66) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[46]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[14]), .ZN(n65) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n92) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[44]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[12]), .ZN(n89) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[43]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[11]), .ZN(n85) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[42]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[10]), .ZN(n86) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[41]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[9]), .ZN(n87) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[40]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[8]), .ZN(n88) );
  INVD2BWP30P140 U68 ( .I(n35), .ZN(n29) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[63]), .ZN(n17) );
  INVD2BWP30P140 U70 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[31]), .ZN(n84) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[62]), .ZN(n18) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[30]), .ZN(n82) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[61]), .ZN(n19) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[29]), .ZN(n81) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[60]), .ZN(n20) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[28]), .ZN(n80) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[59]), .ZN(n21) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[27]), .ZN(n79) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[58]), .ZN(n22) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[26]), .ZN(n78) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[57]), .ZN(n23) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[25]), .ZN(n77) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[56]), .ZN(n24) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[24]), .ZN(n76) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[55]), .ZN(n25) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[23]), .ZN(n75) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[54]), .ZN(n26) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[53]), .ZN(n27) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[21]), .ZN(n73) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[52]), .ZN(n28) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[20]), .ZN(n72) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[51]), .ZN(n31) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[19]), .ZN(n70) );
  OAI22D1BWP30P140 U96 ( .A1(n32), .A2(n31), .B1(n30), .B2(n70), .ZN(N306) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n40) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n40), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[32]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n64), .B1(n45), .B2(n36), .ZN(N287) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[33]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n63), .B1(n45), .B2(n37), .ZN(N288) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[34]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n62), .B1(n45), .B2(n38), .ZN(N289) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[35]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n61), .B1(n45), .B2(n39), .ZN(N290) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[36]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n60), .B1(n45), .B2(n41), .ZN(N291) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[37]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n59), .B1(n45), .B2(n42), .ZN(N292) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[39]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n57), .B1(n45), .B2(n43), .ZN(N294) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[38]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n58), .B1(n45), .B2(n44), .ZN(N293) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n91), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n91), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n91), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n91), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n91), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n91), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n91), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U142 ( .I(n71), .ZN(n83) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n83), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n83), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n83), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n83), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n83), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n83), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n83), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n83), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n83), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n83), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n83), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n83), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_48 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n32), .A2(n16), .B1(n46), .B2(n92), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n32), .A2(n15), .B1(n46), .B2(n89), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n32), .A2(n14), .B1(n46), .B2(n88), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n32), .A2(n13), .B1(n46), .B2(n87), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n32), .A2(n12), .B1(n46), .B2(n86), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n32), .A2(n11), .B1(n46), .B2(n85), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n32), .A2(n10), .B1(n46), .B2(n84), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n32), .A2(n9), .B1(n46), .B2(n83), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n32), .A2(n8), .B1(n46), .B2(n82), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n32), .A2(n7), .B1(n46), .B2(n81), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n32), .A2(n6), .B1(n46), .B2(n80), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n29), .A2(n28), .B1(n30), .B2(n77), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n29), .A2(n27), .B1(n30), .B2(n75), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n29), .A2(n26), .B1(n30), .B2(n74), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n29), .A2(n25), .B1(n30), .B2(n73), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n29), .A2(n24), .B1(n30), .B2(n72), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n29), .A2(n23), .B1(n30), .B2(n71), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n29), .A2(n22), .B1(n30), .B2(n70), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n29), .A2(n21), .B1(n30), .B2(n69), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n29), .A2(n20), .B1(n30), .B2(n68), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n29), .A2(n19), .B1(n30), .B2(n67), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n29), .A2(n18), .B1(n30), .B2(n66), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n29), .A2(n17), .B1(n30), .B2(n65), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[50]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n46) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[18]), .ZN(n80) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[49]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[17]), .ZN(n81) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[48]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[16]), .ZN(n82) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[47]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[15]), .ZN(n83) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[46]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[14]), .ZN(n84) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n85) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[44]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[43]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[11]), .ZN(n87) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[42]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[41]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[9]), .ZN(n89) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[40]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[8]), .ZN(n92) );
  INVD2BWP30P140 U68 ( .I(n35), .ZN(n29) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[63]), .ZN(n17) );
  INVD2BWP30P140 U70 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[31]), .ZN(n65) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[62]), .ZN(n18) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[30]), .ZN(n66) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[61]), .ZN(n19) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[29]), .ZN(n67) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[60]), .ZN(n20) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[28]), .ZN(n68) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[59]), .ZN(n21) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[58]), .ZN(n22) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[26]), .ZN(n70) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[57]), .ZN(n23) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[25]), .ZN(n71) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[56]), .ZN(n24) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[24]), .ZN(n72) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[55]), .ZN(n25) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[23]), .ZN(n73) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[54]), .ZN(n26) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[53]), .ZN(n27) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[21]), .ZN(n75) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[52]), .ZN(n28) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[51]), .ZN(n31) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[19]), .ZN(n79) );
  OAI22D1BWP30P140 U96 ( .A1(n32), .A2(n31), .B1(n30), .B2(n79), .ZN(N306) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n40) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n40), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[32]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n64), .B1(n45), .B2(n36), .ZN(N287) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[33]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n63), .B1(n45), .B2(n37), .ZN(N288) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[34]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n62), .B1(n45), .B2(n38), .ZN(N289) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[35]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n61), .B1(n45), .B2(n39), .ZN(N290) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[36]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n60), .B1(n45), .B2(n41), .ZN(N291) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[37]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n59), .B1(n45), .B2(n42), .ZN(N292) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[38]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n58), .B1(n45), .B2(n43), .ZN(N293) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[39]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n57), .B1(n45), .B2(n44), .ZN(N294) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_49 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n75), .ZN(n91) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n75) );
  OAI22D1BWP30P140 U5 ( .A1(n20), .A2(n19), .B1(n30), .B2(n89), .ZN(N306) );
  ND2OPTIBD1BWP30P140 U6 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U7 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U8 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U9 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U10 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U11 ( .A1(n20), .A2(n16), .B1(n46), .B2(n74), .ZN(N295) );
  OAI22D1BWP30P140 U12 ( .A1(n20), .A2(n15), .B1(n46), .B2(n73), .ZN(N296) );
  OAI22D1BWP30P140 U13 ( .A1(n20), .A2(n14), .B1(n46), .B2(n72), .ZN(N297) );
  OAI22D1BWP30P140 U14 ( .A1(n20), .A2(n13), .B1(n46), .B2(n71), .ZN(N298) );
  OAI22D1BWP30P140 U15 ( .A1(n20), .A2(n12), .B1(n46), .B2(n70), .ZN(N299) );
  OAI22D1BWP30P140 U16 ( .A1(n20), .A2(n11), .B1(n46), .B2(n69), .ZN(N300) );
  OAI22D1BWP30P140 U17 ( .A1(n20), .A2(n10), .B1(n46), .B2(n68), .ZN(N301) );
  OAI22D1BWP30P140 U18 ( .A1(n20), .A2(n9), .B1(n46), .B2(n67), .ZN(N302) );
  OAI22D1BWP30P140 U19 ( .A1(n20), .A2(n8), .B1(n46), .B2(n66), .ZN(N303) );
  OAI22D1BWP30P140 U20 ( .A1(n20), .A2(n7), .B1(n46), .B2(n65), .ZN(N304) );
  OAI22D1BWP30P140 U21 ( .A1(n20), .A2(n6), .B1(n46), .B2(n92), .ZN(N305) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n18), .B1(n30), .B2(n88), .ZN(N307) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n17), .B1(n30), .B2(n86), .ZN(N308) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n21), .B1(n30), .B2(n85), .ZN(N309) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n31), .B1(n30), .B2(n84), .ZN(N310) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n29), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n28), .B1(n30), .B2(n82), .ZN(N312) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n27), .B1(n30), .B2(n81), .ZN(N313) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n26), .B1(n30), .B2(n80), .ZN(N314) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n25), .B1(n30), .B2(n79), .ZN(N315) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n24), .B1(n30), .B2(n78), .ZN(N316) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n23), .B1(n30), .B2(n77), .ZN(N317) );
  OAI22D1BWP30P140 U33 ( .A1(n32), .A2(n22), .B1(n30), .B2(n76), .ZN(N318) );
  INVD1BWP30P140 U34 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U35 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U36 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U38 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U39 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U41 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U42 ( .I(n35), .ZN(n20) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[50]), .ZN(n6) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U45 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U46 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U47 ( .I(n33), .ZN(n46) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[18]), .ZN(n92) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[49]), .ZN(n7) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[17]), .ZN(n65) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[48]), .ZN(n8) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[16]), .ZN(n66) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[47]), .ZN(n9) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[15]), .ZN(n67) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[46]), .ZN(n10) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[14]), .ZN(n68) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n69) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[44]), .ZN(n12) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[12]), .ZN(n70) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[43]), .ZN(n13) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[11]), .ZN(n71) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[42]), .ZN(n14) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[10]), .ZN(n72) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[41]), .ZN(n15) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[9]), .ZN(n73) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[40]), .ZN(n16) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[8]), .ZN(n74) );
  INVD2BWP30P140 U69 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[53]), .ZN(n17) );
  INVD2BWP30P140 U71 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[21]), .ZN(n86) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n18) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n88) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[51]), .ZN(n19) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[19]), .ZN(n89) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n85) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[63]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[31]), .ZN(n76) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[62]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[30]), .ZN(n77) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[61]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[29]), .ZN(n78) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[60]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[28]), .ZN(n79) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n80) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[58]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[26]), .ZN(n81) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[57]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[25]), .ZN(n82) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[56]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[55]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[23]), .ZN(n84) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n40) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n40), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[32]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n64), .B1(n45), .B2(n36), .ZN(N287) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[33]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n63), .B1(n45), .B2(n37), .ZN(N288) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[34]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n62), .B1(n45), .B2(n38), .ZN(N289) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[35]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n61), .B1(n45), .B2(n39), .ZN(N290) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[36]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n60), .B1(n45), .B2(n41), .ZN(N291) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[37]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n59), .B1(n45), .B2(n42), .ZN(N292) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[38]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n58), .B1(n45), .B2(n43), .ZN(N293) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[39]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n57), .B1(n45), .B2(n44), .ZN(N294) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n91), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n91), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n91), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n91), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n91), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n91), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n91), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  INVD2BWP30P140 U146 ( .I(n75), .ZN(n87) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n87), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n87), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n87), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n87), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n87), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n87), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n87), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n87), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n87), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U156 ( .A1(n85), .A2(n87), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U157 ( .A1(n86), .A2(n87), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n87), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_50 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n74), .ZN(n91) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n74) );
  OAI22D1BWP30P140 U5 ( .A1(n32), .A2(n31), .B1(n30), .B2(n88), .ZN(N306) );
  ND2OPTIBD1BWP30P140 U6 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U7 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U8 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U9 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U10 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U11 ( .A1(n32), .A2(n16), .B1(n46), .B2(n73), .ZN(N295) );
  OAI22D1BWP30P140 U12 ( .A1(n32), .A2(n15), .B1(n46), .B2(n72), .ZN(N296) );
  OAI22D1BWP30P140 U13 ( .A1(n32), .A2(n14), .B1(n46), .B2(n71), .ZN(N297) );
  OAI22D1BWP30P140 U14 ( .A1(n32), .A2(n13), .B1(n46), .B2(n70), .ZN(N298) );
  OAI22D1BWP30P140 U15 ( .A1(n32), .A2(n12), .B1(n46), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U16 ( .A1(n32), .A2(n11), .B1(n46), .B2(n68), .ZN(N300) );
  OAI22D1BWP30P140 U17 ( .A1(n32), .A2(n10), .B1(n46), .B2(n67), .ZN(N301) );
  OAI22D1BWP30P140 U18 ( .A1(n32), .A2(n9), .B1(n46), .B2(n66), .ZN(N302) );
  OAI22D1BWP30P140 U19 ( .A1(n32), .A2(n8), .B1(n46), .B2(n65), .ZN(N303) );
  OAI22D1BWP30P140 U20 ( .A1(n32), .A2(n7), .B1(n46), .B2(n92), .ZN(N304) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n6), .B1(n46), .B2(n89), .ZN(N305) );
  OAI22D1BWP30P140 U22 ( .A1(n29), .A2(n28), .B1(n30), .B2(n87), .ZN(N307) );
  OAI22D1BWP30P140 U23 ( .A1(n29), .A2(n27), .B1(n30), .B2(n85), .ZN(N308) );
  OAI22D1BWP30P140 U24 ( .A1(n29), .A2(n26), .B1(n30), .B2(n84), .ZN(N309) );
  OAI22D1BWP30P140 U25 ( .A1(n29), .A2(n25), .B1(n30), .B2(n83), .ZN(N310) );
  OAI22D1BWP30P140 U26 ( .A1(n29), .A2(n24), .B1(n30), .B2(n82), .ZN(N311) );
  OAI22D1BWP30P140 U27 ( .A1(n29), .A2(n23), .B1(n30), .B2(n81), .ZN(N312) );
  OAI22D1BWP30P140 U28 ( .A1(n29), .A2(n22), .B1(n30), .B2(n80), .ZN(N313) );
  OAI22D1BWP30P140 U29 ( .A1(n29), .A2(n21), .B1(n30), .B2(n79), .ZN(N314) );
  OAI22D1BWP30P140 U30 ( .A1(n29), .A2(n20), .B1(n30), .B2(n78), .ZN(N315) );
  OAI22D1BWP30P140 U31 ( .A1(n29), .A2(n19), .B1(n30), .B2(n77), .ZN(N316) );
  OAI22D1BWP30P140 U32 ( .A1(n29), .A2(n18), .B1(n30), .B2(n76), .ZN(N317) );
  OAI22D1BWP30P140 U33 ( .A1(n29), .A2(n17), .B1(n30), .B2(n75), .ZN(N318) );
  INVD1BWP30P140 U34 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U35 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U36 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U38 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U39 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U41 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U42 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[50]), .ZN(n6) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U45 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U46 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U47 ( .I(n33), .ZN(n46) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[18]), .ZN(n89) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[49]), .ZN(n7) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[17]), .ZN(n92) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[48]), .ZN(n8) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[16]), .ZN(n65) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[47]), .ZN(n9) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[15]), .ZN(n66) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[46]), .ZN(n10) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[14]), .ZN(n67) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n68) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[44]), .ZN(n12) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[43]), .ZN(n13) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[11]), .ZN(n70) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[42]), .ZN(n14) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[10]), .ZN(n71) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[41]), .ZN(n15) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[9]), .ZN(n72) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[40]), .ZN(n16) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[8]), .ZN(n73) );
  INVD2BWP30P140 U69 ( .I(n35), .ZN(n29) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[63]), .ZN(n17) );
  INVD2BWP30P140 U71 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[31]), .ZN(n75) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[62]), .ZN(n18) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[30]), .ZN(n76) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[61]), .ZN(n19) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[29]), .ZN(n77) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[60]), .ZN(n20) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[28]), .ZN(n78) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[59]), .ZN(n21) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[27]), .ZN(n79) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[58]), .ZN(n22) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[26]), .ZN(n80) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n23) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n81) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[56]), .ZN(n24) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[24]), .ZN(n82) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[55]), .ZN(n25) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[23]), .ZN(n83) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[54]), .ZN(n26) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[22]), .ZN(n84) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[53]), .ZN(n27) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[21]), .ZN(n85) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[52]), .ZN(n28) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[20]), .ZN(n87) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[51]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[19]), .ZN(n88) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n40) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n40), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[32]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n64), .B1(n45), .B2(n36), .ZN(N287) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[33]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n63), .B1(n45), .B2(n37), .ZN(N288) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[34]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n62), .B1(n45), .B2(n38), .ZN(N289) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[35]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n61), .B1(n45), .B2(n39), .ZN(N290) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[36]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n60), .B1(n45), .B2(n41), .ZN(N291) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[37]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n59), .B1(n45), .B2(n42), .ZN(N292) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[38]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n58), .B1(n45), .B2(n43), .ZN(N293) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[39]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n57), .B1(n45), .B2(n44), .ZN(N294) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n91), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n91), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n91), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n91), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n91), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n91), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n91), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  INVD2BWP30P140 U145 ( .I(n74), .ZN(n86) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n86), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n86), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n86), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n86), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n86), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n86), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n86), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n86), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n86), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n86), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U156 ( .A1(n85), .A2(n86), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n86), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_51 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n67), .ZN(n82) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n67) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n6), .B1(n46), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n7), .B1(n46), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n8), .B1(n46), .B2(n83), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n9), .B1(n46), .B2(n81), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n10), .B1(n46), .B2(n80), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n11), .B1(n46), .B2(n79), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n12), .B1(n46), .B2(n78), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n13), .B1(n46), .B2(n77), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n14), .B1(n46), .B2(n76), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n15), .B1(n46), .B2(n75), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n16), .B1(n46), .B2(n74), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n19), .B1(n30), .B2(n72), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n20), .B1(n30), .B2(n71), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n21), .B1(n30), .B2(n70), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n22), .B1(n30), .B2(n69), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n23), .B1(n30), .B2(n68), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n24), .B1(n30), .B2(n92), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n25), .B1(n30), .B2(n89), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n26), .B1(n30), .B2(n88), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n27), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n28), .B1(n30), .B2(n86), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n29), .B1(n30), .B2(n85), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n31), .B1(n30), .B2(n84), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n46) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[10]), .ZN(n83) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[11]), .ZN(n81) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n80) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n79) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[14]), .ZN(n78) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n77) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[16]), .ZN(n76) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[17]), .ZN(n75) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[18]), .ZN(n74) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n73) );
  OAI22D1BWP30P140 U71 ( .A1(n18), .A2(n17), .B1(n30), .B2(n73), .ZN(N306) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n72) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n71) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n70) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n69) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n68) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n92) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n89) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n88) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n86) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n85) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n84) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n43) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n43), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[6]), .ZN(n64) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[38]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n46), .A2(n64), .B1(n45), .B2(n36), .ZN(N293) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[37]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n46), .A2(n62), .B1(n45), .B2(n37), .ZN(N292) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[36]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n46), .A2(n61), .B1(n45), .B2(n38), .ZN(N291) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[3]), .ZN(n59) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[35]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n43), .A2(n59), .B1(n45), .B2(n39), .ZN(N290) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[34]), .ZN(n40) );
  OAI22D1BWP30P140 U114 ( .A1(n43), .A2(n60), .B1(n45), .B2(n40), .ZN(N289) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[33]), .ZN(n41) );
  OAI22D1BWP30P140 U117 ( .A1(n43), .A2(n58), .B1(n45), .B2(n41), .ZN(N288) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[32]), .ZN(n42) );
  OAI22D1BWP30P140 U120 ( .A1(n43), .A2(n57), .B1(n45), .B2(n42), .ZN(N287) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[7]), .ZN(n63) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[39]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n63), .B1(n45), .B2(n44), .ZN(N294) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n82), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n82), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n82), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n82), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n82), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n82), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n82), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n82), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n82), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n82), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  INVD2BWP30P140 U138 ( .I(n67), .ZN(n91) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n82), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n82), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n82), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n82), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n82), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n82), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n82), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n82), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n82), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n82), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_52 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n6), .B1(n40), .B2(n92), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n7), .B1(n40), .B2(n89), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n8), .B1(n40), .B2(n88), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n9), .B1(n40), .B2(n87), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n10), .B1(n40), .B2(n86), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n11), .B1(n40), .B2(n85), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n12), .B1(n40), .B2(n84), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n13), .B1(n40), .B2(n83), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n14), .B1(n40), .B2(n82), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n15), .B1(n40), .B2(n81), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n16), .B1(n40), .B2(n80), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n19), .B1(n30), .B2(n77), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n20), .B1(n30), .B2(n75), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n21), .B1(n30), .B2(n74), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n22), .B1(n30), .B2(n73), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n23), .B1(n30), .B2(n72), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n24), .B1(n30), .B2(n71), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n25), .B1(n30), .B2(n70), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n26), .B1(n30), .B2(n69), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n27), .B1(n30), .B2(n68), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n28), .B1(n30), .B2(n67), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n29), .B1(n30), .B2(n66), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n31), .B1(n30), .B2(n65), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[8]), .ZN(n92) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[9]), .ZN(n89) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[11]), .ZN(n87) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n85) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[14]), .ZN(n84) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n83) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[16]), .ZN(n82) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[17]), .ZN(n81) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[18]), .ZN(n80) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n79) );
  OAI22D1BWP30P140 U71 ( .A1(n18), .A2(n17), .B1(n30), .B2(n79), .ZN(N306) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n75) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n73) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n72) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n71) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n70) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n68) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n67) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n66) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n65) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n57), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n58), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n59), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n60), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n61), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n62), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n63), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_53 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n66), .ZN(n91) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n66) );
  OAI22D1BWP30P140 U5 ( .A1(n18), .A2(n6), .B1(n40), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U6 ( .A1(n18), .A2(n7), .B1(n40), .B2(n92), .ZN(N296) );
  OAI22D1BWP30P140 U7 ( .A1(n18), .A2(n8), .B1(n40), .B2(n87), .ZN(N297) );
  OAI22D1BWP30P140 U8 ( .A1(n18), .A2(n9), .B1(n40), .B2(n86), .ZN(N298) );
  OAI22D1BWP30P140 U9 ( .A1(n18), .A2(n10), .B1(n40), .B2(n85), .ZN(N299) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n11), .B1(n40), .B2(n84), .ZN(N300) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n12), .B1(n40), .B2(n83), .ZN(N301) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n13), .B1(n40), .B2(n82), .ZN(N302) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n14), .B1(n40), .B2(n81), .ZN(N303) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n15), .B1(n40), .B2(n80), .ZN(N304) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n16), .B1(n40), .B2(n79), .ZN(N305) );
  OAI22D1BWP30P140 U16 ( .A1(n32), .A2(n19), .B1(n30), .B2(n77), .ZN(N307) );
  OAI22D1BWP30P140 U17 ( .A1(n32), .A2(n20), .B1(n30), .B2(n76), .ZN(N308) );
  OAI22D1BWP30P140 U18 ( .A1(n32), .A2(n21), .B1(n30), .B2(n75), .ZN(N309) );
  OAI22D1BWP30P140 U19 ( .A1(n32), .A2(n22), .B1(n30), .B2(n74), .ZN(N310) );
  OAI22D1BWP30P140 U20 ( .A1(n32), .A2(n23), .B1(n30), .B2(n73), .ZN(N311) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n24), .B1(n30), .B2(n72), .ZN(N312) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n25), .B1(n30), .B2(n71), .ZN(N313) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n26), .B1(n30), .B2(n70), .ZN(N314) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n27), .B1(n30), .B2(n69), .ZN(N315) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n28), .B1(n30), .B2(n68), .ZN(N316) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n29), .B1(n30), .B2(n67), .ZN(N317) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n31), .B1(n30), .B2(n89), .ZN(N318) );
  ND2OPTIBD1BWP30P140 U28 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U29 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U30 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U31 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U32 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U33 ( .A1(n18), .A2(n17), .B1(n30), .B2(n78), .ZN(N306) );
  INVD1BWP30P140 U34 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U35 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U36 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U38 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U39 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U41 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U42 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U45 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U46 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U47 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n92) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n87) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n86) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n85) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n84) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[14]), .ZN(n83) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[15]), .ZN(n82) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n81) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n80) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n79) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U70 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n76) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n75) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n74) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n73) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n72) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n71) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n70) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n69) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n68) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n67) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n89) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n61) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n61), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n62) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n62), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n63) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n63), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n64) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n64), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n60), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n59), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n58), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n57), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n91), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n91), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n91), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n91), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n91), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n91), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n91), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  INVD2BWP30P140 U137 ( .I(n66), .ZN(n88) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n88), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n88), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n88), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n88), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n88), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n88), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n88), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n88), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n88), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n88), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n88), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n85), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n86), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n87), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n88), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_54 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  OAI22D1BWP30P140 U5 ( .A1(n18), .A2(n6), .B1(n40), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U6 ( .A1(n18), .A2(n7), .B1(n40), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U7 ( .A1(n18), .A2(n8), .B1(n40), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U8 ( .A1(n18), .A2(n9), .B1(n40), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U9 ( .A1(n18), .A2(n10), .B1(n40), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n11), .B1(n40), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n12), .B1(n40), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n13), .B1(n40), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n14), .B1(n40), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n15), .B1(n40), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n16), .B1(n40), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U16 ( .A1(n32), .A2(n19), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U17 ( .A1(n32), .A2(n20), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U18 ( .A1(n32), .A2(n21), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U19 ( .A1(n32), .A2(n22), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U20 ( .A1(n32), .A2(n23), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n24), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n25), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n26), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n27), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n28), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n29), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n31), .B1(n30), .B2(n92), .ZN(N318) );
  ND2OPTIBD1BWP30P140 U28 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U29 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U30 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U31 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U32 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U33 ( .A1(n18), .A2(n17), .B1(n30), .B2(n77), .ZN(N306) );
  INVD1BWP30P140 U34 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U35 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U36 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U38 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U39 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U41 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U42 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U45 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U46 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U47 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U70 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n77) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n57), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n58), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n59), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n60), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n61), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n62), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n63), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_55 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n67), .ZN(n91) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n67) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n6), .B1(n40), .B2(n68), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n7), .B1(n40), .B2(n69), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n8), .B1(n40), .B2(n70), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n9), .B1(n40), .B2(n71), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n10), .B1(n40), .B2(n72), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n11), .B1(n40), .B2(n73), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n12), .B1(n40), .B2(n74), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n13), .B1(n40), .B2(n75), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n14), .B1(n40), .B2(n76), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n15), .B1(n40), .B2(n77), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n16), .B1(n40), .B2(n78), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n19), .B1(n30), .B2(n81), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n20), .B1(n30), .B2(n82), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n21), .B1(n30), .B2(n83), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n22), .B1(n30), .B2(n84), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n23), .B1(n30), .B2(n85), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n24), .B1(n30), .B2(n86), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n25), .B1(n30), .B2(n87), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n26), .B1(n30), .B2(n88), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n27), .B1(n30), .B2(n89), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n28), .B1(n30), .B2(n92), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n29), .B1(n30), .B2(n65), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n31), .B1(n30), .B2(n66), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[8]), .ZN(n68) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[9]), .ZN(n69) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[10]), .ZN(n70) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[11]), .ZN(n71) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n72) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n73) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[14]), .ZN(n74) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n75) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[16]), .ZN(n76) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[17]), .ZN(n77) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[18]), .ZN(n78) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n80) );
  OAI22D1BWP30P140 U71 ( .A1(n18), .A2(n17), .B1(n30), .B2(n80), .ZN(N306) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n81) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n82) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n83) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n84) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n85) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n86) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n87) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n88) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n89) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n92) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n65) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n66) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n57), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n64) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n64), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n63) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n63), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n62), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n61), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n60), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n59), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n58) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n58), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n91), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n91), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n91), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n91), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n91), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n91), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n91), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  INVD2BWP30P140 U138 ( .I(n67), .ZN(n79) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n79), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n79), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n79), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n79), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n79), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n79), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n79), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n79), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n79), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n79), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n79), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n79), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_56 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n6), .B1(n40), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n7), .B1(n40), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n8), .B1(n40), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n9), .B1(n40), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n10), .B1(n40), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n11), .B1(n40), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n12), .B1(n40), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n13), .B1(n40), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n14), .B1(n40), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n15), .B1(n40), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n16), .B1(n40), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n19), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n20), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n21), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n22), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n23), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n24), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n25), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n26), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n27), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n28), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n29), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n31), .B1(n30), .B2(n92), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n77) );
  OAI22D1BWP30P140 U71 ( .A1(n18), .A2(n17), .B1(n30), .B2(n77), .ZN(N306) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n64), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n63), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n62), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n61), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n60), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n59), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n58), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n57), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_57 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  OAI22D1BWP30P140 U5 ( .A1(n18), .A2(n17), .B1(n30), .B2(n77), .ZN(N306) );
  ND2OPTIBD1BWP30P140 U6 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U7 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U8 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U9 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U10 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n6), .B1(n46), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n7), .B1(n46), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n8), .B1(n46), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n9), .B1(n46), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n10), .B1(n46), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n11), .B1(n46), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n12), .B1(n46), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n13), .B1(n46), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n14), .B1(n46), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n15), .B1(n46), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U21 ( .A1(n18), .A2(n16), .B1(n46), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n19), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n20), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n21), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n22), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n23), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n24), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n25), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n26), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n27), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n28), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n29), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U33 ( .A1(n32), .A2(n31), .B1(n30), .B2(n92), .ZN(N318) );
  INVD1BWP30P140 U34 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U35 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U36 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U38 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U39 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U41 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U42 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U45 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U46 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U47 ( .I(n33), .ZN(n46) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U70 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n77) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n43) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n43), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[38]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n46), .A2(n63), .B1(n45), .B2(n36), .ZN(N293) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[37]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n46), .A2(n62), .B1(n45), .B2(n37), .ZN(N292) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[36]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n46), .A2(n61), .B1(n45), .B2(n38), .ZN(N291) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[35]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n43), .A2(n60), .B1(n45), .B2(n39), .ZN(N290) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[34]), .ZN(n40) );
  OAI22D1BWP30P140 U114 ( .A1(n43), .A2(n59), .B1(n45), .B2(n40), .ZN(N289) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[33]), .ZN(n41) );
  OAI22D1BWP30P140 U117 ( .A1(n43), .A2(n58), .B1(n45), .B2(n41), .ZN(N288) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[32]), .ZN(n42) );
  OAI22D1BWP30P140 U120 ( .A1(n43), .A2(n57), .B1(n45), .B2(n42), .ZN(N287) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[39]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N294) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_58 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  OAI22D1BWP30P140 U5 ( .A1(n18), .A2(n17), .B1(n30), .B2(n77), .ZN(N306) );
  ND2OPTIBD1BWP30P140 U6 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U7 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U8 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U9 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U10 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n6), .B1(n40), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n7), .B1(n40), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n8), .B1(n40), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n9), .B1(n40), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n10), .B1(n40), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n11), .B1(n40), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n12), .B1(n40), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n13), .B1(n40), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n14), .B1(n40), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n15), .B1(n40), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U21 ( .A1(n18), .A2(n16), .B1(n40), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n19), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n20), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n21), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n22), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n23), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n24), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n25), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n26), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n27), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n28), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n29), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U33 ( .A1(n32), .A2(n31), .B1(n30), .B2(n92), .ZN(N318) );
  INVD1BWP30P140 U34 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U35 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U36 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U38 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U39 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U41 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U42 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U45 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U46 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U47 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U70 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n77) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n64), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n63), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n60) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n60), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n62), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n61), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n59), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n58), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n57), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_59 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n71), .ZN(n91) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n71) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n6), .B1(n40), .B2(n85), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n7), .B1(n40), .B2(n86), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n8), .B1(n40), .B2(n87), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n9), .B1(n40), .B2(n88), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n10), .B1(n40), .B2(n89), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n11), .B1(n40), .B2(n92), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n12), .B1(n40), .B2(n65), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n13), .B1(n40), .B2(n66), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n14), .B1(n40), .B2(n67), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n15), .B1(n40), .B2(n68), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n16), .B1(n40), .B2(n69), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n19), .B1(n30), .B2(n72), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n20), .B1(n30), .B2(n73), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n21), .B1(n30), .B2(n74), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n22), .B1(n30), .B2(n75), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n23), .B1(n30), .B2(n76), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n24), .B1(n30), .B2(n77), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n25), .B1(n30), .B2(n78), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n26), .B1(n30), .B2(n79), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n27), .B1(n30), .B2(n80), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n28), .B1(n30), .B2(n81), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n29), .B1(n30), .B2(n82), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n31), .B1(n30), .B2(n84), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[8]), .ZN(n85) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[9]), .ZN(n86) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[10]), .ZN(n87) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[11]), .ZN(n88) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n89) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n92) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[14]), .ZN(n65) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n66) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[16]), .ZN(n67) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[17]), .ZN(n68) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[18]), .ZN(n69) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n70) );
  OAI22D1BWP30P140 U71 ( .A1(n18), .A2(n17), .B1(n30), .B2(n70), .ZN(N306) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n72) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n73) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n75) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n76) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n77) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n78) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n79) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n80) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n81) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n82) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n84) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n64), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n63), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n62), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n61), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n60), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n59), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n58), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n57), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n91), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n91), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n91), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n91), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n91), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n91), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n91), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U142 ( .I(n71), .ZN(n83) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n83), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n83), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n83), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n83), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n83), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n83), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n83), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n83), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n83), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n83), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n83), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n83), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_60 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n28), .A2(n6), .B1(n40), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n28), .A2(n7), .B1(n40), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n28), .A2(n8), .B1(n40), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n28), .A2(n9), .B1(n40), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n28), .A2(n10), .B1(n40), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n28), .A2(n11), .B1(n40), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n28), .A2(n12), .B1(n40), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n28), .A2(n13), .B1(n40), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n28), .A2(n14), .B1(n40), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n28), .A2(n15), .B1(n40), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n28), .A2(n16), .B1(n40), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n29), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n31), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n26), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n17), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n18), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n19), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n20), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n21), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n22), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n23), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n24), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n25), .B1(n30), .B2(n92), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n28) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD2BWP30P140 U68 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[55]), .ZN(n17) );
  INVD2BWP30P140 U70 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[56]), .ZN(n18) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[57]), .ZN(n19) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[58]), .ZN(n20) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[59]), .ZN(n21) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[60]), .ZN(n22) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[61]), .ZN(n23) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[62]), .ZN(n24) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[63]), .ZN(n25) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[54]), .ZN(n26) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[51]), .ZN(n27) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[19]), .ZN(n77) );
  OAI22D1BWP30P140 U92 ( .A1(n28), .A2(n27), .B1(n30), .B2(n77), .ZN(N306) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[52]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[53]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n57), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n58), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n59), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n60), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n61), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n62), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n63), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_61 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  OAI22D1BWP30P140 U5 ( .A1(n18), .A2(n6), .B1(n40), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U6 ( .A1(n18), .A2(n7), .B1(n40), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U7 ( .A1(n18), .A2(n8), .B1(n40), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U8 ( .A1(n18), .A2(n9), .B1(n40), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U9 ( .A1(n18), .A2(n10), .B1(n40), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n11), .B1(n40), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n12), .B1(n40), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n13), .B1(n40), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n14), .B1(n40), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n15), .B1(n40), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n16), .B1(n40), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U16 ( .A1(n32), .A2(n19), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U17 ( .A1(n32), .A2(n20), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U18 ( .A1(n32), .A2(n21), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U19 ( .A1(n32), .A2(n22), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U20 ( .A1(n32), .A2(n23), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n24), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n25), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n26), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n27), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n28), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n29), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n31), .B1(n30), .B2(n92), .ZN(N318) );
  ND2OPTIBD1BWP30P140 U28 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U29 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U30 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U31 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U32 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U33 ( .A1(n18), .A2(n17), .B1(n30), .B2(n77), .ZN(N306) );
  INVD1BWP30P140 U34 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U35 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U36 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U38 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U39 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U41 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U42 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U45 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U46 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U47 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U70 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n77) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n64), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n63), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n62), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n61), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n60), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n59), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n58), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n57), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_62 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  OAI22D1BWP30P140 U5 ( .A1(n18), .A2(n6), .B1(n40), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U6 ( .A1(n18), .A2(n7), .B1(n40), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U7 ( .A1(n18), .A2(n8), .B1(n40), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U8 ( .A1(n18), .A2(n9), .B1(n40), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U9 ( .A1(n18), .A2(n10), .B1(n40), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n11), .B1(n40), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n12), .B1(n40), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n13), .B1(n40), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n14), .B1(n40), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n15), .B1(n40), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n16), .B1(n40), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U16 ( .A1(n32), .A2(n19), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U17 ( .A1(n32), .A2(n20), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U18 ( .A1(n32), .A2(n21), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U19 ( .A1(n32), .A2(n22), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U20 ( .A1(n32), .A2(n23), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n24), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n25), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n26), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n27), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n28), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n29), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n31), .B1(n30), .B2(n92), .ZN(N318) );
  ND2OPTIBD1BWP30P140 U28 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U29 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U30 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U31 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U32 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U33 ( .A1(n18), .A2(n17), .B1(n30), .B2(n77), .ZN(N306) );
  INVD1BWP30P140 U34 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U35 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U36 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U38 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U39 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U41 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U42 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U45 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U46 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U47 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U70 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n77) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n62) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n62), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n61) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n61), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n64) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n64), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n63) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n63), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n59) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n59), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n60), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n58), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n57), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_63 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n16), .B1(n40), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n15), .B1(n40), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n14), .B1(n40), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n13), .B1(n40), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n6), .B1(n40), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n7), .B1(n40), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n8), .B1(n40), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n9), .B1(n40), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n10), .B1(n40), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n11), .B1(n40), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n12), .B1(n40), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n19), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n20), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n21), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n22), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n23), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n24), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n25), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n26), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n27), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n28), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n29), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n31), .B1(n30), .B2(n92), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[44]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[45]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[46]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[47]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[48]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[49]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[50]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[43]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[42]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[41]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[40]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n77) );
  OAI22D1BWP30P140 U71 ( .A1(n18), .A2(n17), .B1(n30), .B2(n77), .ZN(N306) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n64), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n63), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n62), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n61), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n60), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n59), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n58), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n57), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_64 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n6), .B1(n40), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n7), .B1(n40), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n8), .B1(n40), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n9), .B1(n40), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n10), .B1(n40), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n11), .B1(n40), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n12), .B1(n40), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n13), .B1(n40), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n14), .B1(n40), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n15), .B1(n40), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n16), .B1(n40), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n19), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n20), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n21), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n22), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n23), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n24), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n25), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n26), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n27), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n28), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n29), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n31), .B1(n30), .B2(n92), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n77) );
  OAI22D1BWP30P140 U71 ( .A1(n18), .A2(n17), .B1(n30), .B2(n77), .ZN(N306) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n64), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n63), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n62), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n61), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n60), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n59), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n58), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n57), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_65 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  OAI22D1BWP30P140 U5 ( .A1(n18), .A2(n6), .B1(n40), .B2(n92), .ZN(N295) );
  OAI22D1BWP30P140 U6 ( .A1(n18), .A2(n7), .B1(n40), .B2(n89), .ZN(N296) );
  OAI22D1BWP30P140 U7 ( .A1(n18), .A2(n8), .B1(n40), .B2(n88), .ZN(N297) );
  OAI22D1BWP30P140 U8 ( .A1(n18), .A2(n9), .B1(n40), .B2(n87), .ZN(N298) );
  OAI22D1BWP30P140 U9 ( .A1(n18), .A2(n10), .B1(n40), .B2(n86), .ZN(N299) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n11), .B1(n40), .B2(n85), .ZN(N300) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n12), .B1(n40), .B2(n84), .ZN(N301) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n13), .B1(n40), .B2(n83), .ZN(N302) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n14), .B1(n40), .B2(n82), .ZN(N303) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n15), .B1(n40), .B2(n81), .ZN(N304) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n16), .B1(n40), .B2(n80), .ZN(N305) );
  OAI22D1BWP30P140 U16 ( .A1(n32), .A2(n19), .B1(n30), .B2(n77), .ZN(N307) );
  OAI22D1BWP30P140 U17 ( .A1(n32), .A2(n20), .B1(n30), .B2(n75), .ZN(N308) );
  OAI22D1BWP30P140 U18 ( .A1(n32), .A2(n21), .B1(n30), .B2(n74), .ZN(N309) );
  OAI22D1BWP30P140 U19 ( .A1(n32), .A2(n22), .B1(n30), .B2(n73), .ZN(N310) );
  OAI22D1BWP30P140 U20 ( .A1(n32), .A2(n23), .B1(n30), .B2(n72), .ZN(N311) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n24), .B1(n30), .B2(n71), .ZN(N312) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n25), .B1(n30), .B2(n70), .ZN(N313) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n26), .B1(n30), .B2(n69), .ZN(N314) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n27), .B1(n30), .B2(n68), .ZN(N315) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n28), .B1(n30), .B2(n67), .ZN(N316) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n29), .B1(n30), .B2(n66), .ZN(N317) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n31), .B1(n30), .B2(n65), .ZN(N318) );
  ND2OPTIBD1BWP30P140 U28 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U29 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U30 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U31 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U32 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U33 ( .A1(n18), .A2(n17), .B1(n30), .B2(n79), .ZN(N306) );
  INVD1BWP30P140 U34 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U35 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U36 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U38 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U39 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U41 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U42 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U45 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U46 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U47 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n92) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n89) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n87) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n85) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[14]), .ZN(n84) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[15]), .ZN(n83) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n82) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n81) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n80) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U70 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n79) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n75) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n73) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n72) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n71) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n70) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n68) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n67) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n66) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n65) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n57), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n58), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n59), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n60), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n61), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n62), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n63), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_66 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n69), .ZN(n85) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n69) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n26), .A2(n14), .B1(n40), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n26), .A2(n16), .B1(n40), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n26), .A2(n13), .B1(n40), .B2(n68), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n26), .A2(n11), .B1(n40), .B2(n78), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n26), .A2(n15), .B1(n40), .B2(n79), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n26), .A2(n9), .B1(n40), .B2(n67), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n26), .A2(n6), .B1(n40), .B2(n86), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n26), .A2(n7), .B1(n40), .B2(n84), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n26), .A2(n10), .B1(n40), .B2(n83), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n26), .A2(n8), .B1(n40), .B2(n82), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n26), .A2(n12), .B1(n40), .B2(n81), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n22), .B1(n30), .B2(n77), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n23), .B1(n30), .B2(n76), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n31), .B1(n30), .B2(n75), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n24), .B1(n30), .B2(n74), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n28), .B1(n30), .B2(n73), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n27), .B1(n30), .B2(n72), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n29), .B1(n30), .B2(n71), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n21), .B1(n30), .B2(n70), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n17), .B1(n30), .B2(n92), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n18), .B1(n30), .B2(n89), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n19), .B1(n30), .B2(n88), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n20), .B1(n30), .B2(n87), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n26) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[46]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[14]), .ZN(n86) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[47]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[15]), .ZN(n84) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[49]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[17]), .ZN(n82) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[45]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[13]), .ZN(n67) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[48]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[16]), .ZN(n83) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[43]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[11]), .ZN(n78) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[50]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[18]), .ZN(n81) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[42]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[10]), .ZN(n68) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[40]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[44]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[12]), .ZN(n79) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[41]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD2BWP30P140 U68 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[60]), .ZN(n17) );
  INVD2BWP30P140 U70 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[28]), .ZN(n92) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[61]), .ZN(n18) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[29]), .ZN(n89) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[62]), .ZN(n19) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[30]), .ZN(n88) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[63]), .ZN(n20) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[31]), .ZN(n87) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[59]), .ZN(n21) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[27]), .ZN(n70) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[52]), .ZN(n22) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[53]), .ZN(n23) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[21]), .ZN(n76) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[55]), .ZN(n24) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[23]), .ZN(n74) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[51]), .ZN(n25) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[19]), .ZN(n80) );
  OAI22D1BWP30P140 U88 ( .A1(n26), .A2(n25), .B1(n30), .B2(n80), .ZN(N306) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[57]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[25]), .ZN(n72) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[56]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[24]), .ZN(n73) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[58]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[26]), .ZN(n71) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[54]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[22]), .ZN(n75) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n57), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n58), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n59), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n60), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n61), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n62), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n63), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n85), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n85), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n85), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n85), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n85), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n85), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n85), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n85), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n85), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n85), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n85), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n85), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  INVD2BWP30P140 U140 ( .I(n69), .ZN(n91) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n85), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n85), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n85), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n85), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n85), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n85), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n85), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n85), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_67 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  OAI22D1BWP30P140 U5 ( .A1(n18), .A2(n6), .B1(n40), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U6 ( .A1(n18), .A2(n7), .B1(n40), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U7 ( .A1(n18), .A2(n8), .B1(n40), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U8 ( .A1(n18), .A2(n9), .B1(n40), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U9 ( .A1(n18), .A2(n10), .B1(n40), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n11), .B1(n40), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n12), .B1(n40), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n13), .B1(n40), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n14), .B1(n40), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n15), .B1(n40), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n16), .B1(n40), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U16 ( .A1(n32), .A2(n19), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U17 ( .A1(n32), .A2(n20), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U18 ( .A1(n32), .A2(n21), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U19 ( .A1(n32), .A2(n22), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U20 ( .A1(n32), .A2(n23), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n24), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n25), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n26), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n27), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n28), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n29), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n31), .B1(n30), .B2(n92), .ZN(N318) );
  ND2OPTIBD1BWP30P140 U28 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U29 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U30 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U31 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U32 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U33 ( .A1(n18), .A2(n17), .B1(n30), .B2(n77), .ZN(N306) );
  INVD1BWP30P140 U34 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U35 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U36 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U38 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U39 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U41 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U42 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U45 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U46 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U47 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U70 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n77) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n57), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n58), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n59), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n60), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n61), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n62), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n63), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_68 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n6), .B1(n40), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n7), .B1(n40), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n8), .B1(n40), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n9), .B1(n40), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n10), .B1(n40), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n11), .B1(n40), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n12), .B1(n40), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n13), .B1(n40), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n14), .B1(n40), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n15), .B1(n40), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n16), .B1(n40), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n19), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n20), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n21), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n22), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n23), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n24), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n25), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n26), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n27), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n28), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n29), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n31), .B1(n30), .B2(n92), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n77) );
  OAI22D1BWP30P140 U71 ( .A1(n18), .A2(n17), .B1(n30), .B2(n77), .ZN(N306) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n57), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n58), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n59), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n60), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n61), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n62), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n63), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_69 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n76), .ZN(n91) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n76) );
  OAI22D1BWP30P140 U5 ( .A1(n18), .A2(n17), .B1(n30), .B2(n89), .ZN(N306) );
  ND2OPTIBD1BWP30P140 U6 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U7 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U8 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U9 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U10 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n6), .B1(n40), .B2(n77), .ZN(N295) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n7), .B1(n40), .B2(n78), .ZN(N296) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n8), .B1(n40), .B2(n79), .ZN(N297) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n9), .B1(n40), .B2(n80), .ZN(N298) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n10), .B1(n40), .B2(n81), .ZN(N299) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n11), .B1(n40), .B2(n82), .ZN(N300) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n12), .B1(n40), .B2(n83), .ZN(N301) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n13), .B1(n40), .B2(n84), .ZN(N302) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n14), .B1(n40), .B2(n85), .ZN(N303) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n15), .B1(n40), .B2(n86), .ZN(N304) );
  OAI22D1BWP30P140 U21 ( .A1(n18), .A2(n16), .B1(n40), .B2(n87), .ZN(N305) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n19), .B1(n30), .B2(n92), .ZN(N307) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n20), .B1(n30), .B2(n75), .ZN(N308) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n21), .B1(n30), .B2(n74), .ZN(N309) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n22), .B1(n30), .B2(n65), .ZN(N310) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n23), .B1(n30), .B2(n66), .ZN(N311) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n24), .B1(n30), .B2(n67), .ZN(N312) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n25), .B1(n30), .B2(n68), .ZN(N313) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n26), .B1(n30), .B2(n69), .ZN(N314) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n27), .B1(n30), .B2(n70), .ZN(N315) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n28), .B1(n30), .B2(n71), .ZN(N316) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n29), .B1(n30), .B2(n72), .ZN(N317) );
  OAI22D1BWP30P140 U33 ( .A1(n32), .A2(n31), .B1(n30), .B2(n73), .ZN(N318) );
  INVD1BWP30P140 U34 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U35 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U36 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U38 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U39 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U41 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U42 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U45 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U46 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U47 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n77) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n78) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n79) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n80) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n81) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n82) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[14]), .ZN(n83) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[15]), .ZN(n84) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n85) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n86) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n87) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U70 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n89) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n92) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n75) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n65) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n66) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n67) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n68) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n70) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n71) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n72) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n73) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n64), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n63), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n62), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n61), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n60), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n59), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n58), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n57), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n91), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n91), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n91), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n91), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n91), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n91), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n91), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  INVD2BWP30P140 U147 ( .I(n76), .ZN(n88) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n88), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n88), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n88), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n88), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n88), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n88), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n88), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n88), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U156 ( .A1(n85), .A2(n88), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U157 ( .A1(n86), .A2(n88), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U158 ( .A1(n87), .A2(n88), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n88), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_70 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U6 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n6), .B1(n40), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n7), .B1(n40), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n8), .B1(n40), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n9), .B1(n40), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n10), .B1(n40), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n11), .B1(n40), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n12), .B1(n40), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n13), .B1(n40), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n14), .B1(n40), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n15), .B1(n40), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n16), .B1(n40), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n19), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n20), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n21), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n22), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n23), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n24), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n25), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U28 ( .A1(n32), .A2(n26), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U29 ( .A1(n32), .A2(n27), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U30 ( .A1(n32), .A2(n28), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U31 ( .A1(n32), .A2(n29), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U32 ( .A1(n32), .A2(n31), .B1(n30), .B2(n92), .ZN(N318) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U34 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n77) );
  OAI22D1BWP30P140 U71 ( .A1(n18), .A2(n17), .B1(n30), .B2(n77), .ZN(N306) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n40), .A2(n64), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n40), .A2(n63), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n40), .A2(n62), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n40), .A2(n61), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n46), .A2(n60), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n59), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n58), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n57), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_71 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n78), .ZN(n76) );
  INVD2BWP30P140 U4 ( .I(n56), .ZN(n78) );
  OAI22D1BWP30P140 U5 ( .A1(n18), .A2(n6), .B1(n41), .B2(n65), .ZN(N295) );
  OAI22D1BWP30P140 U6 ( .A1(n18), .A2(n7), .B1(n41), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U7 ( .A1(n18), .A2(n8), .B1(n41), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U8 ( .A1(n18), .A2(n9), .B1(n41), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U9 ( .A1(n18), .A2(n10), .B1(n41), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n11), .B1(n41), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n12), .B1(n41), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n13), .B1(n41), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n14), .B1(n41), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n15), .B1(n41), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n16), .B1(n41), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U16 ( .A1(n32), .A2(n19), .B1(n30), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U17 ( .A1(n32), .A2(n20), .B1(n30), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U18 ( .A1(n32), .A2(n21), .B1(n30), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U19 ( .A1(n32), .A2(n22), .B1(n30), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U20 ( .A1(n32), .A2(n23), .B1(n30), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U21 ( .A1(n32), .A2(n24), .B1(n30), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U22 ( .A1(n32), .A2(n25), .B1(n30), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U23 ( .A1(n32), .A2(n26), .B1(n30), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U24 ( .A1(n32), .A2(n27), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U25 ( .A1(n32), .A2(n28), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U26 ( .A1(n32), .A2(n29), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U27 ( .A1(n32), .A2(n31), .B1(n30), .B2(n92), .ZN(N318) );
  ND2OPTIBD1BWP30P140 U28 ( .A1(n55), .A2(n54), .ZN(n56) );
  MUX2ND0BWP30P140 U29 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  NR2D1BWP30P140 U30 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD1BWP30P140 U31 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U32 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U33 ( .A1(n18), .A2(n17), .B1(n30), .B2(n77), .ZN(N306) );
  INVD1BWP30P140 U34 ( .I(rst), .ZN(n1) );
  ND2D1BWP30P140 U35 ( .A1(n1), .A2(i_en), .ZN(n51) );
  NR2D1BWP30P140 U36 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n53) );
  INVD1BWP30P140 U38 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U39 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U41 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U42 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U45 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U46 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U47 ( .I(n33), .ZN(n41) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U70 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n77) );
  INVD2BWP30P140 U72 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U97 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U98 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[0]), .ZN(n63) );
  INVD2BWP30P140 U100 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[32]), .ZN(n36) );
  OAI22D1BWP30P140 U102 ( .A1(n46), .A2(n63), .B1(n45), .B2(n36), .ZN(N287) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[7]), .ZN(n62) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[39]), .ZN(n37) );
  OAI22D1BWP30P140 U105 ( .A1(n41), .A2(n62), .B1(n45), .B2(n37), .ZN(N294) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[6]), .ZN(n61) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[38]), .ZN(n38) );
  OAI22D1BWP30P140 U108 ( .A1(n41), .A2(n61), .B1(n45), .B2(n38), .ZN(N293) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[37]), .ZN(n39) );
  OAI22D1BWP30P140 U111 ( .A1(n41), .A2(n59), .B1(n45), .B2(n39), .ZN(N292) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[4]), .ZN(n57) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[36]), .ZN(n40) );
  OAI22D1BWP30P140 U114 ( .A1(n41), .A2(n57), .B1(n45), .B2(n40), .ZN(N291) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[3]), .ZN(n58) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[35]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n46), .A2(n58), .B1(n45), .B2(n42), .ZN(N290) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[34]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n46), .A2(n60), .B1(n45), .B2(n43), .ZN(N289) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[1]), .ZN(n64) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[33]), .ZN(n44) );
  OAI22D1BWP30P140 U123 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N288) );
  INVD1BWP30P140 U124 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U125 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U127 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n76), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n76), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n76), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n76), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n76), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n76), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n76), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n76), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_72 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  INVD2BWP30P140 U3 ( .I(n6), .ZN(n25) );
  ND2OPTIBD1BWP30P140 U4 ( .A1(n55), .A2(n54), .ZN(n56) );
  NR2D1BWP30P140 U5 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD2BWP30P140 U6 ( .I(n25), .ZN(n21) );
  INVD1BWP30P140 U7 ( .I(n56), .ZN(n78) );
  ND2D1BWP30P140 U8 ( .A1(n2), .A2(i_en), .ZN(n51) );
  INVD1BWP30P140 U9 ( .I(i_cmd[0]), .ZN(n22) );
  CKBD1BWP30P140 U10 ( .I(n56), .Z(n1) );
  INVD1BWP30P140 U11 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U12 ( .A1(n45), .A2(n7), .B1(n21), .B2(n77), .ZN(N306) );
  OAI22D1BWP30P140 U13 ( .A1(n20), .A2(n8), .B1(n21), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U14 ( .A1(n20), .A2(n9), .B1(n21), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U15 ( .A1(n20), .A2(n10), .B1(n21), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U16 ( .A1(n20), .A2(n11), .B1(n21), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U17 ( .A1(n20), .A2(n12), .B1(n21), .B2(n83), .ZN(N311) );
  OAI22D1BWP30P140 U18 ( .A1(n20), .A2(n13), .B1(n21), .B2(n84), .ZN(N312) );
  OAI22D1BWP30P140 U19 ( .A1(n20), .A2(n14), .B1(n21), .B2(n85), .ZN(N313) );
  OAI22D1BWP30P140 U20 ( .A1(n20), .A2(n15), .B1(n21), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U21 ( .A1(n20), .A2(n16), .B1(n21), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U22 ( .A1(n20), .A2(n17), .B1(n21), .B2(n92), .ZN(N316) );
  OAI22D1BWP30P140 U23 ( .A1(n20), .A2(n18), .B1(n21), .B2(n88), .ZN(N317) );
  OAI22D1BWP30P140 U24 ( .A1(n20), .A2(n19), .B1(n21), .B2(n89), .ZN(N318) );
  INVD1BWP30P140 U25 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U26 ( .A1(n51), .A2(n22), .ZN(n4) );
  INVD1BWP30P140 U27 ( .I(i_valid[0]), .ZN(n53) );
  INVD2BWP30P140 U28 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U29 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U30 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U31 ( .I(n5), .ZN(n23) );
  INVD3BWP30P140 U32 ( .I(n23), .ZN(n45) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[51]), .ZN(n7) );
  INR2D1BWP30P140 U34 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U35 ( .A1(n47), .A2(n22), .ZN(n6) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[19]), .ZN(n77) );
  INVD2BWP30P140 U37 ( .I(n23), .ZN(n20) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[52]), .ZN(n8) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[53]), .ZN(n9) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[54]), .ZN(n10) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[55]), .ZN(n11) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[56]), .ZN(n12) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[24]), .ZN(n83) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[57]), .ZN(n13) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[25]), .ZN(n84) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[58]), .ZN(n14) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[26]), .ZN(n85) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[59]), .ZN(n15) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[60]), .ZN(n16) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[61]), .ZN(n17) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[29]), .ZN(n92) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[62]), .ZN(n18) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[30]), .ZN(n88) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[63]), .ZN(n19) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[31]), .ZN(n89) );
  OAI31D1BWP30P140 U62 ( .A1(n51), .A2(n52), .A3(n22), .B(n21), .ZN(N353) );
  INVD2BWP30P140 U63 ( .I(n25), .ZN(n46) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD2BWP30P140 U65 ( .I(n23), .ZN(n38) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[36]), .ZN(n24) );
  OAI22D1BWP30P140 U67 ( .A1(n46), .A2(n62), .B1(n38), .B2(n24), .ZN(N291) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[3]), .ZN(n64) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[35]), .ZN(n26) );
  OAI22D1BWP30P140 U70 ( .A1(n46), .A2(n64), .B1(n38), .B2(n26), .ZN(N290) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[2]), .ZN(n58) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[34]), .ZN(n27) );
  OAI22D1BWP30P140 U73 ( .A1(n46), .A2(n58), .B1(n38), .B2(n27), .ZN(N289) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[1]), .ZN(n61) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[33]), .ZN(n28) );
  OAI22D1BWP30P140 U76 ( .A1(n46), .A2(n61), .B1(n38), .B2(n28), .ZN(N288) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[0]), .ZN(n59) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[32]), .ZN(n29) );
  OAI22D1BWP30P140 U79 ( .A1(n46), .A2(n59), .B1(n38), .B2(n29), .ZN(N287) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[7]), .ZN(n60) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[39]), .ZN(n30) );
  OAI22D1BWP30P140 U82 ( .A1(n46), .A2(n60), .B1(n38), .B2(n30), .ZN(N294) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[6]), .ZN(n57) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[38]), .ZN(n31) );
  OAI22D1BWP30P140 U85 ( .A1(n46), .A2(n57), .B1(n38), .B2(n31), .ZN(N293) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[5]), .ZN(n63) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[37]), .ZN(n32) );
  OAI22D1BWP30P140 U88 ( .A1(n46), .A2(n63), .B1(n45), .B2(n32), .ZN(N292) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[40]), .ZN(n33) );
  OAI22D1BWP30P140 U91 ( .A1(n46), .A2(n65), .B1(n45), .B2(n33), .ZN(N295) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[41]), .ZN(n34) );
  OAI22D1BWP30P140 U94 ( .A1(n46), .A2(n66), .B1(n45), .B2(n34), .ZN(N296) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[42]), .ZN(n35) );
  OAI22D1BWP30P140 U97 ( .A1(n46), .A2(n67), .B1(n45), .B2(n35), .ZN(N297) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[43]), .ZN(n36) );
  OAI22D1BWP30P140 U100 ( .A1(n46), .A2(n68), .B1(n45), .B2(n36), .ZN(N298) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[44]), .ZN(n37) );
  OAI22D1BWP30P140 U103 ( .A1(n46), .A2(n69), .B1(n38), .B2(n37), .ZN(N299) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[45]), .ZN(n39) );
  OAI22D1BWP30P140 U106 ( .A1(n46), .A2(n70), .B1(n45), .B2(n39), .ZN(N300) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[46]), .ZN(n40) );
  OAI22D1BWP30P140 U109 ( .A1(n46), .A2(n71), .B1(n45), .B2(n40), .ZN(N301) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[47]), .ZN(n41) );
  OAI22D1BWP30P140 U112 ( .A1(n46), .A2(n72), .B1(n45), .B2(n41), .ZN(N302) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[48]), .ZN(n42) );
  OAI22D1BWP30P140 U115 ( .A1(n46), .A2(n73), .B1(n45), .B2(n42), .ZN(N303) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[49]), .ZN(n43) );
  OAI22D1BWP30P140 U118 ( .A1(n46), .A2(n74), .B1(n45), .B2(n43), .ZN(N304) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[50]), .ZN(n44) );
  OAI22D1BWP30P140 U121 ( .A1(n46), .A2(n75), .B1(n45), .B2(n44), .ZN(N305) );
  INVD1BWP30P140 U122 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U123 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U125 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MUX2NUD1BWP30P140 U126 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  MOAI22D1BWP30P140 U127 ( .A1(n57), .A2(n1), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n1), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n1), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n1), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n1), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n1), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n1), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n1), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  INVD2BWP30P140 U135 ( .I(n78), .ZN(n76) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_73 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  INVD2BWP30P140 U3 ( .I(n6), .ZN(n26) );
  INVD2BWP30P140 U4 ( .I(n26), .ZN(n21) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n55), .A2(n54), .ZN(n56) );
  NR2D1BWP30P140 U6 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  OAI22D1BWP30P140 U7 ( .A1(n20), .A2(n8), .B1(n21), .B2(n85), .ZN(N307) );
  OAI22D1BWP30P140 U8 ( .A1(n20), .A2(n9), .B1(n21), .B2(n86), .ZN(N308) );
  OAI22D1BWP30P140 U9 ( .A1(n20), .A2(n10), .B1(n21), .B2(n87), .ZN(N309) );
  OAI22D1BWP30P140 U10 ( .A1(n20), .A2(n11), .B1(n21), .B2(n88), .ZN(N310) );
  OAI22D1BWP30P140 U11 ( .A1(n20), .A2(n12), .B1(n21), .B2(n89), .ZN(N311) );
  OAI22D1BWP30P140 U12 ( .A1(n20), .A2(n13), .B1(n21), .B2(n92), .ZN(N312) );
  OAI22D1BWP30P140 U13 ( .A1(n20), .A2(n14), .B1(n21), .B2(n65), .ZN(N313) );
  OAI22D1BWP30P140 U14 ( .A1(n20), .A2(n15), .B1(n21), .B2(n66), .ZN(N314) );
  OAI22D1BWP30P140 U15 ( .A1(n20), .A2(n16), .B1(n21), .B2(n67), .ZN(N315) );
  OAI22D1BWP30P140 U16 ( .A1(n20), .A2(n17), .B1(n21), .B2(n68), .ZN(N316) );
  OAI22D1BWP30P140 U17 ( .A1(n20), .A2(n18), .B1(n21), .B2(n69), .ZN(N317) );
  OAI22D1BWP30P140 U18 ( .A1(n20), .A2(n19), .B1(n21), .B2(n70), .ZN(N318) );
  INVD1BWP30P140 U19 ( .I(n56), .ZN(n71) );
  ND2D1BWP30P140 U20 ( .A1(n2), .A2(i_en), .ZN(n51) );
  INVD1BWP30P140 U21 ( .I(i_cmd[0]), .ZN(n22) );
  CKBD1BWP30P140 U22 ( .I(n56), .Z(n1) );
  INVD1BWP30P140 U23 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U24 ( .A1(n45), .A2(n7), .B1(n21), .B2(n84), .ZN(N306) );
  INVD1BWP30P140 U25 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U26 ( .A1(n51), .A2(n22), .ZN(n4) );
  INVD1BWP30P140 U27 ( .I(i_valid[0]), .ZN(n53) );
  INVD2BWP30P140 U28 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U29 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U30 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U31 ( .I(n5), .ZN(n23) );
  INVD3BWP30P140 U32 ( .I(n23), .ZN(n45) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[51]), .ZN(n7) );
  INR2D1BWP30P140 U34 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U35 ( .A1(n47), .A2(n22), .ZN(n6) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[19]), .ZN(n84) );
  INVD2BWP30P140 U37 ( .I(n23), .ZN(n20) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[52]), .ZN(n8) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[20]), .ZN(n85) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[53]), .ZN(n9) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[21]), .ZN(n86) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[54]), .ZN(n10) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[22]), .ZN(n87) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[55]), .ZN(n11) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[23]), .ZN(n88) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[56]), .ZN(n12) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[24]), .ZN(n89) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[57]), .ZN(n13) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[25]), .ZN(n92) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[58]), .ZN(n14) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[26]), .ZN(n65) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[59]), .ZN(n15) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[27]), .ZN(n66) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[60]), .ZN(n16) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[28]), .ZN(n67) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[61]), .ZN(n17) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[29]), .ZN(n68) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[62]), .ZN(n18) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[30]), .ZN(n69) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[63]), .ZN(n19) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[31]), .ZN(n70) );
  OAI31D1BWP30P140 U62 ( .A1(n51), .A2(n52), .A3(n22), .B(n21), .ZN(N353) );
  INVD2BWP30P140 U63 ( .I(n26), .ZN(n46) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD2BWP30P140 U65 ( .I(n23), .ZN(n38) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[39]), .ZN(n24) );
  OAI22D1BWP30P140 U67 ( .A1(n46), .A2(n57), .B1(n38), .B2(n24), .ZN(N294) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[38]), .ZN(n25) );
  OAI22D1BWP30P140 U70 ( .A1(n46), .A2(n58), .B1(n38), .B2(n25), .ZN(N293) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[35]), .ZN(n27) );
  OAI22D1BWP30P140 U73 ( .A1(n46), .A2(n61), .B1(n38), .B2(n27), .ZN(N290) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[34]), .ZN(n28) );
  OAI22D1BWP30P140 U76 ( .A1(n46), .A2(n62), .B1(n38), .B2(n28), .ZN(N289) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[33]), .ZN(n29) );
  OAI22D1BWP30P140 U79 ( .A1(n46), .A2(n63), .B1(n38), .B2(n29), .ZN(N288) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[37]), .ZN(n30) );
  OAI22D1BWP30P140 U82 ( .A1(n46), .A2(n59), .B1(n38), .B2(n30), .ZN(N292) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[36]), .ZN(n31) );
  OAI22D1BWP30P140 U85 ( .A1(n46), .A2(n60), .B1(n38), .B2(n31), .ZN(N291) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[32]), .ZN(n32) );
  OAI22D1BWP30P140 U88 ( .A1(n46), .A2(n64), .B1(n45), .B2(n32), .ZN(N287) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[9]), .ZN(n73) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[41]), .ZN(n33) );
  OAI22D1BWP30P140 U91 ( .A1(n46), .A2(n73), .B1(n45), .B2(n33), .ZN(N296) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[11]), .ZN(n75) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[43]), .ZN(n34) );
  OAI22D1BWP30P140 U94 ( .A1(n46), .A2(n75), .B1(n45), .B2(n34), .ZN(N298) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[12]), .ZN(n76) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[44]), .ZN(n35) );
  OAI22D1BWP30P140 U97 ( .A1(n46), .A2(n76), .B1(n45), .B2(n35), .ZN(N299) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[13]), .ZN(n77) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[45]), .ZN(n36) );
  OAI22D1BWP30P140 U100 ( .A1(n46), .A2(n77), .B1(n45), .B2(n36), .ZN(N300) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[14]), .ZN(n78) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[46]), .ZN(n37) );
  OAI22D1BWP30P140 U103 ( .A1(n46), .A2(n78), .B1(n38), .B2(n37), .ZN(N301) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[15]), .ZN(n79) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[47]), .ZN(n39) );
  OAI22D1BWP30P140 U106 ( .A1(n46), .A2(n79), .B1(n45), .B2(n39), .ZN(N302) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[16]), .ZN(n80) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[48]), .ZN(n40) );
  OAI22D1BWP30P140 U109 ( .A1(n46), .A2(n80), .B1(n45), .B2(n40), .ZN(N303) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[17]), .ZN(n81) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[49]), .ZN(n41) );
  OAI22D1BWP30P140 U112 ( .A1(n46), .A2(n81), .B1(n45), .B2(n41), .ZN(N304) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[18]), .ZN(n82) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[50]), .ZN(n42) );
  OAI22D1BWP30P140 U115 ( .A1(n46), .A2(n82), .B1(n45), .B2(n42), .ZN(N305) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[8]), .ZN(n72) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[40]), .ZN(n43) );
  OAI22D1BWP30P140 U118 ( .A1(n46), .A2(n72), .B1(n45), .B2(n43), .ZN(N295) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[10]), .ZN(n74) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[42]), .ZN(n44) );
  OAI22D1BWP30P140 U121 ( .A1(n46), .A2(n74), .B1(n45), .B2(n44), .ZN(N297) );
  INVD1BWP30P140 U122 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U123 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U125 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MUX2NUD1BWP30P140 U126 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  MOAI22D1BWP30P140 U127 ( .A1(n57), .A2(n1), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n1), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n1), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n1), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n1), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n1), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n1), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n1), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  INVD2BWP30P140 U135 ( .I(n71), .ZN(n91) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  INVD2BWP30P140 U142 ( .I(n71), .ZN(n83) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n83), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n83), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n83), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n83), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n83), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n83), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n83), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n83), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n83), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n83), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n83), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n83), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_74 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  INVD2BWP30P140 U3 ( .I(n6), .ZN(n28) );
  ND2OPTIBD1BWP30P140 U4 ( .A1(n55), .A2(n54), .ZN(n56) );
  NR2D1BWP30P140 U5 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  INVD2BWP30P140 U6 ( .I(n28), .ZN(n21) );
  INVD1BWP30P140 U7 ( .I(n56), .ZN(n67) );
  ND2D1BWP30P140 U8 ( .A1(n2), .A2(i_en), .ZN(n51) );
  INVD1BWP30P140 U9 ( .I(i_cmd[0]), .ZN(n22) );
  CKBD1BWP30P140 U10 ( .I(n56), .Z(n1) );
  INVD1BWP30P140 U11 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U12 ( .A1(n45), .A2(n20), .B1(n21), .B2(n77), .ZN(N306) );
  OAI22D1BWP30P140 U13 ( .A1(n19), .A2(n18), .B1(n21), .B2(n76), .ZN(N307) );
  OAI22D1BWP30P140 U14 ( .A1(n19), .A2(n17), .B1(n21), .B2(n75), .ZN(N308) );
  OAI22D1BWP30P140 U15 ( .A1(n19), .A2(n16), .B1(n21), .B2(n74), .ZN(N309) );
  OAI22D1BWP30P140 U16 ( .A1(n19), .A2(n15), .B1(n21), .B2(n73), .ZN(N310) );
  OAI22D1BWP30P140 U17 ( .A1(n19), .A2(n14), .B1(n21), .B2(n72), .ZN(N311) );
  OAI22D1BWP30P140 U18 ( .A1(n19), .A2(n13), .B1(n21), .B2(n71), .ZN(N312) );
  OAI22D1BWP30P140 U19 ( .A1(n19), .A2(n12), .B1(n21), .B2(n70), .ZN(N313) );
  OAI22D1BWP30P140 U20 ( .A1(n19), .A2(n11), .B1(n21), .B2(n69), .ZN(N314) );
  OAI22D1BWP30P140 U21 ( .A1(n19), .A2(n10), .B1(n21), .B2(n68), .ZN(N315) );
  OAI22D1BWP30P140 U22 ( .A1(n19), .A2(n9), .B1(n21), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U23 ( .A1(n19), .A2(n8), .B1(n21), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U24 ( .A1(n19), .A2(n7), .B1(n21), .B2(n92), .ZN(N318) );
  INVD1BWP30P140 U25 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U26 ( .A1(n51), .A2(n22), .ZN(n4) );
  INVD1BWP30P140 U27 ( .I(i_valid[0]), .ZN(n53) );
  INVD2BWP30P140 U28 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U29 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U30 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U31 ( .I(n5), .ZN(n23) );
  INVD2BWP30P140 U32 ( .I(n23), .ZN(n19) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[63]), .ZN(n7) );
  INR2D1BWP30P140 U34 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U35 ( .A1(n47), .A2(n22), .ZN(n6) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[62]), .ZN(n8) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[61]), .ZN(n9) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[60]), .ZN(n10) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[28]), .ZN(n68) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[59]), .ZN(n11) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[58]), .ZN(n12) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[26]), .ZN(n70) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[57]), .ZN(n13) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[25]), .ZN(n71) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[56]), .ZN(n14) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[24]), .ZN(n72) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[55]), .ZN(n15) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[23]), .ZN(n73) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[54]), .ZN(n16) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[53]), .ZN(n17) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[21]), .ZN(n75) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[52]), .ZN(n18) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[20]), .ZN(n76) );
  INVD3BWP30P140 U59 ( .I(n23), .ZN(n45) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[51]), .ZN(n20) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[19]), .ZN(n77) );
  OAI31D1BWP30P140 U62 ( .A1(n51), .A2(n52), .A3(n22), .B(n21), .ZN(N353) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD2BWP30P140 U64 ( .I(n23), .ZN(n38) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[35]), .ZN(n24) );
  OAI22D1BWP30P140 U66 ( .A1(n46), .A2(n61), .B1(n38), .B2(n24), .ZN(N290) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[32]), .ZN(n25) );
  OAI22D1BWP30P140 U69 ( .A1(n46), .A2(n64), .B1(n38), .B2(n25), .ZN(N287) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[33]), .ZN(n26) );
  OAI22D1BWP30P140 U72 ( .A1(n46), .A2(n63), .B1(n38), .B2(n26), .ZN(N288) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[34]), .ZN(n27) );
  OAI22D1BWP30P140 U75 ( .A1(n46), .A2(n62), .B1(n38), .B2(n27), .ZN(N289) );
  INVD2BWP30P140 U76 ( .I(n28), .ZN(n46) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[36]), .ZN(n29) );
  OAI22D1BWP30P140 U79 ( .A1(n46), .A2(n60), .B1(n38), .B2(n29), .ZN(N291) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[37]), .ZN(n30) );
  OAI22D1BWP30P140 U82 ( .A1(n46), .A2(n59), .B1(n38), .B2(n30), .ZN(N292) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[38]), .ZN(n31) );
  OAI22D1BWP30P140 U85 ( .A1(n46), .A2(n58), .B1(n38), .B2(n31), .ZN(N293) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[39]), .ZN(n32) );
  OAI22D1BWP30P140 U88 ( .A1(n46), .A2(n57), .B1(n45), .B2(n32), .ZN(N294) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[18]), .ZN(n78) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[50]), .ZN(n33) );
  OAI22D1BWP30P140 U91 ( .A1(n46), .A2(n78), .B1(n45), .B2(n33), .ZN(N305) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[17]), .ZN(n79) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[49]), .ZN(n34) );
  OAI22D1BWP30P140 U94 ( .A1(n46), .A2(n79), .B1(n45), .B2(n34), .ZN(N304) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[16]), .ZN(n80) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[48]), .ZN(n35) );
  OAI22D1BWP30P140 U97 ( .A1(n46), .A2(n80), .B1(n45), .B2(n35), .ZN(N303) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[15]), .ZN(n81) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[47]), .ZN(n36) );
  OAI22D1BWP30P140 U100 ( .A1(n46), .A2(n81), .B1(n45), .B2(n36), .ZN(N302) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[14]), .ZN(n82) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[46]), .ZN(n37) );
  OAI22D1BWP30P140 U103 ( .A1(n46), .A2(n82), .B1(n38), .B2(n37), .ZN(N301) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[13]), .ZN(n83) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[45]), .ZN(n39) );
  OAI22D1BWP30P140 U106 ( .A1(n46), .A2(n83), .B1(n45), .B2(n39), .ZN(N300) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[12]), .ZN(n84) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[44]), .ZN(n40) );
  OAI22D1BWP30P140 U109 ( .A1(n46), .A2(n84), .B1(n45), .B2(n40), .ZN(N299) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[11]), .ZN(n85) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[43]), .ZN(n41) );
  OAI22D1BWP30P140 U112 ( .A1(n46), .A2(n85), .B1(n45), .B2(n41), .ZN(N298) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[10]), .ZN(n87) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[42]), .ZN(n42) );
  OAI22D1BWP30P140 U115 ( .A1(n46), .A2(n87), .B1(n45), .B2(n42), .ZN(N297) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[9]), .ZN(n65) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[41]), .ZN(n43) );
  OAI22D1BWP30P140 U118 ( .A1(n46), .A2(n65), .B1(n45), .B2(n43), .ZN(N296) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[40]), .ZN(n44) );
  OAI22D1BWP30P140 U121 ( .A1(n46), .A2(n66), .B1(n45), .B2(n44), .ZN(N295) );
  INVD1BWP30P140 U122 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U123 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U125 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MUX2NUD1BWP30P140 U126 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  MOAI22D1BWP30P140 U127 ( .A1(n57), .A2(n1), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n1), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n1), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n1), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n1), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n1), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n1), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n1), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  INVD2BWP30P140 U135 ( .I(n67), .ZN(n86) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n86), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n86), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  INVD2BWP30P140 U138 ( .I(n67), .ZN(n91) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n86), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n86), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n86), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n86), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n86), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n86), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n86), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n86), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U156 ( .A1(n85), .A2(n86), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n86), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_75 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n45), .A2(n19), .B1(n20), .B2(n80), .ZN(N306) );
  INVD3BWP30P140 U4 ( .I(n28), .ZN(n20) );
  INVD1BWP30P140 U5 ( .I(n5), .ZN(n28) );
  ND2OPTIBD1BWP30P140 U6 ( .A1(n47), .A2(n21), .ZN(n5) );
  OAI22D1BWP30P140 U7 ( .A1(n18), .A2(n17), .B1(n20), .B2(n78), .ZN(N307) );
  OAI22D1BWP30P140 U8 ( .A1(n18), .A2(n16), .B1(n20), .B2(n76), .ZN(N308) );
  OAI22D1BWP30P140 U9 ( .A1(n18), .A2(n15), .B1(n20), .B2(n75), .ZN(N309) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n14), .B1(n20), .B2(n74), .ZN(N310) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n13), .B1(n20), .B2(n73), .ZN(N311) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n12), .B1(n20), .B2(n72), .ZN(N312) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n11), .B1(n20), .B2(n71), .ZN(N313) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n10), .B1(n20), .B2(n70), .ZN(N314) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n9), .B1(n20), .B2(n69), .ZN(N315) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n8), .B1(n20), .B2(n68), .ZN(N316) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n7), .B1(n20), .B2(n67), .ZN(N317) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n6), .B1(n20), .B2(n66), .ZN(N318) );
  ND2D1BWP30P140 U19 ( .A1(n1), .A2(i_en), .ZN(n51) );
  INVD1BWP30P140 U20 ( .I(n91), .ZN(n49) );
  INVD1BWP30P140 U21 ( .I(rst), .ZN(n1) );
  INVD1P5BWP30P140 U22 ( .I(i_cmd[0]), .ZN(n21) );
  NR2D1BWP30P140 U23 ( .A1(n51), .A2(n21), .ZN(n3) );
  INVD1BWP30P140 U24 ( .I(i_valid[0]), .ZN(n53) );
  INVD2BWP30P140 U25 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U26 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U27 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U28 ( .I(n4), .ZN(n22) );
  INVD2BWP30P140 U29 ( .I(n22), .ZN(n18) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[63]), .ZN(n6) );
  INR2D1BWP30P140 U31 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[31]), .ZN(n66) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[62]), .ZN(n7) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[30]), .ZN(n67) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[61]), .ZN(n8) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[29]), .ZN(n68) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[60]), .ZN(n9) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[28]), .ZN(n69) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[59]), .ZN(n10) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[27]), .ZN(n70) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[58]), .ZN(n11) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[26]), .ZN(n71) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[57]), .ZN(n12) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[25]), .ZN(n72) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[56]), .ZN(n13) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[24]), .ZN(n73) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[55]), .ZN(n14) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[23]), .ZN(n74) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[54]), .ZN(n15) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[22]), .ZN(n75) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[53]), .ZN(n16) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[21]), .ZN(n76) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[52]), .ZN(n17) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[20]), .ZN(n78) );
  INVD3BWP30P140 U55 ( .I(n22), .ZN(n45) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[51]), .ZN(n19) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[19]), .ZN(n80) );
  OAI31D1BWP30P140 U58 ( .A1(n51), .A2(n52), .A3(n21), .B(n20), .ZN(N353) );
  INVD1BWP30P140 U59 ( .I(n28), .ZN(n27) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD2BWP30P140 U61 ( .I(n22), .ZN(n38) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[32]), .ZN(n23) );
  OAI22D1BWP30P140 U63 ( .A1(n27), .A2(n57), .B1(n38), .B2(n23), .ZN(N287) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[33]), .ZN(n24) );
  OAI22D1BWP30P140 U66 ( .A1(n27), .A2(n58), .B1(n38), .B2(n24), .ZN(N288) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[34]), .ZN(n25) );
  OAI22D1BWP30P140 U69 ( .A1(n27), .A2(n59), .B1(n38), .B2(n25), .ZN(N289) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[35]), .ZN(n26) );
  OAI22D1BWP30P140 U72 ( .A1(n27), .A2(n60), .B1(n38), .B2(n26), .ZN(N290) );
  INVD2BWP30P140 U73 ( .I(n28), .ZN(n46) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[36]), .ZN(n29) );
  OAI22D1BWP30P140 U76 ( .A1(n46), .A2(n62), .B1(n38), .B2(n29), .ZN(N291) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[5]), .ZN(n61) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[37]), .ZN(n30) );
  OAI22D1BWP30P140 U79 ( .A1(n46), .A2(n61), .B1(n38), .B2(n30), .ZN(N292) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[38]), .ZN(n31) );
  OAI22D1BWP30P140 U82 ( .A1(n46), .A2(n63), .B1(n38), .B2(n31), .ZN(N293) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[7]), .ZN(n65) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[39]), .ZN(n32) );
  OAI22D1BWP30P140 U85 ( .A1(n46), .A2(n65), .B1(n45), .B2(n32), .ZN(N294) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[18]), .ZN(n81) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[50]), .ZN(n33) );
  OAI22D1BWP30P140 U88 ( .A1(n46), .A2(n81), .B1(n45), .B2(n33), .ZN(N305) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[17]), .ZN(n82) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[49]), .ZN(n34) );
  OAI22D1BWP30P140 U91 ( .A1(n46), .A2(n82), .B1(n45), .B2(n34), .ZN(N304) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[16]), .ZN(n83) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[48]), .ZN(n35) );
  OAI22D1BWP30P140 U94 ( .A1(n46), .A2(n83), .B1(n45), .B2(n35), .ZN(N303) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[15]), .ZN(n84) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[47]), .ZN(n36) );
  OAI22D1BWP30P140 U97 ( .A1(n46), .A2(n84), .B1(n45), .B2(n36), .ZN(N302) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[14]), .ZN(n85) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[46]), .ZN(n37) );
  OAI22D1BWP30P140 U100 ( .A1(n46), .A2(n85), .B1(n38), .B2(n37), .ZN(N301) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[13]), .ZN(n86) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[45]), .ZN(n39) );
  OAI22D1BWP30P140 U103 ( .A1(n46), .A2(n86), .B1(n45), .B2(n39), .ZN(N300) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[12]), .ZN(n87) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[44]), .ZN(n40) );
  OAI22D1BWP30P140 U106 ( .A1(n46), .A2(n87), .B1(n45), .B2(n40), .ZN(N299) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[11]), .ZN(n88) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[43]), .ZN(n41) );
  OAI22D1BWP30P140 U109 ( .A1(n46), .A2(n88), .B1(n45), .B2(n41), .ZN(N298) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[10]), .ZN(n89) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[42]), .ZN(n42) );
  OAI22D1BWP30P140 U112 ( .A1(n46), .A2(n89), .B1(n45), .B2(n42), .ZN(N297) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[9]), .ZN(n90) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[41]), .ZN(n43) );
  OAI22D1BWP30P140 U115 ( .A1(n46), .A2(n90), .B1(n45), .B2(n43), .ZN(N296) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[8]), .ZN(n93) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[40]), .ZN(n44) );
  OAI22D1BWP30P140 U118 ( .A1(n46), .A2(n93), .B1(n45), .B2(n44), .ZN(N295) );
  INVD1BWP30P140 U119 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U120 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U121 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n91) );
  OAI21D1BWP30P140 U122 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  NR2D1BWP30P140 U123 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  MUX2NUD1BWP30P140 U124 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n55), .A2(n54), .ZN(n56) );
  INVD2BWP30P140 U126 ( .I(n56), .ZN(n79) );
  INVD1BWP30P140 U127 ( .I(n79), .ZN(n64) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n64), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n64), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n64), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n64), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n64), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n64), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n64), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n64), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  INVD2BWP30P140 U136 ( .I(n79), .ZN(n77) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n77), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n77), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n77), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n77), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n77), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n77), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n77), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n77), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n77), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n77), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n77), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n77), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  INVD2BWP30P140 U149 ( .I(n79), .ZN(n92) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n92), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_76 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  INVD2BWP30P140 U3 ( .I(n27), .ZN(n20) );
  INVD2BWP30P140 U4 ( .I(i_cmd[0]), .ZN(n21) );
  CKAN2D1BWP30P140 U5 ( .A1(i_valid[0]), .A2(n47), .Z(n46) );
  INVD1BWP30P140 U6 ( .I(n5), .ZN(n27) );
  ND2OPTIBD1BWP30P140 U7 ( .A1(n46), .A2(n21), .ZN(n5) );
  ND2D1BWP30P140 U8 ( .A1(n1), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n48) );
  OAI22D1BWP30P140 U10 ( .A1(n44), .A2(n19), .B1(n20), .B2(n79), .ZN(N306) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n17), .B1(n20), .B2(n77), .ZN(N307) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n16), .B1(n20), .B2(n75), .ZN(N308) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n15), .B1(n20), .B2(n74), .ZN(N309) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n14), .B1(n20), .B2(n73), .ZN(N310) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n13), .B1(n20), .B2(n72), .ZN(N311) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n12), .B1(n20), .B2(n71), .ZN(N312) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n11), .B1(n20), .B2(n70), .ZN(N313) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n10), .B1(n20), .B2(n69), .ZN(N314) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n9), .B1(n20), .B2(n68), .ZN(N315) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n8), .B1(n20), .B2(n67), .ZN(N316) );
  OAI22D1BWP30P140 U21 ( .A1(n18), .A2(n7), .B1(n20), .B2(n66), .ZN(N317) );
  OAI22D1BWP30P140 U22 ( .A1(n18), .A2(n6), .B1(n20), .B2(n65), .ZN(N318) );
  INVD1BWP30P140 U23 ( .I(rst), .ZN(n1) );
  NR2D1BWP30P140 U24 ( .A1(n50), .A2(n21), .ZN(n3) );
  INVD1BWP30P140 U25 ( .I(i_valid[0]), .ZN(n52) );
  INVD2BWP30P140 U26 ( .I(i_valid[1]), .ZN(n51) );
  MUX2NUD1BWP30P140 U27 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U28 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U29 ( .I(n4), .ZN(n22) );
  INVD2BWP30P140 U30 ( .I(n22), .ZN(n18) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[63]), .ZN(n6) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[31]), .ZN(n65) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[62]), .ZN(n7) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[30]), .ZN(n66) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[61]), .ZN(n8) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[29]), .ZN(n67) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[60]), .ZN(n9) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[28]), .ZN(n68) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[59]), .ZN(n10) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[58]), .ZN(n11) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[26]), .ZN(n70) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[57]), .ZN(n12) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[25]), .ZN(n71) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[56]), .ZN(n13) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[24]), .ZN(n72) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[55]), .ZN(n14) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[23]), .ZN(n73) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[54]), .ZN(n15) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[53]), .ZN(n16) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[21]), .ZN(n75) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[52]), .ZN(n17) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD3BWP30P140 U55 ( .I(n22), .ZN(n44) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[51]), .ZN(n19) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[19]), .ZN(n79) );
  OAI31D1BWP30P140 U58 ( .A1(n50), .A2(n51), .A3(n21), .B(n20), .ZN(N353) );
  INVD2BWP30P140 U59 ( .I(n27), .ZN(n45) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD2BWP30P140 U61 ( .I(n22), .ZN(n37) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[36]), .ZN(n23) );
  OAI22D1BWP30P140 U63 ( .A1(n45), .A2(n60), .B1(n37), .B2(n23), .ZN(N291) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[5]), .ZN(n61) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[37]), .ZN(n24) );
  OAI22D1BWP30P140 U66 ( .A1(n45), .A2(n61), .B1(n37), .B2(n24), .ZN(N292) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[6]), .ZN(n62) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[38]), .ZN(n25) );
  OAI22D1BWP30P140 U69 ( .A1(n45), .A2(n62), .B1(n37), .B2(n25), .ZN(N293) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[39]), .ZN(n26) );
  OAI22D1BWP30P140 U72 ( .A1(n45), .A2(n64), .B1(n37), .B2(n26), .ZN(N294) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[3]), .ZN(n59) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[35]), .ZN(n28) );
  OAI22D1BWP30P140 U75 ( .A1(n45), .A2(n59), .B1(n37), .B2(n28), .ZN(N290) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[2]), .ZN(n58) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[34]), .ZN(n29) );
  OAI22D1BWP30P140 U78 ( .A1(n20), .A2(n58), .B1(n37), .B2(n29), .ZN(N289) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[1]), .ZN(n57) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[33]), .ZN(n30) );
  OAI22D1BWP30P140 U81 ( .A1(n45), .A2(n57), .B1(n37), .B2(n30), .ZN(N288) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[0]), .ZN(n56) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[32]), .ZN(n31) );
  OAI22D1BWP30P140 U84 ( .A1(n20), .A2(n56), .B1(n44), .B2(n31), .ZN(N287) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[18]), .ZN(n80) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[50]), .ZN(n32) );
  OAI22D1BWP30P140 U87 ( .A1(n45), .A2(n80), .B1(n44), .B2(n32), .ZN(N305) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[17]), .ZN(n81) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[49]), .ZN(n33) );
  OAI22D1BWP30P140 U90 ( .A1(n45), .A2(n81), .B1(n44), .B2(n33), .ZN(N304) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[16]), .ZN(n82) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[48]), .ZN(n34) );
  OAI22D1BWP30P140 U93 ( .A1(n45), .A2(n82), .B1(n44), .B2(n34), .ZN(N303) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[15]), .ZN(n83) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[47]), .ZN(n35) );
  OAI22D1BWP30P140 U96 ( .A1(n45), .A2(n83), .B1(n44), .B2(n35), .ZN(N302) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[14]), .ZN(n84) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[46]), .ZN(n36) );
  OAI22D1BWP30P140 U99 ( .A1(n45), .A2(n84), .B1(n37), .B2(n36), .ZN(N301) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[13]), .ZN(n85) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[45]), .ZN(n38) );
  OAI22D1BWP30P140 U102 ( .A1(n45), .A2(n85), .B1(n44), .B2(n38), .ZN(N300) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[44]), .ZN(n39) );
  OAI22D1BWP30P140 U105 ( .A1(n45), .A2(n86), .B1(n44), .B2(n39), .ZN(N299) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[11]), .ZN(n87) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[43]), .ZN(n40) );
  OAI22D1BWP30P140 U108 ( .A1(n45), .A2(n87), .B1(n44), .B2(n40), .ZN(N298) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[42]), .ZN(n41) );
  OAI22D1BWP30P140 U111 ( .A1(n45), .A2(n88), .B1(n44), .B2(n41), .ZN(N297) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[9]), .ZN(n89) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[41]), .ZN(n42) );
  OAI22D1BWP30P140 U114 ( .A1(n45), .A2(n89), .B1(n44), .B2(n42), .ZN(N296) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[8]), .ZN(n92) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[40]), .ZN(n43) );
  OAI22D1BWP30P140 U117 ( .A1(n45), .A2(n92), .B1(n44), .B2(n43), .ZN(N295) );
  INVD1BWP30P140 U118 ( .I(n46), .ZN(n49) );
  INVD1BWP30P140 U119 ( .I(n50), .ZN(n47) );
  AN3D4BWP30P140 U120 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n47), .Z(n90) );
  OAI21D1BWP30P140 U121 ( .A1(n49), .A2(i_cmd[1]), .B(n48), .ZN(N354) );
  NR2D1BWP30P140 U122 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  MUX2NUD1BWP30P140 U123 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U124 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U125 ( .I(n55), .ZN(n78) );
  INVD1BWP30P140 U126 ( .I(n78), .ZN(n63) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  INVD2BWP30P140 U135 ( .I(n78), .ZN(n76) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_77 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  INVD2BWP30P140 U3 ( .I(n26), .ZN(n20) );
  INVD2BWP30P140 U4 ( .I(i_cmd[0]), .ZN(n21) );
  CKAN2D1BWP30P140 U5 ( .A1(i_valid[0]), .A2(n47), .Z(n46) );
  INVD1BWP30P140 U6 ( .I(n5), .ZN(n26) );
  ND2OPTIBD1BWP30P140 U7 ( .A1(n46), .A2(n21), .ZN(n5) );
  OAI22D1BWP30P140 U8 ( .A1(n44), .A2(n19), .B1(n20), .B2(n81), .ZN(N306) );
  ND2D1BWP30P140 U9 ( .A1(n1), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U10 ( .I(n90), .ZN(n48) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n17), .B1(n20), .B2(n80), .ZN(N307) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n16), .B1(n20), .B2(n78), .ZN(N308) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n15), .B1(n20), .B2(n77), .ZN(N309) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n14), .B1(n20), .B2(n73), .ZN(N310) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n13), .B1(n20), .B2(n72), .ZN(N311) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n12), .B1(n20), .B2(n71), .ZN(N312) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n11), .B1(n20), .B2(n70), .ZN(N313) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n10), .B1(n20), .B2(n69), .ZN(N314) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n9), .B1(n20), .B2(n68), .ZN(N315) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n8), .B1(n20), .B2(n67), .ZN(N316) );
  OAI22D1BWP30P140 U21 ( .A1(n18), .A2(n7), .B1(n20), .B2(n66), .ZN(N317) );
  OAI22D1BWP30P140 U22 ( .A1(n18), .A2(n6), .B1(n20), .B2(n65), .ZN(N318) );
  INVD1BWP30P140 U23 ( .I(rst), .ZN(n1) );
  NR2D1BWP30P140 U24 ( .A1(n50), .A2(n21), .ZN(n3) );
  INVD1BWP30P140 U25 ( .I(i_valid[0]), .ZN(n52) );
  INVD2BWP30P140 U26 ( .I(i_valid[1]), .ZN(n51) );
  MUX2NUD1BWP30P140 U27 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U28 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U29 ( .I(n4), .ZN(n22) );
  INVD2BWP30P140 U30 ( .I(n22), .ZN(n18) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[63]), .ZN(n6) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[31]), .ZN(n65) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[62]), .ZN(n7) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[30]), .ZN(n66) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[61]), .ZN(n8) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[29]), .ZN(n67) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[60]), .ZN(n9) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[28]), .ZN(n68) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[59]), .ZN(n10) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[58]), .ZN(n11) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[26]), .ZN(n70) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[57]), .ZN(n12) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[25]), .ZN(n71) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[56]), .ZN(n13) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[24]), .ZN(n72) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[55]), .ZN(n14) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[23]), .ZN(n73) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[54]), .ZN(n15) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[22]), .ZN(n77) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[53]), .ZN(n16) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[21]), .ZN(n78) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[52]), .ZN(n17) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD3BWP30P140 U55 ( .I(n22), .ZN(n44) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[51]), .ZN(n19) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[19]), .ZN(n81) );
  OAI31D1BWP30P140 U58 ( .A1(n50), .A2(n51), .A3(n21), .B(n20), .ZN(N353) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD2BWP30P140 U60 ( .I(n22), .ZN(n37) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[32]), .ZN(n23) );
  OAI22D1BWP30P140 U62 ( .A1(n45), .A2(n64), .B1(n37), .B2(n23), .ZN(N287) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[2]), .ZN(n61) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[34]), .ZN(n24) );
  OAI22D1BWP30P140 U65 ( .A1(n20), .A2(n61), .B1(n37), .B2(n24), .ZN(N289) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[35]), .ZN(n25) );
  OAI22D1BWP30P140 U68 ( .A1(n45), .A2(n60), .B1(n37), .B2(n25), .ZN(N290) );
  INVD2BWP30P140 U69 ( .I(n26), .ZN(n45) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[36]), .ZN(n27) );
  OAI22D1BWP30P140 U72 ( .A1(n45), .A2(n59), .B1(n37), .B2(n27), .ZN(N291) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[5]), .ZN(n58) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[37]), .ZN(n28) );
  OAI22D1BWP30P140 U75 ( .A1(n45), .A2(n58), .B1(n37), .B2(n28), .ZN(N292) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[6]), .ZN(n57) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[38]), .ZN(n29) );
  OAI22D1BWP30P140 U78 ( .A1(n45), .A2(n57), .B1(n37), .B2(n29), .ZN(N293) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[39]), .ZN(n30) );
  OAI22D1BWP30P140 U81 ( .A1(n45), .A2(n56), .B1(n37), .B2(n30), .ZN(N294) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[1]), .ZN(n62) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[33]), .ZN(n31) );
  OAI22D1BWP30P140 U84 ( .A1(n20), .A2(n62), .B1(n44), .B2(n31), .ZN(N288) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[16]), .ZN(n84) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[48]), .ZN(n32) );
  OAI22D1BWP30P140 U87 ( .A1(n45), .A2(n84), .B1(n44), .B2(n32), .ZN(N303) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[10]), .ZN(n92) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[42]), .ZN(n33) );
  OAI22D1BWP30P140 U90 ( .A1(n45), .A2(n92), .B1(n44), .B2(n33), .ZN(N297) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[11]), .ZN(n89) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[43]), .ZN(n34) );
  OAI22D1BWP30P140 U93 ( .A1(n45), .A2(n89), .B1(n44), .B2(n34), .ZN(N298) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[9]), .ZN(n76) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[41]), .ZN(n35) );
  OAI22D1BWP30P140 U96 ( .A1(n45), .A2(n76), .B1(n44), .B2(n35), .ZN(N296) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[8]), .ZN(n75) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[40]), .ZN(n36) );
  OAI22D1BWP30P140 U99 ( .A1(n45), .A2(n75), .B1(n37), .B2(n36), .ZN(N295) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[15]), .ZN(n85) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[47]), .ZN(n38) );
  OAI22D1BWP30P140 U102 ( .A1(n45), .A2(n85), .B1(n44), .B2(n38), .ZN(N302) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[14]), .ZN(n86) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[46]), .ZN(n39) );
  OAI22D1BWP30P140 U105 ( .A1(n45), .A2(n86), .B1(n44), .B2(n39), .ZN(N301) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[13]), .ZN(n87) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[45]), .ZN(n40) );
  OAI22D1BWP30P140 U108 ( .A1(n45), .A2(n87), .B1(n44), .B2(n40), .ZN(N300) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[12]), .ZN(n88) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[44]), .ZN(n41) );
  OAI22D1BWP30P140 U111 ( .A1(n45), .A2(n88), .B1(n44), .B2(n41), .ZN(N299) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[17]), .ZN(n83) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[49]), .ZN(n42) );
  OAI22D1BWP30P140 U114 ( .A1(n45), .A2(n83), .B1(n44), .B2(n42), .ZN(N304) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[18]), .ZN(n82) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[50]), .ZN(n43) );
  OAI22D1BWP30P140 U117 ( .A1(n45), .A2(n82), .B1(n44), .B2(n43), .ZN(N305) );
  INVD1BWP30P140 U118 ( .I(n46), .ZN(n49) );
  INVD1BWP30P140 U119 ( .I(n50), .ZN(n47) );
  AN3D4BWP30P140 U120 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n47), .Z(n90) );
  OAI21D1BWP30P140 U121 ( .A1(n49), .A2(i_cmd[1]), .B(n48), .ZN(N354) );
  NR2D1BWP30P140 U122 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  MUX2NUD1BWP30P140 U123 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U124 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U125 ( .I(n55), .ZN(n74) );
  INVD1BWP30P140 U126 ( .I(n74), .ZN(n63) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n63), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  INVD2BWP30P140 U135 ( .I(n74), .ZN(n79) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n79), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n79), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n79), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n79), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n79), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n79), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n79), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n79), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n79), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  INVD2BWP30P140 U145 ( .I(n74), .ZN(n91) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n79), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n79), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n79), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_78 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  INVD2BWP30P140 U3 ( .I(n27), .ZN(n20) );
  INVD2BWP30P140 U4 ( .I(i_cmd[0]), .ZN(n21) );
  CKAN2D1BWP30P140 U5 ( .A1(i_valid[0]), .A2(n47), .Z(n46) );
  INVD1BWP30P140 U6 ( .I(n5), .ZN(n27) );
  ND2OPTIBD1BWP30P140 U7 ( .A1(n46), .A2(n21), .ZN(n5) );
  ND2D1BWP30P140 U8 ( .A1(n1), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n48) );
  OAI22D1BWP30P140 U10 ( .A1(n44), .A2(n6), .B1(n20), .B2(n77), .ZN(N306) );
  OAI22D1BWP30P140 U11 ( .A1(n19), .A2(n7), .B1(n20), .B2(n79), .ZN(N307) );
  OAI22D1BWP30P140 U12 ( .A1(n19), .A2(n8), .B1(n20), .B2(n80), .ZN(N308) );
  OAI22D1BWP30P140 U13 ( .A1(n19), .A2(n9), .B1(n20), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U14 ( .A1(n19), .A2(n10), .B1(n20), .B2(n82), .ZN(N310) );
  OAI22D1BWP30P140 U15 ( .A1(n19), .A2(n11), .B1(n20), .B2(n92), .ZN(N311) );
  OAI22D1BWP30P140 U16 ( .A1(n19), .A2(n12), .B1(n20), .B2(n89), .ZN(N312) );
  OAI22D1BWP30P140 U17 ( .A1(n19), .A2(n13), .B1(n20), .B2(n88), .ZN(N313) );
  OAI22D1BWP30P140 U18 ( .A1(n19), .A2(n14), .B1(n20), .B2(n87), .ZN(N314) );
  OAI22D1BWP30P140 U19 ( .A1(n19), .A2(n15), .B1(n20), .B2(n86), .ZN(N315) );
  OAI22D1BWP30P140 U20 ( .A1(n19), .A2(n16), .B1(n20), .B2(n85), .ZN(N316) );
  OAI22D1BWP30P140 U21 ( .A1(n19), .A2(n17), .B1(n20), .B2(n84), .ZN(N317) );
  OAI22D1BWP30P140 U22 ( .A1(n19), .A2(n18), .B1(n20), .B2(n83), .ZN(N318) );
  INVD1BWP30P140 U23 ( .I(rst), .ZN(n1) );
  NR2D1BWP30P140 U24 ( .A1(n50), .A2(n21), .ZN(n3) );
  INVD1BWP30P140 U25 ( .I(i_valid[0]), .ZN(n52) );
  INVD2BWP30P140 U26 ( .I(i_valid[1]), .ZN(n51) );
  MUX2NUD1BWP30P140 U27 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U28 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U29 ( .I(n4), .ZN(n22) );
  INVD3BWP30P140 U30 ( .I(n22), .ZN(n44) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[51]), .ZN(n6) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[19]), .ZN(n77) );
  INVD2BWP30P140 U33 ( .I(n22), .ZN(n19) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[52]), .ZN(n7) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[20]), .ZN(n79) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[53]), .ZN(n8) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[54]), .ZN(n9) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[55]), .ZN(n10) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[23]), .ZN(n82) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[56]), .ZN(n11) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[24]), .ZN(n92) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[57]), .ZN(n12) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[25]), .ZN(n89) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[58]), .ZN(n13) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[26]), .ZN(n88) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[59]), .ZN(n14) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[27]), .ZN(n87) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[60]), .ZN(n15) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[28]), .ZN(n86) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[61]), .ZN(n16) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[29]), .ZN(n85) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[62]), .ZN(n17) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[30]), .ZN(n84) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[63]), .ZN(n18) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[31]), .ZN(n83) );
  OAI31D1BWP30P140 U58 ( .A1(n50), .A2(n51), .A3(n21), .B(n20), .ZN(N353) );
  INVD2BWP30P140 U59 ( .I(n27), .ZN(n45) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[7]), .ZN(n58) );
  INVD2BWP30P140 U61 ( .I(n22), .ZN(n37) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[39]), .ZN(n23) );
  OAI22D1BWP30P140 U63 ( .A1(n45), .A2(n58), .B1(n37), .B2(n23), .ZN(N294) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[6]), .ZN(n57) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[38]), .ZN(n24) );
  OAI22D1BWP30P140 U66 ( .A1(n45), .A2(n57), .B1(n37), .B2(n24), .ZN(N293) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[5]), .ZN(n64) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[37]), .ZN(n25) );
  OAI22D1BWP30P140 U69 ( .A1(n45), .A2(n64), .B1(n37), .B2(n25), .ZN(N292) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[4]), .ZN(n56) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[36]), .ZN(n26) );
  OAI22D1BWP30P140 U72 ( .A1(n45), .A2(n56), .B1(n37), .B2(n26), .ZN(N291) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[3]), .ZN(n59) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[35]), .ZN(n28) );
  OAI22D1BWP30P140 U75 ( .A1(n45), .A2(n59), .B1(n37), .B2(n28), .ZN(N290) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[34]), .ZN(n29) );
  OAI22D1BWP30P140 U78 ( .A1(n20), .A2(n60), .B1(n37), .B2(n29), .ZN(N289) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[1]), .ZN(n61) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[33]), .ZN(n30) );
  OAI22D1BWP30P140 U81 ( .A1(n45), .A2(n61), .B1(n37), .B2(n30), .ZN(N288) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[0]), .ZN(n62) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[32]), .ZN(n31) );
  OAI22D1BWP30P140 U84 ( .A1(n20), .A2(n62), .B1(n44), .B2(n31), .ZN(N287) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[8]), .ZN(n65) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[40]), .ZN(n32) );
  OAI22D1BWP30P140 U87 ( .A1(n45), .A2(n65), .B1(n44), .B2(n32), .ZN(N295) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[41]), .ZN(n33) );
  OAI22D1BWP30P140 U90 ( .A1(n45), .A2(n66), .B1(n44), .B2(n33), .ZN(N296) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[42]), .ZN(n34) );
  OAI22D1BWP30P140 U93 ( .A1(n45), .A2(n67), .B1(n44), .B2(n34), .ZN(N297) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[43]), .ZN(n35) );
  OAI22D1BWP30P140 U96 ( .A1(n45), .A2(n68), .B1(n44), .B2(n35), .ZN(N298) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[44]), .ZN(n36) );
  OAI22D1BWP30P140 U99 ( .A1(n45), .A2(n69), .B1(n37), .B2(n36), .ZN(N299) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[45]), .ZN(n38) );
  OAI22D1BWP30P140 U102 ( .A1(n45), .A2(n70), .B1(n44), .B2(n38), .ZN(N300) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[46]), .ZN(n39) );
  OAI22D1BWP30P140 U105 ( .A1(n45), .A2(n71), .B1(n44), .B2(n39), .ZN(N301) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[47]), .ZN(n40) );
  OAI22D1BWP30P140 U108 ( .A1(n45), .A2(n72), .B1(n44), .B2(n40), .ZN(N302) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[48]), .ZN(n41) );
  OAI22D1BWP30P140 U111 ( .A1(n45), .A2(n73), .B1(n44), .B2(n41), .ZN(N303) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[49]), .ZN(n42) );
  OAI22D1BWP30P140 U114 ( .A1(n45), .A2(n74), .B1(n44), .B2(n42), .ZN(N304) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[50]), .ZN(n43) );
  OAI22D1BWP30P140 U117 ( .A1(n45), .A2(n75), .B1(n44), .B2(n43), .ZN(N305) );
  INVD1BWP30P140 U118 ( .I(n46), .ZN(n49) );
  INVD1BWP30P140 U119 ( .I(n50), .ZN(n47) );
  AN3D4BWP30P140 U120 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n47), .Z(n90) );
  OAI21D1BWP30P140 U121 ( .A1(n49), .A2(i_cmd[1]), .B(n48), .ZN(N354) );
  NR2D1BWP30P140 U122 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  MUX2NUD1BWP30P140 U123 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U124 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U125 ( .I(n55), .ZN(n78) );
  INVD1BWP30P140 U126 ( .I(n78), .ZN(n63) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  INVD2BWP30P140 U135 ( .I(n78), .ZN(n76) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_79 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n45), .A2(n19), .B1(n20), .B2(n68), .ZN(N306) );
  INVD3BWP30P140 U4 ( .I(n25), .ZN(n20) );
  INVD1BWP30P140 U5 ( .I(n5), .ZN(n25) );
  ND2OPTIBD1BWP30P140 U6 ( .A1(n47), .A2(n21), .ZN(n5) );
  OAI22D1BWP30P140 U7 ( .A1(n18), .A2(n17), .B1(n20), .B2(n70), .ZN(N307) );
  OAI22D1BWP30P140 U8 ( .A1(n18), .A2(n16), .B1(n20), .B2(n71), .ZN(N308) );
  OAI22D1BWP30P140 U9 ( .A1(n18), .A2(n15), .B1(n20), .B2(n78), .ZN(N309) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n14), .B1(n20), .B2(n79), .ZN(N310) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n13), .B1(n20), .B2(n80), .ZN(N311) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n12), .B1(n20), .B2(n83), .ZN(N312) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n11), .B1(n20), .B2(n84), .ZN(N313) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n10), .B1(n20), .B2(n85), .ZN(N314) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n9), .B1(n20), .B2(n86), .ZN(N315) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n8), .B1(n20), .B2(n87), .ZN(N316) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n7), .B1(n20), .B2(n88), .ZN(N317) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n6), .B1(n20), .B2(n90), .ZN(N318) );
  ND2D1BWP30P140 U19 ( .A1(n1), .A2(i_en), .ZN(n51) );
  INVD1BWP30P140 U20 ( .I(n91), .ZN(n49) );
  INVD1BWP30P140 U21 ( .I(rst), .ZN(n1) );
  INVD1P5BWP30P140 U22 ( .I(i_cmd[0]), .ZN(n21) );
  NR2D1BWP30P140 U23 ( .A1(n51), .A2(n21), .ZN(n3) );
  INVD1BWP30P140 U24 ( .I(i_valid[0]), .ZN(n53) );
  INVD2BWP30P140 U25 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U26 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U27 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U28 ( .I(n4), .ZN(n22) );
  INVD2BWP30P140 U29 ( .I(n22), .ZN(n18) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[63]), .ZN(n6) );
  INR2D1BWP30P140 U31 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[31]), .ZN(n90) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[62]), .ZN(n7) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[30]), .ZN(n88) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[61]), .ZN(n8) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[29]), .ZN(n87) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[60]), .ZN(n9) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[28]), .ZN(n86) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[59]), .ZN(n10) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[27]), .ZN(n85) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[58]), .ZN(n11) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[26]), .ZN(n84) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[57]), .ZN(n12) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[25]), .ZN(n83) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[56]), .ZN(n13) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[24]), .ZN(n80) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[55]), .ZN(n14) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[23]), .ZN(n79) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[54]), .ZN(n15) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[22]), .ZN(n78) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[53]), .ZN(n16) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[21]), .ZN(n71) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[52]), .ZN(n17) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[20]), .ZN(n70) );
  INVD3BWP30P140 U55 ( .I(n22), .ZN(n45) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[51]), .ZN(n19) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[19]), .ZN(n68) );
  OAI31D1BWP30P140 U58 ( .A1(n51), .A2(n52), .A3(n21), .B(n20), .ZN(N353) );
  INVD1BWP30P140 U59 ( .I(n25), .ZN(n31) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD2BWP30P140 U61 ( .I(n22), .ZN(n38) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[32]), .ZN(n23) );
  OAI22D1BWP30P140 U63 ( .A1(n31), .A2(n57), .B1(n38), .B2(n23), .ZN(N287) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[33]), .ZN(n24) );
  OAI22D1BWP30P140 U66 ( .A1(n31), .A2(n58), .B1(n38), .B2(n24), .ZN(N288) );
  INVD2BWP30P140 U67 ( .I(n25), .ZN(n46) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[36]), .ZN(n26) );
  OAI22D1BWP30P140 U70 ( .A1(n46), .A2(n61), .B1(n38), .B2(n26), .ZN(N291) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[37]), .ZN(n27) );
  OAI22D1BWP30P140 U73 ( .A1(n46), .A2(n62), .B1(n38), .B2(n27), .ZN(N292) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[7]), .ZN(n65) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[39]), .ZN(n28) );
  OAI22D1BWP30P140 U76 ( .A1(n46), .A2(n65), .B1(n38), .B2(n28), .ZN(N294) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[34]), .ZN(n29) );
  OAI22D1BWP30P140 U79 ( .A1(n31), .A2(n59), .B1(n38), .B2(n29), .ZN(N289) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[35]), .ZN(n30) );
  OAI22D1BWP30P140 U82 ( .A1(n31), .A2(n60), .B1(n38), .B2(n30), .ZN(N290) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[38]), .ZN(n32) );
  OAI22D1BWP30P140 U85 ( .A1(n46), .A2(n63), .B1(n45), .B2(n32), .ZN(N293) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[18]), .ZN(n67) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[50]), .ZN(n33) );
  OAI22D1BWP30P140 U88 ( .A1(n46), .A2(n67), .B1(n45), .B2(n33), .ZN(N305) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[17]), .ZN(n93) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[49]), .ZN(n34) );
  OAI22D1BWP30P140 U91 ( .A1(n46), .A2(n93), .B1(n45), .B2(n34), .ZN(N304) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[16]), .ZN(n66) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[48]), .ZN(n35) );
  OAI22D1BWP30P140 U94 ( .A1(n46), .A2(n66), .B1(n45), .B2(n35), .ZN(N303) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[47]), .ZN(n36) );
  OAI22D1BWP30P140 U97 ( .A1(n46), .A2(n72), .B1(n45), .B2(n36), .ZN(N302) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[14]), .ZN(n73) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[46]), .ZN(n37) );
  OAI22D1BWP30P140 U100 ( .A1(n46), .A2(n73), .B1(n38), .B2(n37), .ZN(N301) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[13]), .ZN(n74) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[45]), .ZN(n39) );
  OAI22D1BWP30P140 U103 ( .A1(n46), .A2(n74), .B1(n45), .B2(n39), .ZN(N300) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[12]), .ZN(n75) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[44]), .ZN(n40) );
  OAI22D1BWP30P140 U106 ( .A1(n46), .A2(n75), .B1(n45), .B2(n40), .ZN(N299) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[11]), .ZN(n76) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[43]), .ZN(n41) );
  OAI22D1BWP30P140 U109 ( .A1(n46), .A2(n76), .B1(n45), .B2(n41), .ZN(N298) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[10]), .ZN(n77) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[42]), .ZN(n42) );
  OAI22D1BWP30P140 U112 ( .A1(n46), .A2(n77), .B1(n45), .B2(n42), .ZN(N297) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[9]), .ZN(n81) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[41]), .ZN(n43) );
  OAI22D1BWP30P140 U115 ( .A1(n46), .A2(n81), .B1(n45), .B2(n43), .ZN(N296) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[8]), .ZN(n82) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[40]), .ZN(n44) );
  OAI22D1BWP30P140 U118 ( .A1(n46), .A2(n82), .B1(n45), .B2(n44), .ZN(N295) );
  INVD1BWP30P140 U119 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U120 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U121 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n91) );
  OAI21D1BWP30P140 U122 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  NR2D1BWP30P140 U123 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  MUX2NUD1BWP30P140 U124 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n55), .A2(n54), .ZN(n56) );
  INVD2BWP30P140 U126 ( .I(n56), .ZN(n69) );
  INVD1BWP30P140 U127 ( .I(n69), .ZN(n64) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n64), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n64), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n64), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n64), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n64), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n64), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n64), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n64), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  INVD2BWP30P140 U136 ( .I(n69), .ZN(n92) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n92), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n92), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n92), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  INVD2BWP30P140 U140 ( .I(n69), .ZN(n89) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n89), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n89), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n92), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n92), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n92), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n92), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n92), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n92), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n89), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n89), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n89), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n92), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n92), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n89), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n89), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n85), .A2(n89), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n86), .A2(n89), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n87), .A2(n89), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n88), .A2(n89), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n89), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_80 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  INVD2BWP30P140 U3 ( .I(n24), .ZN(n20) );
  INVD2BWP30P140 U4 ( .I(i_cmd[0]), .ZN(n21) );
  CKAN2D1BWP30P140 U5 ( .A1(i_valid[0]), .A2(n47), .Z(n46) );
  INVD1BWP30P140 U6 ( .I(n5), .ZN(n24) );
  ND2OPTIBD1BWP30P140 U7 ( .A1(n46), .A2(n21), .ZN(n5) );
  ND2D1BWP30P140 U8 ( .A1(n1), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n48) );
  OAI22D1BWP30P140 U10 ( .A1(n44), .A2(n19), .B1(n20), .B2(n79), .ZN(N306) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n17), .B1(n20), .B2(n77), .ZN(N307) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n16), .B1(n20), .B2(n75), .ZN(N308) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n15), .B1(n20), .B2(n74), .ZN(N309) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n14), .B1(n20), .B2(n73), .ZN(N310) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n13), .B1(n20), .B2(n72), .ZN(N311) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n12), .B1(n20), .B2(n71), .ZN(N312) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n11), .B1(n20), .B2(n70), .ZN(N313) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n10), .B1(n20), .B2(n69), .ZN(N314) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n9), .B1(n20), .B2(n68), .ZN(N315) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n8), .B1(n20), .B2(n67), .ZN(N316) );
  OAI22D1BWP30P140 U21 ( .A1(n18), .A2(n7), .B1(n20), .B2(n66), .ZN(N317) );
  OAI22D1BWP30P140 U22 ( .A1(n18), .A2(n6), .B1(n20), .B2(n65), .ZN(N318) );
  INVD1BWP30P140 U23 ( .I(rst), .ZN(n1) );
  NR2D1BWP30P140 U24 ( .A1(n50), .A2(n21), .ZN(n3) );
  INVD1BWP30P140 U25 ( .I(i_valid[0]), .ZN(n52) );
  INVD2BWP30P140 U26 ( .I(i_valid[1]), .ZN(n51) );
  MUX2NUD1BWP30P140 U27 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U28 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U29 ( .I(n4), .ZN(n22) );
  INVD2BWP30P140 U30 ( .I(n22), .ZN(n18) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[63]), .ZN(n6) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[31]), .ZN(n65) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[62]), .ZN(n7) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[30]), .ZN(n66) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[61]), .ZN(n8) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[29]), .ZN(n67) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[60]), .ZN(n9) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[28]), .ZN(n68) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[59]), .ZN(n10) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[58]), .ZN(n11) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[26]), .ZN(n70) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[57]), .ZN(n12) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[25]), .ZN(n71) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[56]), .ZN(n13) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[24]), .ZN(n72) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[55]), .ZN(n14) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[23]), .ZN(n73) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[54]), .ZN(n15) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[53]), .ZN(n16) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[21]), .ZN(n75) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[52]), .ZN(n17) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD3BWP30P140 U55 ( .I(n22), .ZN(n44) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[51]), .ZN(n19) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[19]), .ZN(n79) );
  OAI31D1BWP30P140 U58 ( .A1(n50), .A2(n51), .A3(n21), .B(n20), .ZN(N353) );
  INVD2BWP30P140 U59 ( .I(n24), .ZN(n45) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[5]), .ZN(n58) );
  INVD2BWP30P140 U61 ( .I(n22), .ZN(n37) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[37]), .ZN(n23) );
  OAI22D1BWP30P140 U63 ( .A1(n45), .A2(n58), .B1(n37), .B2(n23), .ZN(N292) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[1]), .ZN(n62) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[33]), .ZN(n25) );
  OAI22D1BWP30P140 U66 ( .A1(n45), .A2(n62), .B1(n37), .B2(n25), .ZN(N288) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[36]), .ZN(n26) );
  OAI22D1BWP30P140 U69 ( .A1(n45), .A2(n59), .B1(n37), .B2(n26), .ZN(N291) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[32]), .ZN(n27) );
  OAI22D1BWP30P140 U72 ( .A1(n20), .A2(n64), .B1(n37), .B2(n27), .ZN(N287) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[6]), .ZN(n57) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[38]), .ZN(n28) );
  OAI22D1BWP30P140 U75 ( .A1(n45), .A2(n57), .B1(n37), .B2(n28), .ZN(N293) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[35]), .ZN(n29) );
  OAI22D1BWP30P140 U78 ( .A1(n45), .A2(n60), .B1(n37), .B2(n29), .ZN(N290) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[2]), .ZN(n61) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[34]), .ZN(n30) );
  OAI22D1BWP30P140 U81 ( .A1(n20), .A2(n61), .B1(n37), .B2(n30), .ZN(N289) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[39]), .ZN(n31) );
  OAI22D1BWP30P140 U84 ( .A1(n45), .A2(n56), .B1(n44), .B2(n31), .ZN(N294) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[18]), .ZN(n80) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[50]), .ZN(n32) );
  OAI22D1BWP30P140 U87 ( .A1(n45), .A2(n80), .B1(n44), .B2(n32), .ZN(N305) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[17]), .ZN(n81) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[49]), .ZN(n33) );
  OAI22D1BWP30P140 U90 ( .A1(n45), .A2(n81), .B1(n44), .B2(n33), .ZN(N304) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[16]), .ZN(n82) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[48]), .ZN(n34) );
  OAI22D1BWP30P140 U93 ( .A1(n45), .A2(n82), .B1(n44), .B2(n34), .ZN(N303) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[15]), .ZN(n83) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[47]), .ZN(n35) );
  OAI22D1BWP30P140 U96 ( .A1(n45), .A2(n83), .B1(n44), .B2(n35), .ZN(N302) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[14]), .ZN(n84) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[46]), .ZN(n36) );
  OAI22D1BWP30P140 U99 ( .A1(n45), .A2(n84), .B1(n37), .B2(n36), .ZN(N301) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[44]), .ZN(n38) );
  OAI22D1BWP30P140 U102 ( .A1(n45), .A2(n86), .B1(n44), .B2(n38), .ZN(N299) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[11]), .ZN(n87) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[43]), .ZN(n39) );
  OAI22D1BWP30P140 U105 ( .A1(n45), .A2(n87), .B1(n44), .B2(n39), .ZN(N298) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[42]), .ZN(n40) );
  OAI22D1BWP30P140 U108 ( .A1(n45), .A2(n88), .B1(n44), .B2(n40), .ZN(N297) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[9]), .ZN(n89) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[41]), .ZN(n41) );
  OAI22D1BWP30P140 U111 ( .A1(n45), .A2(n89), .B1(n44), .B2(n41), .ZN(N296) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[8]), .ZN(n92) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[40]), .ZN(n42) );
  OAI22D1BWP30P140 U114 ( .A1(n45), .A2(n92), .B1(n44), .B2(n42), .ZN(N295) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[13]), .ZN(n85) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[45]), .ZN(n43) );
  OAI22D1BWP30P140 U117 ( .A1(n45), .A2(n85), .B1(n44), .B2(n43), .ZN(N300) );
  INVD1BWP30P140 U118 ( .I(n46), .ZN(n49) );
  INVD1BWP30P140 U119 ( .I(n50), .ZN(n47) );
  AN3D4BWP30P140 U120 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n47), .Z(n90) );
  OAI21D1BWP30P140 U121 ( .A1(n49), .A2(i_cmd[1]), .B(n48), .ZN(N354) );
  NR2D1BWP30P140 U122 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  MUX2NUD1BWP30P140 U123 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U124 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U125 ( .I(n55), .ZN(n78) );
  INVD1BWP30P140 U126 ( .I(n78), .ZN(n63) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n63), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  INVD2BWP30P140 U135 ( .I(n78), .ZN(n76) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n76), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n76), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n76), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n76), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n76), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n76), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n76), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n76), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n76), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n76), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n76), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U147 ( .A1(n77), .A2(n76), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  INVD2BWP30P140 U148 ( .I(n78), .ZN(n91) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_81 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n45), .A2(n19), .B1(n20), .B2(n86), .ZN(N306) );
  INVD3BWP30P140 U4 ( .I(n27), .ZN(n20) );
  INVD1BWP30P140 U5 ( .I(n5), .ZN(n27) );
  ND2OPTIBD1BWP30P140 U6 ( .A1(n47), .A2(n21), .ZN(n5) );
  OAI22D1BWP30P140 U7 ( .A1(n18), .A2(n17), .B1(n20), .B2(n77), .ZN(N307) );
  OAI22D1BWP30P140 U8 ( .A1(n18), .A2(n16), .B1(n20), .B2(n76), .ZN(N308) );
  OAI22D1BWP30P140 U9 ( .A1(n18), .A2(n15), .B1(n20), .B2(n75), .ZN(N309) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n14), .B1(n20), .B2(n74), .ZN(N310) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n13), .B1(n20), .B2(n69), .ZN(N311) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n12), .B1(n20), .B2(n68), .ZN(N312) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n11), .B1(n20), .B2(n67), .ZN(N313) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n10), .B1(n20), .B2(n66), .ZN(N314) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n9), .B1(n20), .B2(n73), .ZN(N315) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n8), .B1(n20), .B2(n72), .ZN(N316) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n7), .B1(n20), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n6), .B1(n20), .B2(n87), .ZN(N318) );
  ND2D1BWP30P140 U19 ( .A1(n1), .A2(i_en), .ZN(n51) );
  INVD1BWP30P140 U20 ( .I(n91), .ZN(n49) );
  INVD1BWP30P140 U21 ( .I(rst), .ZN(n1) );
  INVD1P5BWP30P140 U22 ( .I(i_cmd[0]), .ZN(n21) );
  NR2D1BWP30P140 U23 ( .A1(n51), .A2(n21), .ZN(n3) );
  INVD1BWP30P140 U24 ( .I(i_valid[0]), .ZN(n53) );
  INVD2BWP30P140 U25 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U26 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U27 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U28 ( .I(n4), .ZN(n22) );
  INVD2BWP30P140 U29 ( .I(n22), .ZN(n18) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[63]), .ZN(n6) );
  INR2D1BWP30P140 U31 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[31]), .ZN(n87) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[62]), .ZN(n7) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[61]), .ZN(n8) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[29]), .ZN(n72) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[60]), .ZN(n9) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[28]), .ZN(n73) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[59]), .ZN(n10) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[27]), .ZN(n66) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[58]), .ZN(n11) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[26]), .ZN(n67) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[57]), .ZN(n12) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[25]), .ZN(n68) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[56]), .ZN(n13) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[24]), .ZN(n69) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[55]), .ZN(n14) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[23]), .ZN(n74) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[54]), .ZN(n15) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[22]), .ZN(n75) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[53]), .ZN(n16) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[21]), .ZN(n76) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[52]), .ZN(n17) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD3BWP30P140 U55 ( .I(n22), .ZN(n45) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[51]), .ZN(n19) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[19]), .ZN(n86) );
  OAI31D1BWP30P140 U58 ( .A1(n51), .A2(n52), .A3(n21), .B(n20), .ZN(N353) );
  INVD2BWP30P140 U59 ( .I(n27), .ZN(n46) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[7]), .ZN(n65) );
  INVD2BWP30P140 U61 ( .I(n22), .ZN(n38) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[39]), .ZN(n23) );
  OAI22D1BWP30P140 U63 ( .A1(n46), .A2(n65), .B1(n38), .B2(n23), .ZN(N294) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[38]), .ZN(n24) );
  OAI22D1BWP30P140 U66 ( .A1(n46), .A2(n63), .B1(n38), .B2(n24), .ZN(N293) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[37]), .ZN(n25) );
  OAI22D1BWP30P140 U69 ( .A1(n46), .A2(n62), .B1(n38), .B2(n25), .ZN(N292) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[36]), .ZN(n26) );
  OAI22D1BWP30P140 U72 ( .A1(n46), .A2(n61), .B1(n38), .B2(n26), .ZN(N291) );
  INVD1BWP30P140 U73 ( .I(n27), .ZN(n32) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[35]), .ZN(n28) );
  OAI22D1BWP30P140 U76 ( .A1(n32), .A2(n60), .B1(n38), .B2(n28), .ZN(N290) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[34]), .ZN(n29) );
  OAI22D1BWP30P140 U79 ( .A1(n32), .A2(n59), .B1(n38), .B2(n29), .ZN(N289) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[33]), .ZN(n30) );
  OAI22D1BWP30P140 U82 ( .A1(n32), .A2(n58), .B1(n38), .B2(n30), .ZN(N288) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[32]), .ZN(n31) );
  OAI22D1BWP30P140 U85 ( .A1(n32), .A2(n57), .B1(n45), .B2(n31), .ZN(N287) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[18]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[50]), .ZN(n33) );
  OAI22D1BWP30P140 U88 ( .A1(n46), .A2(n85), .B1(n45), .B2(n33), .ZN(N305) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[17]), .ZN(n84) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[49]), .ZN(n34) );
  OAI22D1BWP30P140 U91 ( .A1(n46), .A2(n84), .B1(n45), .B2(n34), .ZN(N304) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[16]), .ZN(n83) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[48]), .ZN(n35) );
  OAI22D1BWP30P140 U94 ( .A1(n46), .A2(n83), .B1(n45), .B2(n35), .ZN(N303) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[15]), .ZN(n82) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[47]), .ZN(n36) );
  OAI22D1BWP30P140 U97 ( .A1(n46), .A2(n82), .B1(n45), .B2(n36), .ZN(N302) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[14]), .ZN(n81) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[46]), .ZN(n37) );
  OAI22D1BWP30P140 U100 ( .A1(n46), .A2(n81), .B1(n38), .B2(n37), .ZN(N301) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[13]), .ZN(n80) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[45]), .ZN(n39) );
  OAI22D1BWP30P140 U103 ( .A1(n46), .A2(n80), .B1(n45), .B2(n39), .ZN(N300) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[12]), .ZN(n79) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[44]), .ZN(n40) );
  OAI22D1BWP30P140 U106 ( .A1(n46), .A2(n79), .B1(n45), .B2(n40), .ZN(N299) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[11]), .ZN(n78) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[43]), .ZN(n41) );
  OAI22D1BWP30P140 U109 ( .A1(n46), .A2(n78), .B1(n45), .B2(n41), .ZN(N298) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[10]), .ZN(n71) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[42]), .ZN(n42) );
  OAI22D1BWP30P140 U112 ( .A1(n46), .A2(n71), .B1(n45), .B2(n42), .ZN(N297) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[9]), .ZN(n90) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[41]), .ZN(n43) );
  OAI22D1BWP30P140 U115 ( .A1(n46), .A2(n90), .B1(n45), .B2(n43), .ZN(N296) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[8]), .ZN(n93) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[40]), .ZN(n44) );
  OAI22D1BWP30P140 U118 ( .A1(n46), .A2(n93), .B1(n45), .B2(n44), .ZN(N295) );
  INVD1BWP30P140 U119 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U120 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U121 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n91) );
  OAI21D1BWP30P140 U122 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  NR2D1BWP30P140 U123 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  MUX2NUD1BWP30P140 U124 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n55), .A2(n54), .ZN(n56) );
  INVD2BWP30P140 U126 ( .I(n56), .ZN(n70) );
  INVD1BWP30P140 U127 ( .I(n70), .ZN(n64) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n64), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n64), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n64), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n64), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n64), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n64), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n64), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n64), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  INVD2BWP30P140 U136 ( .I(n70), .ZN(n88) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n88), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n88), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n88), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n88), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  INVD2BWP30P140 U141 ( .I(n70), .ZN(n92) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n92), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n88), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n88), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n88), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n88), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n88), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n88), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n92), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n92), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n92), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n92), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n92), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n92), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n92), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U156 ( .A1(n85), .A2(n92), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U157 ( .A1(n86), .A2(n92), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U158 ( .A1(n87), .A2(n88), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n88), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_82 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  INVD2BWP30P140 U3 ( .I(n27), .ZN(n20) );
  INVD2BWP30P140 U4 ( .I(i_cmd[0]), .ZN(n21) );
  CKAN2D1BWP30P140 U5 ( .A1(i_valid[0]), .A2(n47), .Z(n46) );
  INVD1BWP30P140 U6 ( .I(n5), .ZN(n27) );
  ND2OPTIBD1BWP30P140 U7 ( .A1(n46), .A2(n21), .ZN(n5) );
  ND2D1BWP30P140 U8 ( .A1(n1), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n48) );
  OAI22D1BWP30P140 U10 ( .A1(n44), .A2(n19), .B1(n20), .B2(n92), .ZN(N306) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n17), .B1(n20), .B2(n89), .ZN(N307) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n16), .B1(n20), .B2(n83), .ZN(N308) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n15), .B1(n20), .B2(n79), .ZN(N309) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n14), .B1(n20), .B2(n78), .ZN(N310) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n13), .B1(n20), .B2(n77), .ZN(N311) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n12), .B1(n20), .B2(n76), .ZN(N312) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n11), .B1(n20), .B2(n75), .ZN(N313) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n10), .B1(n20), .B2(n74), .ZN(N314) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n9), .B1(n20), .B2(n73), .ZN(N315) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n8), .B1(n20), .B2(n72), .ZN(N316) );
  OAI22D1BWP30P140 U21 ( .A1(n18), .A2(n7), .B1(n20), .B2(n70), .ZN(N317) );
  OAI22D1BWP30P140 U22 ( .A1(n18), .A2(n6), .B1(n20), .B2(n69), .ZN(N318) );
  INVD1BWP30P140 U23 ( .I(rst), .ZN(n1) );
  NR2D1BWP30P140 U24 ( .A1(n50), .A2(n21), .ZN(n3) );
  INVD1BWP30P140 U25 ( .I(i_valid[0]), .ZN(n52) );
  INVD2BWP30P140 U26 ( .I(i_valid[1]), .ZN(n51) );
  MUX2NUD1BWP30P140 U27 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U28 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U29 ( .I(n4), .ZN(n22) );
  INVD2BWP30P140 U30 ( .I(n22), .ZN(n18) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[63]), .ZN(n6) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[31]), .ZN(n69) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[62]), .ZN(n7) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[30]), .ZN(n70) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[61]), .ZN(n8) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[29]), .ZN(n72) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[60]), .ZN(n9) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[28]), .ZN(n73) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[59]), .ZN(n10) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[27]), .ZN(n74) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[58]), .ZN(n11) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[26]), .ZN(n75) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[57]), .ZN(n12) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[25]), .ZN(n76) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[56]), .ZN(n13) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[24]), .ZN(n77) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[55]), .ZN(n14) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[23]), .ZN(n78) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[54]), .ZN(n15) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[22]), .ZN(n79) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[53]), .ZN(n16) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[21]), .ZN(n83) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[52]), .ZN(n17) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[20]), .ZN(n89) );
  INVD3BWP30P140 U55 ( .I(n22), .ZN(n44) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[51]), .ZN(n19) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[19]), .ZN(n92) );
  OAI31D1BWP30P140 U58 ( .A1(n50), .A2(n51), .A3(n21), .B(n20), .ZN(N353) );
  INVD2BWP30P140 U59 ( .I(n27), .ZN(n45) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD2BWP30P140 U61 ( .I(n22), .ZN(n37) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[39]), .ZN(n23) );
  OAI22D1BWP30P140 U63 ( .A1(n45), .A2(n56), .B1(n37), .B2(n23), .ZN(N294) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[6]), .ZN(n57) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[38]), .ZN(n24) );
  OAI22D1BWP30P140 U66 ( .A1(n45), .A2(n57), .B1(n37), .B2(n24), .ZN(N293) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[5]), .ZN(n58) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[37]), .ZN(n25) );
  OAI22D1BWP30P140 U69 ( .A1(n45), .A2(n58), .B1(n37), .B2(n25), .ZN(N292) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[36]), .ZN(n26) );
  OAI22D1BWP30P140 U72 ( .A1(n45), .A2(n59), .B1(n37), .B2(n26), .ZN(N291) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[35]), .ZN(n28) );
  OAI22D1BWP30P140 U75 ( .A1(n45), .A2(n60), .B1(n37), .B2(n28), .ZN(N290) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[2]), .ZN(n61) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[34]), .ZN(n29) );
  OAI22D1BWP30P140 U78 ( .A1(n20), .A2(n61), .B1(n37), .B2(n29), .ZN(N289) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[1]), .ZN(n62) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[33]), .ZN(n30) );
  OAI22D1BWP30P140 U81 ( .A1(n45), .A2(n62), .B1(n37), .B2(n30), .ZN(N288) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[32]), .ZN(n31) );
  OAI22D1BWP30P140 U84 ( .A1(n20), .A2(n64), .B1(n44), .B2(n31), .ZN(N287) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[18]), .ZN(n84) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[50]), .ZN(n32) );
  OAI22D1BWP30P140 U87 ( .A1(n45), .A2(n84), .B1(n44), .B2(n32), .ZN(N305) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[17]), .ZN(n87) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[49]), .ZN(n33) );
  OAI22D1BWP30P140 U90 ( .A1(n45), .A2(n87), .B1(n44), .B2(n33), .ZN(N304) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[16]), .ZN(n86) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[48]), .ZN(n34) );
  OAI22D1BWP30P140 U93 ( .A1(n45), .A2(n86), .B1(n44), .B2(n34), .ZN(N303) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[15]), .ZN(n82) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[47]), .ZN(n35) );
  OAI22D1BWP30P140 U96 ( .A1(n45), .A2(n82), .B1(n44), .B2(n35), .ZN(N302) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[14]), .ZN(n85) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[46]), .ZN(n36) );
  OAI22D1BWP30P140 U99 ( .A1(n45), .A2(n85), .B1(n37), .B2(n36), .ZN(N301) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[13]), .ZN(n81) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[45]), .ZN(n38) );
  OAI22D1BWP30P140 U102 ( .A1(n45), .A2(n81), .B1(n44), .B2(n38), .ZN(N300) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[12]), .ZN(n80) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[44]), .ZN(n39) );
  OAI22D1BWP30P140 U105 ( .A1(n45), .A2(n80), .B1(n44), .B2(n39), .ZN(N299) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[11]), .ZN(n65) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[43]), .ZN(n40) );
  OAI22D1BWP30P140 U108 ( .A1(n45), .A2(n65), .B1(n44), .B2(n40), .ZN(N298) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[10]), .ZN(n66) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[42]), .ZN(n41) );
  OAI22D1BWP30P140 U111 ( .A1(n45), .A2(n66), .B1(n44), .B2(n41), .ZN(N297) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[9]), .ZN(n67) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[41]), .ZN(n42) );
  OAI22D1BWP30P140 U114 ( .A1(n45), .A2(n67), .B1(n44), .B2(n42), .ZN(N296) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[8]), .ZN(n71) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[40]), .ZN(n43) );
  OAI22D1BWP30P140 U117 ( .A1(n45), .A2(n71), .B1(n44), .B2(n43), .ZN(N295) );
  INVD1BWP30P140 U118 ( .I(n46), .ZN(n49) );
  INVD1BWP30P140 U119 ( .I(n50), .ZN(n47) );
  AN3D4BWP30P140 U120 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n47), .Z(n90) );
  OAI21D1BWP30P140 U121 ( .A1(n49), .A2(i_cmd[1]), .B(n48), .ZN(N354) );
  NR2D1BWP30P140 U122 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  MUX2NUD1BWP30P140 U123 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U124 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U125 ( .I(n55), .ZN(n68) );
  INVD1BWP30P140 U126 ( .I(n68), .ZN(n63) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n63), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  INVD2BWP30P140 U135 ( .I(n68), .ZN(n91) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  INVD2BWP30P140 U139 ( .I(n68), .ZN(n88) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n88), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n88), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n88), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n88), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n88), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n88), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n88), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n88), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n88), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n88), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n88), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U156 ( .A1(n85), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U157 ( .A1(n86), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U158 ( .A1(n87), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n88), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_83 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n45), .A2(n19), .B1(n20), .B2(n80), .ZN(N306) );
  INVD3BWP30P140 U4 ( .I(n27), .ZN(n20) );
  INVD1BWP30P140 U5 ( .I(n5), .ZN(n27) );
  ND2OPTIBD1BWP30P140 U6 ( .A1(n47), .A2(n21), .ZN(n5) );
  OAI22D1BWP30P140 U7 ( .A1(n18), .A2(n17), .B1(n20), .B2(n81), .ZN(N307) );
  OAI22D1BWP30P140 U8 ( .A1(n18), .A2(n16), .B1(n20), .B2(n82), .ZN(N308) );
  OAI22D1BWP30P140 U9 ( .A1(n18), .A2(n15), .B1(n20), .B2(n83), .ZN(N309) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n14), .B1(n20), .B2(n85), .ZN(N310) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n13), .B1(n20), .B2(n66), .ZN(N311) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n12), .B1(n20), .B2(n67), .ZN(N312) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n11), .B1(n20), .B2(n68), .ZN(N313) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n10), .B1(n20), .B2(n69), .ZN(N314) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n9), .B1(n20), .B2(n70), .ZN(N315) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n8), .B1(n20), .B2(n71), .ZN(N316) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n7), .B1(n20), .B2(n72), .ZN(N317) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n6), .B1(n20), .B2(n73), .ZN(N318) );
  ND2D1BWP30P140 U19 ( .A1(n1), .A2(i_en), .ZN(n51) );
  INVD1BWP30P140 U20 ( .I(n91), .ZN(n49) );
  INVD1BWP30P140 U21 ( .I(rst), .ZN(n1) );
  INVD1P5BWP30P140 U22 ( .I(i_cmd[0]), .ZN(n21) );
  NR2D1BWP30P140 U23 ( .A1(n51), .A2(n21), .ZN(n3) );
  INVD1BWP30P140 U24 ( .I(i_valid[0]), .ZN(n53) );
  INVD2BWP30P140 U25 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U26 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U27 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U28 ( .I(n4), .ZN(n22) );
  INVD2BWP30P140 U29 ( .I(n22), .ZN(n18) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[63]), .ZN(n6) );
  INR2D1BWP30P140 U31 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[31]), .ZN(n73) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[62]), .ZN(n7) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[30]), .ZN(n72) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[61]), .ZN(n8) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[29]), .ZN(n71) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[60]), .ZN(n9) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[28]), .ZN(n70) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[59]), .ZN(n10) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[58]), .ZN(n11) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[26]), .ZN(n68) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[57]), .ZN(n12) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[25]), .ZN(n67) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[56]), .ZN(n13) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[24]), .ZN(n66) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[55]), .ZN(n14) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[23]), .ZN(n85) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[54]), .ZN(n15) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[22]), .ZN(n83) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[53]), .ZN(n16) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[21]), .ZN(n82) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[52]), .ZN(n17) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[20]), .ZN(n81) );
  INVD3BWP30P140 U55 ( .I(n22), .ZN(n45) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[51]), .ZN(n19) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[19]), .ZN(n80) );
  OAI31D1BWP30P140 U58 ( .A1(n51), .A2(n52), .A3(n21), .B(n20), .ZN(N353) );
  INVD2BWP30P140 U59 ( .I(n27), .ZN(n46) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[7]), .ZN(n61) );
  INVD2BWP30P140 U61 ( .I(n22), .ZN(n38) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[39]), .ZN(n23) );
  OAI22D1BWP30P140 U63 ( .A1(n46), .A2(n61), .B1(n38), .B2(n23), .ZN(N294) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[6]), .ZN(n62) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[38]), .ZN(n24) );
  OAI22D1BWP30P140 U66 ( .A1(n46), .A2(n62), .B1(n38), .B2(n24), .ZN(N293) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[5]), .ZN(n63) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[37]), .ZN(n25) );
  OAI22D1BWP30P140 U69 ( .A1(n46), .A2(n63), .B1(n38), .B2(n25), .ZN(N292) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[4]), .ZN(n65) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[36]), .ZN(n26) );
  OAI22D1BWP30P140 U72 ( .A1(n46), .A2(n65), .B1(n38), .B2(n26), .ZN(N291) );
  INVD1BWP30P140 U73 ( .I(n27), .ZN(n32) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[3]), .ZN(n57) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[35]), .ZN(n28) );
  OAI22D1BWP30P140 U76 ( .A1(n32), .A2(n57), .B1(n38), .B2(n28), .ZN(N290) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[34]), .ZN(n29) );
  OAI22D1BWP30P140 U79 ( .A1(n32), .A2(n60), .B1(n38), .B2(n29), .ZN(N289) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[33]), .ZN(n30) );
  OAI22D1BWP30P140 U82 ( .A1(n32), .A2(n59), .B1(n38), .B2(n30), .ZN(N288) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[0]), .ZN(n58) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[32]), .ZN(n31) );
  OAI22D1BWP30P140 U85 ( .A1(n32), .A2(n58), .B1(n45), .B2(n31), .ZN(N287) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[18]), .ZN(n79) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[50]), .ZN(n33) );
  OAI22D1BWP30P140 U88 ( .A1(n46), .A2(n79), .B1(n45), .B2(n33), .ZN(N305) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[17]), .ZN(n78) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[49]), .ZN(n34) );
  OAI22D1BWP30P140 U91 ( .A1(n46), .A2(n78), .B1(n45), .B2(n34), .ZN(N304) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[16]), .ZN(n77) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[48]), .ZN(n35) );
  OAI22D1BWP30P140 U94 ( .A1(n46), .A2(n77), .B1(n45), .B2(n35), .ZN(N303) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[15]), .ZN(n76) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[47]), .ZN(n36) );
  OAI22D1BWP30P140 U97 ( .A1(n46), .A2(n76), .B1(n45), .B2(n36), .ZN(N302) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[14]), .ZN(n75) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[46]), .ZN(n37) );
  OAI22D1BWP30P140 U100 ( .A1(n46), .A2(n75), .B1(n38), .B2(n37), .ZN(N301) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[13]), .ZN(n86) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[45]), .ZN(n39) );
  OAI22D1BWP30P140 U103 ( .A1(n46), .A2(n86), .B1(n45), .B2(n39), .ZN(N300) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[12]), .ZN(n87) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[44]), .ZN(n40) );
  OAI22D1BWP30P140 U106 ( .A1(n46), .A2(n87), .B1(n45), .B2(n40), .ZN(N299) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[11]), .ZN(n88) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[43]), .ZN(n41) );
  OAI22D1BWP30P140 U109 ( .A1(n46), .A2(n88), .B1(n45), .B2(n41), .ZN(N298) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[10]), .ZN(n89) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[42]), .ZN(n42) );
  OAI22D1BWP30P140 U112 ( .A1(n46), .A2(n89), .B1(n45), .B2(n42), .ZN(N297) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[9]), .ZN(n90) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[41]), .ZN(n43) );
  OAI22D1BWP30P140 U115 ( .A1(n46), .A2(n90), .B1(n45), .B2(n43), .ZN(N296) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[8]), .ZN(n93) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[40]), .ZN(n44) );
  OAI22D1BWP30P140 U118 ( .A1(n46), .A2(n93), .B1(n45), .B2(n44), .ZN(N295) );
  INVD1BWP30P140 U119 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U120 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U121 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n91) );
  OAI21D1BWP30P140 U122 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  NR2D1BWP30P140 U123 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  MUX2NUD1BWP30P140 U124 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n55), .A2(n54), .ZN(n56) );
  INVD2BWP30P140 U126 ( .I(n56), .ZN(n74) );
  INVD1BWP30P140 U127 ( .I(n74), .ZN(n64) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n64), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n64), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n64), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n64), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n64), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n64), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n64), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n64), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  INVD2BWP30P140 U136 ( .I(n74), .ZN(n84) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n84), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n84), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n84), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n84), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n84), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n84), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n84), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n84), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
  INVD2BWP30P140 U145 ( .I(n74), .ZN(n92) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n92), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n92), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n92), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n92), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n92), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n92), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n84), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n84), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n84), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n84), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_84 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  INVD2BWP30P140 U3 ( .I(n27), .ZN(n20) );
  INVD2BWP30P140 U4 ( .I(i_cmd[0]), .ZN(n21) );
  CKAN2D1BWP30P140 U5 ( .A1(i_valid[0]), .A2(n47), .Z(n46) );
  INVD1BWP30P140 U6 ( .I(n5), .ZN(n27) );
  ND2OPTIBD1BWP30P140 U7 ( .A1(n46), .A2(n21), .ZN(n5) );
  ND2D1BWP30P140 U8 ( .A1(n1), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U9 ( .I(n90), .ZN(n48) );
  OAI22D1BWP30P140 U10 ( .A1(n44), .A2(n19), .B1(n20), .B2(n81), .ZN(N306) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n17), .B1(n20), .B2(n80), .ZN(N307) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n16), .B1(n20), .B2(n78), .ZN(N308) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n15), .B1(n20), .B2(n77), .ZN(N309) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n14), .B1(n20), .B2(n76), .ZN(N310) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n13), .B1(n20), .B2(n75), .ZN(N311) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n12), .B1(n20), .B2(n74), .ZN(N312) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n11), .B1(n20), .B2(n70), .ZN(N313) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n10), .B1(n20), .B2(n69), .ZN(N314) );
  OAI22D1BWP30P140 U19 ( .A1(n18), .A2(n9), .B1(n20), .B2(n68), .ZN(N315) );
  OAI22D1BWP30P140 U20 ( .A1(n18), .A2(n8), .B1(n20), .B2(n67), .ZN(N316) );
  OAI22D1BWP30P140 U21 ( .A1(n18), .A2(n7), .B1(n20), .B2(n66), .ZN(N317) );
  OAI22D1BWP30P140 U22 ( .A1(n18), .A2(n6), .B1(n20), .B2(n65), .ZN(N318) );
  INVD1BWP30P140 U23 ( .I(rst), .ZN(n1) );
  NR2D1BWP30P140 U24 ( .A1(n50), .A2(n21), .ZN(n3) );
  INVD1BWP30P140 U25 ( .I(i_valid[0]), .ZN(n52) );
  INVD2BWP30P140 U26 ( .I(i_valid[1]), .ZN(n51) );
  MUX2NUD1BWP30P140 U27 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U28 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U29 ( .I(n4), .ZN(n22) );
  INVD2BWP30P140 U30 ( .I(n22), .ZN(n18) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[63]), .ZN(n6) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[31]), .ZN(n65) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[62]), .ZN(n7) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[30]), .ZN(n66) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[61]), .ZN(n8) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[29]), .ZN(n67) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[60]), .ZN(n9) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[28]), .ZN(n68) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[59]), .ZN(n10) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[58]), .ZN(n11) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[26]), .ZN(n70) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[57]), .ZN(n12) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[25]), .ZN(n74) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[56]), .ZN(n13) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[24]), .ZN(n75) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[55]), .ZN(n14) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[23]), .ZN(n76) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[54]), .ZN(n15) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[22]), .ZN(n77) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[53]), .ZN(n16) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[21]), .ZN(n78) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[52]), .ZN(n17) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD3BWP30P140 U55 ( .I(n22), .ZN(n44) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[51]), .ZN(n19) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[19]), .ZN(n81) );
  OAI31D1BWP30P140 U58 ( .A1(n50), .A2(n51), .A3(n21), .B(n20), .ZN(N353) );
  INVD2BWP30P140 U59 ( .I(n27), .ZN(n45) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD2BWP30P140 U61 ( .I(n22), .ZN(n37) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[39]), .ZN(n23) );
  OAI22D1BWP30P140 U63 ( .A1(n45), .A2(n57), .B1(n37), .B2(n23), .ZN(N294) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[6]), .ZN(n56) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[38]), .ZN(n24) );
  OAI22D1BWP30P140 U66 ( .A1(n45), .A2(n56), .B1(n37), .B2(n24), .ZN(N293) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[5]), .ZN(n58) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[37]), .ZN(n25) );
  OAI22D1BWP30P140 U69 ( .A1(n45), .A2(n58), .B1(n37), .B2(n25), .ZN(N292) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[36]), .ZN(n26) );
  OAI22D1BWP30P140 U72 ( .A1(n45), .A2(n59), .B1(n37), .B2(n26), .ZN(N291) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[3]), .ZN(n64) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[35]), .ZN(n28) );
  OAI22D1BWP30P140 U75 ( .A1(n45), .A2(n64), .B1(n37), .B2(n28), .ZN(N290) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[34]), .ZN(n29) );
  OAI22D1BWP30P140 U78 ( .A1(n20), .A2(n60), .B1(n37), .B2(n29), .ZN(N289) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[1]), .ZN(n61) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[33]), .ZN(n30) );
  OAI22D1BWP30P140 U81 ( .A1(n45), .A2(n61), .B1(n37), .B2(n30), .ZN(N288) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[0]), .ZN(n62) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[32]), .ZN(n31) );
  OAI22D1BWP30P140 U84 ( .A1(n20), .A2(n62), .B1(n44), .B2(n31), .ZN(N287) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[18]), .ZN(n82) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[50]), .ZN(n32) );
  OAI22D1BWP30P140 U87 ( .A1(n45), .A2(n82), .B1(n44), .B2(n32), .ZN(N305) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[17]), .ZN(n73) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[49]), .ZN(n33) );
  OAI22D1BWP30P140 U90 ( .A1(n45), .A2(n73), .B1(n44), .B2(n33), .ZN(N304) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[16]), .ZN(n72) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[48]), .ZN(n34) );
  OAI22D1BWP30P140 U93 ( .A1(n45), .A2(n72), .B1(n44), .B2(n34), .ZN(N303) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[15]), .ZN(n84) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[47]), .ZN(n35) );
  OAI22D1BWP30P140 U96 ( .A1(n45), .A2(n84), .B1(n44), .B2(n35), .ZN(N302) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[14]), .ZN(n83) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[46]), .ZN(n36) );
  OAI22D1BWP30P140 U99 ( .A1(n45), .A2(n83), .B1(n37), .B2(n36), .ZN(N301) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[13]), .ZN(n87) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[45]), .ZN(n38) );
  OAI22D1BWP30P140 U102 ( .A1(n45), .A2(n87), .B1(n44), .B2(n38), .ZN(N300) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[12]), .ZN(n88) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[44]), .ZN(n39) );
  OAI22D1BWP30P140 U105 ( .A1(n45), .A2(n88), .B1(n44), .B2(n39), .ZN(N299) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[11]), .ZN(n92) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[43]), .ZN(n40) );
  OAI22D1BWP30P140 U108 ( .A1(n45), .A2(n92), .B1(n44), .B2(n40), .ZN(N298) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[10]), .ZN(n89) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[42]), .ZN(n41) );
  OAI22D1BWP30P140 U111 ( .A1(n45), .A2(n89), .B1(n44), .B2(n41), .ZN(N297) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[8]), .ZN(n85) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[40]), .ZN(n42) );
  OAI22D1BWP30P140 U114 ( .A1(n45), .A2(n85), .B1(n44), .B2(n42), .ZN(N295) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[9]), .ZN(n86) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[41]), .ZN(n43) );
  OAI22D1BWP30P140 U117 ( .A1(n45), .A2(n86), .B1(n44), .B2(n43), .ZN(N296) );
  INVD1BWP30P140 U118 ( .I(n46), .ZN(n49) );
  INVD1BWP30P140 U119 ( .I(n50), .ZN(n47) );
  AN3D4BWP30P140 U120 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n47), .Z(n90) );
  OAI21D1BWP30P140 U121 ( .A1(n49), .A2(i_cmd[1]), .B(n48), .ZN(N354) );
  NR2D1BWP30P140 U122 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  MUX2NUD1BWP30P140 U123 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U124 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U125 ( .I(n55), .ZN(n71) );
  INVD1BWP30P140 U126 ( .I(n71), .ZN(n63) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  INVD2BWP30P140 U135 ( .I(n71), .ZN(n79) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n79), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n79), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n79), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n79), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n79), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n79), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  INVD2BWP30P140 U142 ( .I(n71), .ZN(n91) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n79), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n79), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n79), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n79), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n79), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n79), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_85 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD2BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n45), .A2(n19), .B1(n20), .B2(n83), .ZN(N306) );
  INVD3BWP30P140 U4 ( .I(n27), .ZN(n20) );
  INVD1BWP30P140 U5 ( .I(n5), .ZN(n27) );
  ND2OPTIBD1BWP30P140 U6 ( .A1(n47), .A2(n21), .ZN(n5) );
  OAI22D1BWP30P140 U7 ( .A1(n18), .A2(n17), .B1(n20), .B2(n84), .ZN(N307) );
  OAI22D1BWP30P140 U8 ( .A1(n18), .A2(n16), .B1(n20), .B2(n85), .ZN(N308) );
  OAI22D1BWP30P140 U9 ( .A1(n18), .A2(n15), .B1(n20), .B2(n86), .ZN(N309) );
  OAI22D1BWP30P140 U10 ( .A1(n18), .A2(n14), .B1(n20), .B2(n87), .ZN(N310) );
  OAI22D1BWP30P140 U11 ( .A1(n18), .A2(n13), .B1(n20), .B2(n88), .ZN(N311) );
  OAI22D1BWP30P140 U12 ( .A1(n18), .A2(n12), .B1(n20), .B2(n89), .ZN(N312) );
  OAI22D1BWP30P140 U13 ( .A1(n18), .A2(n11), .B1(n20), .B2(n90), .ZN(N313) );
  OAI22D1BWP30P140 U14 ( .A1(n18), .A2(n10), .B1(n20), .B2(n93), .ZN(N314) );
  OAI22D1BWP30P140 U15 ( .A1(n18), .A2(n9), .B1(n20), .B2(n80), .ZN(N315) );
  OAI22D1BWP30P140 U16 ( .A1(n18), .A2(n8), .B1(n20), .B2(n79), .ZN(N316) );
  OAI22D1BWP30P140 U17 ( .A1(n18), .A2(n7), .B1(n20), .B2(n67), .ZN(N317) );
  OAI22D1BWP30P140 U18 ( .A1(n18), .A2(n6), .B1(n20), .B2(n66), .ZN(N318) );
  ND2D1BWP30P140 U19 ( .A1(n1), .A2(i_en), .ZN(n51) );
  INVD1BWP30P140 U20 ( .I(n91), .ZN(n49) );
  INVD1BWP30P140 U21 ( .I(rst), .ZN(n1) );
  INVD1P5BWP30P140 U22 ( .I(i_cmd[0]), .ZN(n21) );
  NR2D1BWP30P140 U23 ( .A1(n51), .A2(n21), .ZN(n3) );
  INVD1BWP30P140 U24 ( .I(i_valid[0]), .ZN(n53) );
  INVD2BWP30P140 U25 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U26 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U27 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U28 ( .I(n4), .ZN(n22) );
  INVD2BWP30P140 U29 ( .I(n22), .ZN(n18) );
  INVD1BWP30P140 U30 ( .I(i_data_bus[63]), .ZN(n6) );
  INR2D1BWP30P140 U31 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  INVD1BWP30P140 U32 ( .I(i_data_bus[31]), .ZN(n66) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[62]), .ZN(n7) );
  INVD1BWP30P140 U34 ( .I(i_data_bus[30]), .ZN(n67) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[61]), .ZN(n8) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[29]), .ZN(n79) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[60]), .ZN(n9) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[28]), .ZN(n80) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[59]), .ZN(n10) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[27]), .ZN(n93) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[58]), .ZN(n11) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[26]), .ZN(n90) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[57]), .ZN(n12) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[25]), .ZN(n89) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[56]), .ZN(n13) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[24]), .ZN(n88) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[55]), .ZN(n14) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[23]), .ZN(n87) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[54]), .ZN(n15) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[22]), .ZN(n86) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[53]), .ZN(n16) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[21]), .ZN(n85) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[52]), .ZN(n17) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[20]), .ZN(n84) );
  INVD3BWP30P140 U55 ( .I(n22), .ZN(n45) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[51]), .ZN(n19) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[19]), .ZN(n83) );
  OAI31D1BWP30P140 U58 ( .A1(n51), .A2(n52), .A3(n21), .B(n20), .ZN(N353) );
  INVD2BWP30P140 U59 ( .I(n27), .ZN(n46) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD2BWP30P140 U61 ( .I(n22), .ZN(n38) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[39]), .ZN(n23) );
  OAI22D1BWP30P140 U63 ( .A1(n46), .A2(n57), .B1(n38), .B2(n23), .ZN(N294) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[38]), .ZN(n24) );
  OAI22D1BWP30P140 U66 ( .A1(n46), .A2(n58), .B1(n38), .B2(n24), .ZN(N293) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[37]), .ZN(n25) );
  OAI22D1BWP30P140 U69 ( .A1(n46), .A2(n59), .B1(n38), .B2(n25), .ZN(N292) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[36]), .ZN(n26) );
  OAI22D1BWP30P140 U72 ( .A1(n46), .A2(n60), .B1(n38), .B2(n26), .ZN(N291) );
  INVD1BWP30P140 U73 ( .I(n27), .ZN(n32) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[35]), .ZN(n28) );
  OAI22D1BWP30P140 U76 ( .A1(n32), .A2(n61), .B1(n38), .B2(n28), .ZN(N290) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[34]), .ZN(n29) );
  OAI22D1BWP30P140 U79 ( .A1(n32), .A2(n62), .B1(n38), .B2(n29), .ZN(N289) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[33]), .ZN(n30) );
  OAI22D1BWP30P140 U82 ( .A1(n32), .A2(n63), .B1(n38), .B2(n30), .ZN(N288) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[0]), .ZN(n65) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[32]), .ZN(n31) );
  OAI22D1BWP30P140 U85 ( .A1(n32), .A2(n65), .B1(n45), .B2(n31), .ZN(N287) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[18]), .ZN(n81) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[50]), .ZN(n33) );
  OAI22D1BWP30P140 U88 ( .A1(n46), .A2(n81), .B1(n45), .B2(n33), .ZN(N305) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[17]), .ZN(n78) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[49]), .ZN(n34) );
  OAI22D1BWP30P140 U91 ( .A1(n46), .A2(n78), .B1(n45), .B2(n34), .ZN(N304) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[16]), .ZN(n77) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[48]), .ZN(n35) );
  OAI22D1BWP30P140 U94 ( .A1(n46), .A2(n77), .B1(n45), .B2(n35), .ZN(N303) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[15]), .ZN(n76) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[47]), .ZN(n36) );
  OAI22D1BWP30P140 U97 ( .A1(n46), .A2(n76), .B1(n45), .B2(n36), .ZN(N302) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[14]), .ZN(n75) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[46]), .ZN(n37) );
  OAI22D1BWP30P140 U100 ( .A1(n46), .A2(n75), .B1(n38), .B2(n37), .ZN(N301) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[13]), .ZN(n74) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[45]), .ZN(n39) );
  OAI22D1BWP30P140 U103 ( .A1(n46), .A2(n74), .B1(n45), .B2(n39), .ZN(N300) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[12]), .ZN(n73) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[44]), .ZN(n40) );
  OAI22D1BWP30P140 U106 ( .A1(n46), .A2(n73), .B1(n45), .B2(n40), .ZN(N299) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[11]), .ZN(n72) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[43]), .ZN(n41) );
  OAI22D1BWP30P140 U109 ( .A1(n46), .A2(n72), .B1(n45), .B2(n41), .ZN(N298) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[10]), .ZN(n71) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[42]), .ZN(n42) );
  OAI22D1BWP30P140 U112 ( .A1(n46), .A2(n71), .B1(n45), .B2(n42), .ZN(N297) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[9]), .ZN(n70) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[41]), .ZN(n43) );
  OAI22D1BWP30P140 U115 ( .A1(n46), .A2(n70), .B1(n45), .B2(n43), .ZN(N296) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[8]), .ZN(n69) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[40]), .ZN(n44) );
  OAI22D1BWP30P140 U118 ( .A1(n46), .A2(n69), .B1(n45), .B2(n44), .ZN(N295) );
  INVD1BWP30P140 U119 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U120 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U121 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n91) );
  OAI21D1BWP30P140 U122 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  NR2D1BWP30P140 U123 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  MUX2NUD1BWP30P140 U124 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  ND2OPTIBD1BWP30P140 U125 ( .A1(n55), .A2(n54), .ZN(n56) );
  INVD2BWP30P140 U126 ( .I(n56), .ZN(n68) );
  INVD1BWP30P140 U127 ( .I(n68), .ZN(n64) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n64), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n64), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n64), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n64), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n64), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n64), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n64), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n64), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  INVD2BWP30P140 U136 ( .I(n68), .ZN(n92) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n92), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n92), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  INVD2BWP30P140 U139 ( .I(n68), .ZN(n82) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n82), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n82), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n82), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n82), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n82), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n82), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n82), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n82), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n82), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n82), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n92), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n92), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n82), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n82), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_86 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140 U3 ( .I(n29), .ZN(n25) );
  INVD2BWP30P140 U4 ( .I(n5), .ZN(n29) );
  ND2OPTIBD1BWP30P140 U5 ( .A1(n46), .A2(n26), .ZN(n5) );
  ND2D1BWP30P140 U6 ( .A1(n1), .A2(i_en), .ZN(n50) );
  INVD1BWP30P140 U7 ( .I(n90), .ZN(n48) );
  OAI22D1BWP30P140 U8 ( .A1(n44), .A2(n9), .B1(n45), .B2(n75), .ZN(N295) );
  OAI22D1BWP30P140 U9 ( .A1(n44), .A2(n8), .B1(n45), .B2(n74), .ZN(N296) );
  OAI22D1BWP30P140 U10 ( .A1(n44), .A2(n7), .B1(n45), .B2(n69), .ZN(N297) );
  OAI22D1BWP30P140 U11 ( .A1(n44), .A2(n6), .B1(n45), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U12 ( .A1(n44), .A2(n10), .B1(n45), .B2(n71), .ZN(N304) );
  OAI22D1BWP30P140 U13 ( .A1(n44), .A2(n22), .B1(n25), .B2(n73), .ZN(N306) );
  OAI22D1BWP30P140 U14 ( .A1(n24), .A2(n21), .B1(n25), .B2(n77), .ZN(N307) );
  OAI22D1BWP30P140 U15 ( .A1(n24), .A2(n20), .B1(n25), .B2(n78), .ZN(N308) );
  OAI22D1BWP30P140 U16 ( .A1(n24), .A2(n19), .B1(n25), .B2(n79), .ZN(N309) );
  OAI22D1BWP30P140 U17 ( .A1(n24), .A2(n18), .B1(n25), .B2(n80), .ZN(N310) );
  OAI22D1BWP30P140 U18 ( .A1(n24), .A2(n17), .B1(n25), .B2(n81), .ZN(N311) );
  OAI22D1BWP30P140 U19 ( .A1(n24), .A2(n14), .B1(n25), .B2(n82), .ZN(N312) );
  OAI22D1BWP30P140 U20 ( .A1(n24), .A2(n13), .B1(n25), .B2(n83), .ZN(N313) );
  OAI22D1BWP30P140 U21 ( .A1(n24), .A2(n12), .B1(n25), .B2(n84), .ZN(N314) );
  OAI22D1BWP30P140 U22 ( .A1(n24), .A2(n23), .B1(n25), .B2(n85), .ZN(N315) );
  OAI22D1BWP30P140 U23 ( .A1(n24), .A2(n16), .B1(n25), .B2(n86), .ZN(N316) );
  OAI22D1BWP30P140 U24 ( .A1(n24), .A2(n15), .B1(n25), .B2(n92), .ZN(N317) );
  OAI22D1BWP30P140 U25 ( .A1(n24), .A2(n11), .B1(n25), .B2(n87), .ZN(N318) );
  INVD1BWP30P140 U26 ( .I(rst), .ZN(n1) );
  INVD1P5BWP30P140 U27 ( .I(i_cmd[0]), .ZN(n26) );
  NR2D1BWP30P140 U28 ( .A1(n50), .A2(n26), .ZN(n3) );
  INVD1BWP30P140 U29 ( .I(i_valid[0]), .ZN(n52) );
  INVD2BWP30P140 U30 ( .I(i_valid[1]), .ZN(n51) );
  MUX2NUD1BWP30P140 U31 ( .I0(n52), .I1(n51), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U32 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U33 ( .I(n4), .ZN(n27) );
  INVD3BWP30P140 U34 ( .I(n27), .ZN(n44) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[43]), .ZN(n6) );
  INR2D2BWP30P140 U36 ( .A1(i_valid[0]), .B1(n50), .ZN(n46) );
  INVD2BWP30P140 U37 ( .I(n29), .ZN(n45) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[42]), .ZN(n7) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[10]), .ZN(n69) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[41]), .ZN(n8) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[9]), .ZN(n74) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n9) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[8]), .ZN(n75) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[49]), .ZN(n10) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[17]), .ZN(n71) );
  INVD2BWP30P140 U47 ( .I(n27), .ZN(n24) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[63]), .ZN(n11) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[31]), .ZN(n87) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[59]), .ZN(n12) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[27]), .ZN(n84) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[58]), .ZN(n13) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[26]), .ZN(n83) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[57]), .ZN(n14) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[25]), .ZN(n82) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[62]), .ZN(n15) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[30]), .ZN(n92) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[61]), .ZN(n16) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[29]), .ZN(n86) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[56]), .ZN(n17) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[24]), .ZN(n81) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[55]), .ZN(n18) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[23]), .ZN(n80) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[54]), .ZN(n19) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[22]), .ZN(n79) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[21]), .ZN(n78) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[52]), .ZN(n21) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[51]), .ZN(n22) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n73) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[60]), .ZN(n23) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[28]), .ZN(n85) );
  OAI31D1BWP30P140 U74 ( .A1(n50), .A2(n51), .A3(n26), .B(n25), .ZN(N353) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[7]), .ZN(n56) );
  INVD2BWP30P140 U76 ( .I(n27), .ZN(n42) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[39]), .ZN(n28) );
  OAI22D1BWP30P140 U78 ( .A1(n45), .A2(n56), .B1(n42), .B2(n28), .ZN(N294) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[32]), .ZN(n30) );
  OAI22D1BWP30P140 U81 ( .A1(n25), .A2(n64), .B1(n42), .B2(n30), .ZN(N287) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[1]), .ZN(n62) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[33]), .ZN(n31) );
  OAI22D1BWP30P140 U84 ( .A1(n25), .A2(n62), .B1(n42), .B2(n31), .ZN(N288) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[2]), .ZN(n61) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[34]), .ZN(n32) );
  OAI22D1BWP30P140 U87 ( .A1(n25), .A2(n61), .B1(n42), .B2(n32), .ZN(N289) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[5]), .ZN(n58) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[37]), .ZN(n33) );
  OAI22D1BWP30P140 U90 ( .A1(n45), .A2(n58), .B1(n42), .B2(n33), .ZN(N292) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[35]), .ZN(n34) );
  OAI22D1BWP30P140 U93 ( .A1(n25), .A2(n60), .B1(n44), .B2(n34), .ZN(N290) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[6]), .ZN(n57) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[38]), .ZN(n35) );
  OAI22D1BWP30P140 U96 ( .A1(n45), .A2(n57), .B1(n42), .B2(n35), .ZN(N293) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[36]), .ZN(n36) );
  OAI22D1BWP30P140 U99 ( .A1(n45), .A2(n59), .B1(n42), .B2(n36), .ZN(N291) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[18]), .ZN(n72) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[50]), .ZN(n37) );
  OAI22D1BWP30P140 U102 ( .A1(n45), .A2(n72), .B1(n44), .B2(n37), .ZN(N305) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[16]), .ZN(n70) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[48]), .ZN(n38) );
  OAI22D1BWP30P140 U105 ( .A1(n45), .A2(n70), .B1(n44), .B2(n38), .ZN(N303) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[15]), .ZN(n65) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[47]), .ZN(n39) );
  OAI22D1BWP30P140 U108 ( .A1(n45), .A2(n65), .B1(n44), .B2(n39), .ZN(N302) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[14]), .ZN(n89) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[46]), .ZN(n40) );
  OAI22D1BWP30P140 U111 ( .A1(n45), .A2(n89), .B1(n44), .B2(n40), .ZN(N301) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[13]), .ZN(n66) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[45]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n45), .A2(n66), .B1(n42), .B2(n41), .ZN(N300) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[12]), .ZN(n67) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[44]), .ZN(n43) );
  OAI22D1BWP30P140 U117 ( .A1(n45), .A2(n67), .B1(n44), .B2(n43), .ZN(N299) );
  INVD1BWP30P140 U118 ( .I(n46), .ZN(n49) );
  INVD1BWP30P140 U119 ( .I(n50), .ZN(n47) );
  AN3D4BWP30P140 U120 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n47), .Z(n90) );
  OAI21D1BWP30P140 U121 ( .A1(n49), .A2(i_cmd[1]), .B(n48), .ZN(N354) );
  NR2D1BWP30P140 U122 ( .A1(n50), .A2(i_cmd[1]), .ZN(n54) );
  MUX2NUD1BWP30P140 U123 ( .I0(n52), .I1(n51), .S(i_cmd[0]), .ZN(n53) );
  ND2OPTIBD1BWP30P140 U124 ( .A1(n54), .A2(n53), .ZN(n55) );
  INVD2BWP30P140 U125 ( .I(n55), .ZN(n76) );
  INVD1BWP30P140 U126 ( .I(n76), .ZN(n63) );
  MOAI22D1BWP30P140 U127 ( .A1(n56), .A2(n63), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n63), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n63), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n63), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n63), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n63), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n63), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n63), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  INVD2BWP30P140 U135 ( .I(n76), .ZN(n88) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n88), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n88), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n88), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n88), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n88), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n88), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n88), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n88), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n88), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n88), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n88), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  INVD2BWP30P140 U147 ( .I(n76), .ZN(n91) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U156 ( .A1(n85), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U157 ( .A1(n86), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U158 ( .A1(n87), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n88), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_87 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  OAI22D1BWP30P140 U3 ( .A1(n33), .A2(n25), .B1(n1), .B2(n86), .ZN(N314) );
  OAI22D1BWP30P140 U4 ( .A1(n35), .A2(n14), .B1(n47), .B2(n74), .ZN(N300) );
  OAI22D1BWP30P140 U5 ( .A1(n33), .A2(n26), .B1(n1), .B2(n87), .ZN(N313) );
  OAI22D1BWP30P140 U6 ( .A1(n35), .A2(n19), .B1(n47), .B2(n78), .ZN(N296) );
  OAI22D1BWP30P140 U7 ( .A1(n33), .A2(n29), .B1(n1), .B2(n90), .ZN(N310) );
  OAI22D1BWP30P140 U8 ( .A1(n33), .A2(n24), .B1(n2), .B2(n85), .ZN(N315) );
  OAI22D1BWP30P140 U9 ( .A1(n33), .A2(n23), .B1(n47), .B2(n84), .ZN(N316) );
  OAI22D1BWP30P140 U10 ( .A1(n33), .A2(n30), .B1(n1), .B2(n93), .ZN(N309) );
  OAI22D1BWP30P140 U11 ( .A1(n33), .A2(n28), .B1(n2), .B2(n89), .ZN(N311) );
  OAI22D1BWP30P140 U12 ( .A1(n33), .A2(n27), .B1(n47), .B2(n88), .ZN(N312) );
  OAI22D1BWP30P140 U13 ( .A1(n35), .A2(n34), .B1(n1), .B2(n68), .ZN(N306) );
  OAI22D1BWP30P140 U14 ( .A1(n33), .A2(n32), .B1(n2), .B2(n66), .ZN(N307) );
  OAI22D1BWP30P140 U15 ( .A1(n33), .A2(n31), .B1(n47), .B2(n81), .ZN(N308) );
  OAI22D1BWP30P140 U16 ( .A1(n35), .A2(n20), .B1(n2), .B2(n80), .ZN(N295) );
  OAI22D1BWP30P140 U17 ( .A1(n35), .A2(n10), .B1(n2), .B2(n70), .ZN(N304) );
  INVD4BWP30P140 U18 ( .I(n15), .ZN(n1) );
  INVD3BWP30P140 U19 ( .I(n15), .ZN(n2) );
  INVD2BWP30P140 U20 ( .I(n8), .ZN(n15) );
  ND2OPTIBD1BWP30P140 U21 ( .A1(n48), .A2(n36), .ZN(n8) );
  INVD1BWP30P140 U22 ( .I(n57), .ZN(n67) );
  ND2D1BWP30P140 U23 ( .A1(n4), .A2(i_en), .ZN(n52) );
  CKBD1BWP30P140 U24 ( .I(n57), .Z(n3) );
  INVD1BWP30P140 U25 ( .I(n91), .ZN(n50) );
  CKND2D2BWP30P140 U26 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U27 ( .I(rst), .ZN(n4) );
  INVD1P5BWP30P140 U28 ( .I(i_cmd[0]), .ZN(n36) );
  NR2D1BWP30P140 U29 ( .A1(n52), .A2(n36), .ZN(n6) );
  INVD1BWP30P140 U30 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U31 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U32 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n5) );
  ND2OPTIBD1BWP30P140 U33 ( .A1(n6), .A2(n5), .ZN(n7) );
  INVD2BWP30P140 U34 ( .I(n7), .ZN(n37) );
  INVD2BWP30P140 U35 ( .I(n37), .ZN(n35) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[50]), .ZN(n9) );
  INR2D2BWP30P140 U37 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[18]), .ZN(n69) );
  OAI22OPTPBD1BWP30P140 U39 ( .A1(n35), .A2(n9), .B1(n2), .B2(n69), .ZN(N305)
         );
  INVD1BWP30P140 U40 ( .I(i_data_bus[49]), .ZN(n10) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[17]), .ZN(n70) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[48]), .ZN(n11) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[16]), .ZN(n71) );
  OAI22OPTPBD1BWP30P140 U44 ( .A1(n35), .A2(n11), .B1(n2), .B2(n71), .ZN(N303)
         );
  INVD1BWP30P140 U45 ( .I(i_data_bus[47]), .ZN(n12) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[15]), .ZN(n72) );
  OAI22OPTPBD1BWP30P140 U47 ( .A1(n35), .A2(n12), .B1(n1), .B2(n72), .ZN(N302)
         );
  INVD1BWP30P140 U48 ( .I(i_data_bus[46]), .ZN(n13) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[14]), .ZN(n73) );
  OAI22OPTPBD1BWP30P140 U50 ( .A1(n35), .A2(n13), .B1(n1), .B2(n73), .ZN(N301)
         );
  INVD1BWP30P140 U51 ( .I(i_data_bus[45]), .ZN(n14) );
  INVD2BWP30P140 U52 ( .I(n15), .ZN(n47) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[13]), .ZN(n74) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n16) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n75) );
  OAI22OPTPBD1BWP30P140 U56 ( .A1(n35), .A2(n16), .B1(n2), .B2(n75), .ZN(N299)
         );
  INVD1BWP30P140 U57 ( .I(i_data_bus[43]), .ZN(n17) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[11]), .ZN(n76) );
  OAI22OPTPBD1BWP30P140 U59 ( .A1(n35), .A2(n17), .B1(n1), .B2(n76), .ZN(N298)
         );
  INVD1BWP30P140 U60 ( .I(i_data_bus[42]), .ZN(n18) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[10]), .ZN(n77) );
  OAI22OPTPBD1BWP30P140 U62 ( .A1(n35), .A2(n18), .B1(n1), .B2(n77), .ZN(N297)
         );
  INVD1BWP30P140 U63 ( .I(i_data_bus[41]), .ZN(n19) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[9]), .ZN(n78) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[40]), .ZN(n20) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[8]), .ZN(n80) );
  INVD2BWP30P140 U67 ( .I(n37), .ZN(n33) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[63]), .ZN(n21) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[31]), .ZN(n82) );
  OAI22OPTPBD1BWP30P140 U70 ( .A1(n33), .A2(n21), .B1(n1), .B2(n82), .ZN(N318)
         );
  INVD1BWP30P140 U71 ( .I(i_data_bus[62]), .ZN(n22) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[30]), .ZN(n83) );
  OAI22OPTPBD1BWP30P140 U73 ( .A1(n33), .A2(n22), .B1(n1), .B2(n83), .ZN(N317)
         );
  INVD1BWP30P140 U74 ( .I(i_data_bus[61]), .ZN(n23) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[29]), .ZN(n84) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[60]), .ZN(n24) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[28]), .ZN(n85) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[59]), .ZN(n25) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[27]), .ZN(n86) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[58]), .ZN(n26) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[26]), .ZN(n87) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[57]), .ZN(n27) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[25]), .ZN(n88) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[56]), .ZN(n28) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[24]), .ZN(n89) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[55]), .ZN(n29) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[23]), .ZN(n90) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[54]), .ZN(n30) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[22]), .ZN(n93) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[53]), .ZN(n31) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[21]), .ZN(n81) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[52]), .ZN(n32) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[20]), .ZN(n66) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[51]), .ZN(n34) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[19]), .ZN(n68) );
  OAI31D1BWP30P140 U96 ( .A1(n52), .A2(n53), .A3(n36), .B(n47), .ZN(N353) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[5]), .ZN(n63) );
  INVD2BWP30P140 U98 ( .I(n37), .ZN(n46) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U100 ( .A1(n1), .A2(n63), .B1(n46), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[6]), .ZN(n64) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[38]), .ZN(n39) );
  OAI22D1BWP30P140 U103 ( .A1(n2), .A2(n64), .B1(n46), .B2(n39), .ZN(N293) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[7]), .ZN(n65) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[39]), .ZN(n40) );
  OAI22D1BWP30P140 U106 ( .A1(n1), .A2(n65), .B1(n46), .B2(n40), .ZN(N294) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[36]), .ZN(n41) );
  OAI22D1BWP30P140 U109 ( .A1(n1), .A2(n62), .B1(n46), .B2(n41), .ZN(N291) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[35]), .ZN(n42) );
  OAI22D1BWP30P140 U112 ( .A1(n2), .A2(n61), .B1(n46), .B2(n42), .ZN(N290) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[34]), .ZN(n43) );
  OAI22D1BWP30P140 U115 ( .A1(n1), .A2(n60), .B1(n46), .B2(n43), .ZN(N289) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[33]), .ZN(n44) );
  OAI22D1BWP30P140 U118 ( .A1(n1), .A2(n59), .B1(n46), .B2(n44), .ZN(N288) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[0]), .ZN(n58) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[32]), .ZN(n45) );
  OAI22D1BWP30P140 U121 ( .A1(n47), .A2(n58), .B1(n46), .B2(n45), .ZN(N287) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n3), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n3), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n3), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n3), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n3), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n3), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n3), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n3), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  INVD2BWP30P140 U136 ( .I(n67), .ZN(n92) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n92), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  INVD2BWP30P140 U138 ( .I(n67), .ZN(n79) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n79), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n79), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n79), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n79), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n79), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n79), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n79), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n79), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n79), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n79), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n79), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n79), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_88 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD2BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  OAI22D1BWP30P140 U3 ( .A1(n33), .A2(n22), .B1(n1), .B2(n69), .ZN(N317) );
  OAI22D1BWP30P140 U4 ( .A1(n35), .A2(n14), .B1(n47), .B2(n90), .ZN(N302) );
  OAI22D1BWP30P140 U5 ( .A1(n33), .A2(n25), .B1(n1), .B2(n72), .ZN(N314) );
  OAI22D1BWP30P140 U6 ( .A1(n35), .A2(n19), .B1(n47), .B2(n78), .ZN(N298) );
  OAI22D1BWP30P140 U7 ( .A1(n33), .A2(n26), .B1(n1), .B2(n73), .ZN(N313) );
  OAI22D1BWP30P140 U8 ( .A1(n33), .A2(n24), .B1(n2), .B2(n71), .ZN(N315) );
  OAI22D1BWP30P140 U9 ( .A1(n33), .A2(n23), .B1(n47), .B2(n68), .ZN(N318) );
  OAI22D1BWP30P140 U10 ( .A1(n33), .A2(n30), .B1(n1), .B2(n82), .ZN(N309) );
  OAI22D1BWP30P140 U11 ( .A1(n33), .A2(n28), .B1(n2), .B2(n75), .ZN(N311) );
  OAI22D1BWP30P140 U12 ( .A1(n33), .A2(n27), .B1(n47), .B2(n74), .ZN(N312) );
  OAI22D1BWP30P140 U13 ( .A1(n35), .A2(n34), .B1(n1), .B2(n86), .ZN(N306) );
  OAI22D1BWP30P140 U14 ( .A1(n33), .A2(n32), .B1(n2), .B2(n85), .ZN(N307) );
  OAI22D1BWP30P140 U15 ( .A1(n33), .A2(n31), .B1(n47), .B2(n83), .ZN(N308) );
  OAI22D1BWP30P140 U16 ( .A1(n35), .A2(n9), .B1(n2), .B2(n66), .ZN(N295) );
  OAI22D1BWP30P140 U17 ( .A1(n33), .A2(n29), .B1(n1), .B2(n81), .ZN(N310) );
  INVD4BWP30P140 U18 ( .I(n15), .ZN(n1) );
  INVD3BWP30P140 U19 ( .I(n15), .ZN(n2) );
  INVD2BWP30P140 U20 ( .I(n8), .ZN(n15) );
  ND2OPTIBD1BWP30P140 U21 ( .A1(n48), .A2(n36), .ZN(n8) );
  INVD1BWP30P140 U22 ( .I(n57), .ZN(n67) );
  ND2D1BWP30P140 U23 ( .A1(n4), .A2(i_en), .ZN(n52) );
  CKBD1BWP30P140 U24 ( .I(n57), .Z(n3) );
  INVD1BWP30P140 U25 ( .I(n91), .ZN(n50) );
  CKND2D2BWP30P140 U26 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U27 ( .I(rst), .ZN(n4) );
  INVD1P5BWP30P140 U28 ( .I(i_cmd[0]), .ZN(n36) );
  NR2D1BWP30P140 U29 ( .A1(n52), .A2(n36), .ZN(n6) );
  INVD1BWP30P140 U30 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U31 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U32 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n5) );
  ND2OPTIBD1BWP30P140 U33 ( .A1(n6), .A2(n5), .ZN(n7) );
  INVD2BWP30P140 U34 ( .I(n7), .ZN(n37) );
  INVD2BWP30P140 U35 ( .I(n37), .ZN(n35) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[40]), .ZN(n9) );
  INR2D2BWP30P140 U37 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  INVD1BWP30P140 U38 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[50]), .ZN(n10) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[18]), .ZN(n87) );
  OAI22OPTPBD1BWP30P140 U41 ( .A1(n35), .A2(n10), .B1(n2), .B2(n87), .ZN(N305)
         );
  INVD1BWP30P140 U42 ( .I(i_data_bus[49]), .ZN(n11) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[17]), .ZN(n88) );
  OAI22OPTPBD1BWP30P140 U44 ( .A1(n35), .A2(n11), .B1(n2), .B2(n88), .ZN(N304)
         );
  INVD1BWP30P140 U45 ( .I(i_data_bus[48]), .ZN(n12) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[16]), .ZN(n89) );
  OAI22OPTPBD1BWP30P140 U47 ( .A1(n35), .A2(n12), .B1(n1), .B2(n89), .ZN(N303)
         );
  INVD1BWP30P140 U48 ( .I(i_data_bus[41]), .ZN(n13) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[9]), .ZN(n76) );
  OAI22OPTPBD1BWP30P140 U50 ( .A1(n35), .A2(n13), .B1(n1), .B2(n76), .ZN(N296)
         );
  INVD1BWP30P140 U51 ( .I(i_data_bus[47]), .ZN(n14) );
  INVD2BWP30P140 U52 ( .I(n15), .ZN(n47) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[15]), .ZN(n90) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[46]), .ZN(n16) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[14]), .ZN(n93) );
  OAI22OPTPBD1BWP30P140 U56 ( .A1(n35), .A2(n16), .B1(n2), .B2(n93), .ZN(N301)
         );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n17) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n80) );
  OAI22OPTPBD1BWP30P140 U59 ( .A1(n35), .A2(n17), .B1(n1), .B2(n80), .ZN(N300)
         );
  INVD1BWP30P140 U60 ( .I(i_data_bus[44]), .ZN(n18) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[12]), .ZN(n79) );
  OAI22OPTPBD1BWP30P140 U62 ( .A1(n35), .A2(n18), .B1(n1), .B2(n79), .ZN(N299)
         );
  INVD1BWP30P140 U63 ( .I(i_data_bus[43]), .ZN(n19) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[11]), .ZN(n78) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[42]), .ZN(n20) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[10]), .ZN(n77) );
  OAI22OPTPBD1BWP30P140 U67 ( .A1(n35), .A2(n20), .B1(n2), .B2(n77), .ZN(N297)
         );
  INVD2BWP30P140 U68 ( .I(n37), .ZN(n33) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[61]), .ZN(n21) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[29]), .ZN(n70) );
  OAI22OPTPBD1BWP30P140 U71 ( .A1(n33), .A2(n21), .B1(n1), .B2(n70), .ZN(N316)
         );
  INVD1BWP30P140 U72 ( .I(i_data_bus[62]), .ZN(n22) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[30]), .ZN(n69) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[63]), .ZN(n23) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[31]), .ZN(n68) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[60]), .ZN(n24) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[28]), .ZN(n71) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[59]), .ZN(n25) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[27]), .ZN(n72) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[58]), .ZN(n26) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[26]), .ZN(n73) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[57]), .ZN(n27) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[25]), .ZN(n74) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[56]), .ZN(n28) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[24]), .ZN(n75) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[55]), .ZN(n29) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[23]), .ZN(n81) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[54]), .ZN(n30) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[22]), .ZN(n82) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[53]), .ZN(n31) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[21]), .ZN(n83) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[52]), .ZN(n32) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[20]), .ZN(n85) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[51]), .ZN(n34) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[19]), .ZN(n86) );
  OAI31D1BWP30P140 U96 ( .A1(n52), .A2(n53), .A3(n36), .B(n47), .ZN(N353) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[5]), .ZN(n63) );
  INVD2BWP30P140 U98 ( .I(n37), .ZN(n46) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U100 ( .A1(n1), .A2(n63), .B1(n46), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[7]), .ZN(n65) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[39]), .ZN(n39) );
  OAI22D1BWP30P140 U103 ( .A1(n2), .A2(n65), .B1(n46), .B2(n39), .ZN(N294) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[36]), .ZN(n40) );
  OAI22D1BWP30P140 U106 ( .A1(n1), .A2(n62), .B1(n46), .B2(n40), .ZN(N291) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[6]), .ZN(n64) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[38]), .ZN(n41) );
  OAI22D1BWP30P140 U109 ( .A1(n1), .A2(n64), .B1(n46), .B2(n41), .ZN(N293) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[33]), .ZN(n42) );
  OAI22D1BWP30P140 U112 ( .A1(n2), .A2(n59), .B1(n46), .B2(n42), .ZN(N288) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[0]), .ZN(n58) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[32]), .ZN(n43) );
  OAI22D1BWP30P140 U115 ( .A1(n1), .A2(n58), .B1(n46), .B2(n43), .ZN(N287) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[35]), .ZN(n44) );
  OAI22D1BWP30P140 U118 ( .A1(n1), .A2(n61), .B1(n46), .B2(n44), .ZN(N290) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[34]), .ZN(n45) );
  OAI22D1BWP30P140 U121 ( .A1(n47), .A2(n60), .B1(n46), .B2(n45), .ZN(N289) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n3), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n3), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n3), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n3), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n3), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n3), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n3), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n3), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  INVD2BWP30P140 U136 ( .I(n67), .ZN(n92) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n92), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  INVD2BWP30P140 U138 ( .I(n67), .ZN(n84) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n84), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n84), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n84), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n84), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n84), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n84), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n84), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n84), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n92), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n92), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n92), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n92), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n92), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n84), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n84), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n84), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n84), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_89 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n33), .A2(n25), .B1(n1), .B2(n76), .ZN(N314) );
  OAI22D1BWP30P140 U4 ( .A1(n35), .A2(n20), .B1(n2), .B2(n89), .ZN(N305) );
  OAI22D1BWP30P140 U5 ( .A1(n33), .A2(n26), .B1(n1), .B2(n77), .ZN(N315) );
  OAI22D1BWP30P140 U6 ( .A1(n35), .A2(n14), .B1(n42), .B2(n72), .ZN(N296) );
  OAI22D1BWP30P140 U7 ( .A1(n33), .A2(n29), .B1(n1), .B2(n80), .ZN(N318) );
  OAI22D1BWP30P140 U8 ( .A1(n35), .A2(n19), .B1(n42), .B2(n66), .ZN(N302) );
  OAI22D1BWP30P140 U9 ( .A1(n33), .A2(n24), .B1(n2), .B2(n75), .ZN(N313) );
  OAI22D1BWP30P140 U10 ( .A1(n33), .A2(n30), .B1(n1), .B2(n84), .ZN(N309) );
  OAI22D1BWP30P140 U11 ( .A1(n33), .A2(n28), .B1(n2), .B2(n79), .ZN(N317) );
  OAI22D1BWP30P140 U12 ( .A1(n33), .A2(n23), .B1(n42), .B2(n81), .ZN(N312) );
  OAI22D1BWP30P140 U13 ( .A1(n35), .A2(n34), .B1(n1), .B2(n88), .ZN(N306) );
  OAI22D1BWP30P140 U14 ( .A1(n33), .A2(n32), .B1(n2), .B2(n87), .ZN(N307) );
  OAI22D1BWP30P140 U15 ( .A1(n33), .A2(n31), .B1(n42), .B2(n85), .ZN(N308) );
  OAI22D1BWP30P140 U16 ( .A1(n35), .A2(n16), .B1(n2), .B2(n73), .ZN(N295) );
  OAI22D1BWP30P140 U17 ( .A1(n35), .A2(n9), .B1(n2), .B2(n67), .ZN(N301) );
  OAI22D1BWP30P140 U18 ( .A1(n33), .A2(n27), .B1(n42), .B2(n78), .ZN(N316) );
  INVD4BWP30P140 U19 ( .I(n15), .ZN(n1) );
  INVD3BWP30P140 U20 ( .I(n15), .ZN(n2) );
  INVD2BWP30P140 U21 ( .I(n8), .ZN(n15) );
  ND2OPTIBD1BWP30P140 U22 ( .A1(n48), .A2(n36), .ZN(n8) );
  INVD1BWP30P140 U23 ( .I(n57), .ZN(n74) );
  ND2D1BWP30P140 U24 ( .A1(n4), .A2(i_en), .ZN(n52) );
  CKBD1BWP30P140 U25 ( .I(n57), .Z(n3) );
  INVD1BWP30P140 U26 ( .I(n91), .ZN(n50) );
  CKND2D2BWP30P140 U27 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U28 ( .I(rst), .ZN(n4) );
  INVD1P5BWP30P140 U29 ( .I(i_cmd[0]), .ZN(n36) );
  NR2D1BWP30P140 U30 ( .A1(n52), .A2(n36), .ZN(n6) );
  INVD1BWP30P140 U31 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U32 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U33 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n5) );
  ND2OPTIBD1BWP30P140 U34 ( .A1(n6), .A2(n5), .ZN(n7) );
  INVD2BWP30P140 U35 ( .I(n7), .ZN(n37) );
  INVD2BWP30P140 U36 ( .I(n37), .ZN(n35) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[46]), .ZN(n9) );
  INR2D2BWP30P140 U38 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[14]), .ZN(n67) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[45]), .ZN(n10) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[13]), .ZN(n68) );
  OAI22OPTPBD1BWP30P140 U42 ( .A1(n35), .A2(n10), .B1(n2), .B2(n68), .ZN(N300)
         );
  INVD1BWP30P140 U43 ( .I(i_data_bus[44]), .ZN(n11) );
  INVD1BWP30P140 U44 ( .I(i_data_bus[12]), .ZN(n69) );
  OAI22OPTPBD1BWP30P140 U45 ( .A1(n35), .A2(n11), .B1(n2), .B2(n69), .ZN(N299)
         );
  INVD1BWP30P140 U46 ( .I(i_data_bus[43]), .ZN(n12) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[11]), .ZN(n70) );
  OAI22OPTPBD1BWP30P140 U48 ( .A1(n35), .A2(n12), .B1(n1), .B2(n70), .ZN(N298)
         );
  INVD1BWP30P140 U49 ( .I(i_data_bus[42]), .ZN(n13) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[10]), .ZN(n71) );
  OAI22OPTPBD1BWP30P140 U51 ( .A1(n35), .A2(n13), .B1(n1), .B2(n71), .ZN(N297)
         );
  INVD1BWP30P140 U52 ( .I(i_data_bus[41]), .ZN(n14) );
  INVD2BWP30P140 U53 ( .I(n15), .ZN(n42) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[9]), .ZN(n72) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[40]), .ZN(n16) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[8]), .ZN(n73) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[48]), .ZN(n17) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[16]), .ZN(n93) );
  OAI22OPTPBD1BWP30P140 U59 ( .A1(n35), .A2(n17), .B1(n1), .B2(n93), .ZN(N303)
         );
  INVD1BWP30P140 U60 ( .I(i_data_bus[49]), .ZN(n18) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[17]), .ZN(n90) );
  OAI22OPTPBD1BWP30P140 U62 ( .A1(n35), .A2(n18), .B1(n1), .B2(n90), .ZN(N304)
         );
  INVD1BWP30P140 U63 ( .I(i_data_bus[47]), .ZN(n19) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[15]), .ZN(n66) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[50]), .ZN(n20) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[18]), .ZN(n89) );
  INVD2BWP30P140 U67 ( .I(n37), .ZN(n33) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[55]), .ZN(n21) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[23]), .ZN(n83) );
  OAI22OPTPBD1BWP30P140 U70 ( .A1(n33), .A2(n21), .B1(n1), .B2(n83), .ZN(N310)
         );
  INVD1BWP30P140 U71 ( .I(i_data_bus[56]), .ZN(n22) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[24]), .ZN(n82) );
  OAI22OPTPBD1BWP30P140 U73 ( .A1(n33), .A2(n22), .B1(n1), .B2(n82), .ZN(N311)
         );
  INVD1BWP30P140 U74 ( .I(i_data_bus[57]), .ZN(n23) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[25]), .ZN(n81) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[58]), .ZN(n24) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[26]), .ZN(n75) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[59]), .ZN(n25) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[27]), .ZN(n76) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[60]), .ZN(n26) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[28]), .ZN(n77) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[61]), .ZN(n27) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[29]), .ZN(n78) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[62]), .ZN(n28) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[30]), .ZN(n79) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[63]), .ZN(n29) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[31]), .ZN(n80) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[54]), .ZN(n30) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[22]), .ZN(n84) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[53]), .ZN(n31) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[21]), .ZN(n85) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[52]), .ZN(n32) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[20]), .ZN(n87) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[51]), .ZN(n34) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[19]), .ZN(n88) );
  OAI31D1BWP30P140 U96 ( .A1(n52), .A2(n53), .A3(n36), .B(n42), .ZN(N353) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[1]), .ZN(n64) );
  INVD2BWP30P140 U98 ( .I(n37), .ZN(n47) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[33]), .ZN(n38) );
  OAI22D1BWP30P140 U100 ( .A1(n2), .A2(n64), .B1(n47), .B2(n38), .ZN(N288) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[2]), .ZN(n63) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[34]), .ZN(n39) );
  OAI22D1BWP30P140 U103 ( .A1(n1), .A2(n63), .B1(n47), .B2(n39), .ZN(N289) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[3]), .ZN(n62) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[35]), .ZN(n40) );
  OAI22D1BWP30P140 U106 ( .A1(n1), .A2(n62), .B1(n47), .B2(n40), .ZN(N290) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[0]), .ZN(n65) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[32]), .ZN(n41) );
  OAI22D1BWP30P140 U109 ( .A1(n42), .A2(n65), .B1(n47), .B2(n41), .ZN(N287) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[5]), .ZN(n60) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[37]), .ZN(n43) );
  OAI22D1BWP30P140 U112 ( .A1(n1), .A2(n60), .B1(n47), .B2(n43), .ZN(N292) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[6]), .ZN(n59) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[38]), .ZN(n44) );
  OAI22D1BWP30P140 U115 ( .A1(n2), .A2(n59), .B1(n47), .B2(n44), .ZN(N293) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[7]), .ZN(n58) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[39]), .ZN(n45) );
  OAI22D1BWP30P140 U118 ( .A1(n1), .A2(n58), .B1(n47), .B2(n45), .ZN(N294) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[36]), .ZN(n46) );
  OAI22D1BWP30P140 U121 ( .A1(n1), .A2(n61), .B1(n47), .B2(n46), .ZN(N291) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n3), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n3), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n3), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n3), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n3), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n3), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n3), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n3), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  INVD2BWP30P140 U136 ( .I(n74), .ZN(n92) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n92), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n92), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n92), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n92), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n92), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n92), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n92), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n92), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  INVD2BWP30P140 U145 ( .I(n74), .ZN(n86) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n86), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n86), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n86), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n86), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n86), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n86), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n86), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n86), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n86), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n86), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U156 ( .A1(n85), .A2(n86), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n86), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_90 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n19), .A2(n18), .B1(n31), .B2(n78), .ZN(N306) );
  INVD1BWP30P140 U4 ( .I(n57), .ZN(n79) );
  ND2D1BWP30P140 U5 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U6 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U7 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U8 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U9 ( .A1(n19), .A2(n7), .B1(n47), .B2(n66), .ZN(N295) );
  OAI22D1BWP30P140 U10 ( .A1(n19), .A2(n8), .B1(n47), .B2(n67), .ZN(N296) );
  OAI22D1BWP30P140 U11 ( .A1(n19), .A2(n9), .B1(n47), .B2(n68), .ZN(N297) );
  OAI22D1BWP30P140 U12 ( .A1(n19), .A2(n10), .B1(n47), .B2(n69), .ZN(N298) );
  OAI22D1BWP30P140 U13 ( .A1(n19), .A2(n11), .B1(n47), .B2(n70), .ZN(N299) );
  OAI22D1BWP30P140 U14 ( .A1(n19), .A2(n12), .B1(n47), .B2(n71), .ZN(N300) );
  OAI22D1BWP30P140 U15 ( .A1(n19), .A2(n13), .B1(n47), .B2(n72), .ZN(N301) );
  OAI22D1BWP30P140 U16 ( .A1(n19), .A2(n14), .B1(n47), .B2(n73), .ZN(N302) );
  OAI22D1BWP30P140 U17 ( .A1(n19), .A2(n15), .B1(n47), .B2(n74), .ZN(N303) );
  OAI22D1BWP30P140 U18 ( .A1(n19), .A2(n16), .B1(n47), .B2(n75), .ZN(N304) );
  OAI22D1BWP30P140 U19 ( .A1(n19), .A2(n17), .B1(n47), .B2(n76), .ZN(N305) );
  OAI22D1BWP30P140 U20 ( .A1(n33), .A2(n20), .B1(n31), .B2(n80), .ZN(N307) );
  OAI22D1BWP30P140 U21 ( .A1(n33), .A2(n21), .B1(n31), .B2(n81), .ZN(N308) );
  OAI22D1BWP30P140 U22 ( .A1(n33), .A2(n22), .B1(n31), .B2(n82), .ZN(N309) );
  OAI22D1BWP30P140 U23 ( .A1(n33), .A2(n23), .B1(n31), .B2(n83), .ZN(N310) );
  OAI22D1BWP30P140 U24 ( .A1(n33), .A2(n24), .B1(n31), .B2(n84), .ZN(N311) );
  OAI22D1BWP30P140 U25 ( .A1(n33), .A2(n25), .B1(n31), .B2(n85), .ZN(N312) );
  OAI22D1BWP30P140 U26 ( .A1(n33), .A2(n26), .B1(n31), .B2(n86), .ZN(N313) );
  OAI22D1BWP30P140 U27 ( .A1(n33), .A2(n27), .B1(n31), .B2(n87), .ZN(N314) );
  OAI22D1BWP30P140 U28 ( .A1(n33), .A2(n28), .B1(n31), .B2(n88), .ZN(N315) );
  OAI22D1BWP30P140 U29 ( .A1(n33), .A2(n29), .B1(n31), .B2(n89), .ZN(N316) );
  OAI22D1BWP30P140 U30 ( .A1(n33), .A2(n30), .B1(n31), .B2(n90), .ZN(N317) );
  OAI22D1BWP30P140 U31 ( .A1(n33), .A2(n32), .B1(n31), .B2(n93), .ZN(N318) );
  CKND2D2BWP30P140 U32 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U34 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U35 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U36 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U37 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U38 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U39 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U40 ( .I(n36), .ZN(n19) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[40]), .ZN(n7) );
  INR2D1BWP30P140 U42 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U43 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U44 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U45 ( .I(n34), .ZN(n47) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[41]), .ZN(n8) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[9]), .ZN(n67) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[42]), .ZN(n9) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[10]), .ZN(n68) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[43]), .ZN(n10) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[44]), .ZN(n11) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[12]), .ZN(n70) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[13]), .ZN(n71) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[46]), .ZN(n13) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[14]), .ZN(n72) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[47]), .ZN(n14) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[15]), .ZN(n73) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[48]), .ZN(n15) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[16]), .ZN(n74) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[49]), .ZN(n16) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[17]), .ZN(n75) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[50]), .ZN(n17) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[18]), .ZN(n76) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[51]), .ZN(n18) );
  INVD2BWP30P140 U68 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD2BWP30P140 U70 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[52]), .ZN(n20) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[53]), .ZN(n21) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[21]), .ZN(n81) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[54]), .ZN(n22) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[22]), .ZN(n82) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[55]), .ZN(n23) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[23]), .ZN(n83) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[56]), .ZN(n24) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[24]), .ZN(n84) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[57]), .ZN(n25) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[25]), .ZN(n85) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[58]), .ZN(n26) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[26]), .ZN(n86) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[59]), .ZN(n27) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[27]), .ZN(n87) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[60]), .ZN(n28) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[28]), .ZN(n88) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[61]), .ZN(n29) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[29]), .ZN(n89) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[62]), .ZN(n30) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[30]), .ZN(n90) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[63]), .ZN(n32) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[31]), .ZN(n93) );
  INVD1BWP30P140 U95 ( .I(n34), .ZN(n41) );
  OAI31D1BWP30P140 U96 ( .A1(n52), .A2(n53), .A3(n35), .B(n41), .ZN(N353) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[0]), .ZN(n65) );
  INVD2BWP30P140 U98 ( .I(n36), .ZN(n46) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[32]), .ZN(n37) );
  OAI22D1BWP30P140 U100 ( .A1(n41), .A2(n65), .B1(n46), .B2(n37), .ZN(N287) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[1]), .ZN(n64) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[33]), .ZN(n38) );
  OAI22D1BWP30P140 U103 ( .A1(n41), .A2(n64), .B1(n46), .B2(n38), .ZN(N288) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[2]), .ZN(n63) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[34]), .ZN(n39) );
  OAI22D1BWP30P140 U106 ( .A1(n41), .A2(n63), .B1(n46), .B2(n39), .ZN(N289) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[3]), .ZN(n62) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[35]), .ZN(n40) );
  OAI22D1BWP30P140 U109 ( .A1(n41), .A2(n62), .B1(n46), .B2(n40), .ZN(N290) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[36]), .ZN(n42) );
  OAI22D1BWP30P140 U112 ( .A1(n47), .A2(n61), .B1(n46), .B2(n42), .ZN(N291) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[5]), .ZN(n60) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[37]), .ZN(n43) );
  OAI22D1BWP30P140 U115 ( .A1(n47), .A2(n60), .B1(n46), .B2(n43), .ZN(N292) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[6]), .ZN(n59) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[38]), .ZN(n44) );
  OAI22D1BWP30P140 U118 ( .A1(n47), .A2(n59), .B1(n46), .B2(n44), .ZN(N293) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[7]), .ZN(n58) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[39]), .ZN(n45) );
  OAI22D1BWP30P140 U121 ( .A1(n47), .A2(n58), .B1(n46), .B2(n45), .ZN(N294) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  INVD2BWP30P140 U136 ( .I(n79), .ZN(n77) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n77), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n77), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n77), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n77), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n77), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n77), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n77), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n77), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n77), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n77), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n77), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n77), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  INVD2BWP30P140 U149 ( .I(n79), .ZN(n92) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n92), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_91 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  ND2OPTIBD1BWP30P140 U3 ( .A1(n55), .A2(n54), .ZN(n56) );
  OAI22D1BWP30P140 U4 ( .A1(n18), .A2(n17), .B1(n30), .B2(n78), .ZN(N306) );
  INVD2BWP30P140 U5 ( .I(n56), .ZN(n67) );
  INVD3BWP30P140 U6 ( .I(n67), .ZN(n91) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  OAI22D1BWP30P140 U8 ( .A1(n32), .A2(n19), .B1(n30), .B2(n72), .ZN(N307) );
  OAI22D1BWP30P140 U9 ( .A1(n32), .A2(n20), .B1(n30), .B2(n71), .ZN(N308) );
  OAI22D1BWP30P140 U10 ( .A1(n32), .A2(n21), .B1(n30), .B2(n70), .ZN(N309) );
  OAI22D1BWP30P140 U11 ( .A1(n32), .A2(n22), .B1(n30), .B2(n69), .ZN(N310) );
  OAI22D1BWP30P140 U12 ( .A1(n32), .A2(n23), .B1(n30), .B2(n68), .ZN(N311) );
  OAI22D1BWP30P140 U13 ( .A1(n32), .A2(n24), .B1(n30), .B2(n73), .ZN(N312) );
  OAI22D1BWP30P140 U14 ( .A1(n32), .A2(n25), .B1(n30), .B2(n74), .ZN(N313) );
  OAI22D1BWP30P140 U15 ( .A1(n32), .A2(n26), .B1(n30), .B2(n75), .ZN(N314) );
  OAI22D1BWP30P140 U16 ( .A1(n32), .A2(n27), .B1(n30), .B2(n76), .ZN(N315) );
  OAI22D1BWP30P140 U17 ( .A1(n32), .A2(n28), .B1(n30), .B2(n77), .ZN(N316) );
  OAI22D1BWP30P140 U18 ( .A1(n32), .A2(n29), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U19 ( .A1(n32), .A2(n31), .B1(n30), .B2(n92), .ZN(N318) );
  ND2D1BWP30P140 U20 ( .A1(n1), .A2(i_en), .ZN(n51) );
  INVD1BWP30P140 U21 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U22 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U23 ( .A1(n18), .A2(n6), .B1(n40), .B2(n66), .ZN(N295) );
  OAI22D1BWP30P140 U24 ( .A1(n18), .A2(n7), .B1(n40), .B2(n65), .ZN(N296) );
  OAI22D1BWP30P140 U25 ( .A1(n18), .A2(n8), .B1(n40), .B2(n88), .ZN(N297) );
  OAI22D1BWP30P140 U26 ( .A1(n18), .A2(n9), .B1(n40), .B2(n86), .ZN(N298) );
  OAI22D1BWP30P140 U27 ( .A1(n18), .A2(n10), .B1(n40), .B2(n85), .ZN(N299) );
  OAI22D1BWP30P140 U28 ( .A1(n18), .A2(n11), .B1(n40), .B2(n84), .ZN(N300) );
  OAI22D1BWP30P140 U29 ( .A1(n18), .A2(n12), .B1(n40), .B2(n83), .ZN(N301) );
  OAI22D1BWP30P140 U30 ( .A1(n18), .A2(n13), .B1(n40), .B2(n82), .ZN(N302) );
  OAI22D1BWP30P140 U31 ( .A1(n18), .A2(n14), .B1(n40), .B2(n81), .ZN(N303) );
  OAI22D1BWP30P140 U32 ( .A1(n18), .A2(n15), .B1(n40), .B2(n80), .ZN(N304) );
  OAI22D1BWP30P140 U33 ( .A1(n18), .A2(n16), .B1(n40), .B2(n79), .ZN(N305) );
  INVD1BWP30P140 U34 ( .I(rst), .ZN(n1) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD2BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[40]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n40) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[41]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[9]), .ZN(n65) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[42]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[43]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[11]), .ZN(n86) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n85) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[13]), .ZN(n84) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[14]), .ZN(n83) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[15]), .ZN(n82) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[16]), .ZN(n81) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[17]), .ZN(n80) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[18]), .ZN(n79) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD2BWP30P140 U71 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[20]), .ZN(n72) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[21]), .ZN(n71) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[22]), .ZN(n70) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[23]), .ZN(n69) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[24]), .ZN(n68) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[25]), .ZN(n73) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[26]), .ZN(n74) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[27]), .ZN(n75) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[28]), .ZN(n76) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[29]), .ZN(n77) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U96 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U97 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD2BWP30P140 U99 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U101 ( .A1(n40), .A2(n57), .B1(n45), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[6]), .ZN(n58) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U104 ( .A1(n40), .A2(n58), .B1(n45), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[5]), .ZN(n59) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U107 ( .A1(n40), .A2(n59), .B1(n45), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U110 ( .A1(n40), .A2(n60), .B1(n45), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U113 ( .A1(n46), .A2(n61), .B1(n45), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U116 ( .A1(n46), .A2(n62), .B1(n45), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[1]), .ZN(n63) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U119 ( .A1(n46), .A2(n63), .B1(n45), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U122 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U123 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U124 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U125 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U126 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MUX2NUD1BWP30P140 U127 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n91), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n91), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n91), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n91), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n91), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n91), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n91), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  INVD2BWP30P140 U136 ( .I(n67), .ZN(n87) );
  MOAI22D1BWP30P140 U137 ( .A1(n65), .A2(n87), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U138 ( .A1(n66), .A2(n87), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n87), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n87), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n87), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n87), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n87), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n87), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n87), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n85), .A2(n87), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n86), .A2(n87), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n87), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_92 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  OAI22D1BWP30P140 U3 ( .A1(n27), .A2(n26), .B1(n31), .B2(n83), .ZN(N306) );
  INVD1BWP30P140 U4 ( .I(n57), .ZN(n75) );
  ND2D1BWP30P140 U5 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U6 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U7 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U8 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U9 ( .A1(n27), .A2(n7), .B1(n41), .B2(n93), .ZN(N295) );
  OAI22D1BWP30P140 U10 ( .A1(n27), .A2(n16), .B1(n41), .B2(n88), .ZN(N296) );
  OAI22D1BWP30P140 U11 ( .A1(n27), .A2(n17), .B1(n41), .B2(n87), .ZN(N297) );
  OAI22D1BWP30P140 U12 ( .A1(n27), .A2(n10), .B1(n41), .B2(n86), .ZN(N298) );
  OAI22D1BWP30P140 U13 ( .A1(n27), .A2(n8), .B1(n41), .B2(n76), .ZN(N299) );
  OAI22D1BWP30P140 U14 ( .A1(n27), .A2(n11), .B1(n41), .B2(n77), .ZN(N300) );
  OAI22D1BWP30P140 U15 ( .A1(n27), .A2(n9), .B1(n41), .B2(n78), .ZN(N301) );
  OAI22D1BWP30P140 U16 ( .A1(n27), .A2(n12), .B1(n41), .B2(n79), .ZN(N302) );
  OAI22D1BWP30P140 U17 ( .A1(n27), .A2(n13), .B1(n41), .B2(n80), .ZN(N303) );
  OAI22D1BWP30P140 U18 ( .A1(n27), .A2(n14), .B1(n41), .B2(n81), .ZN(N304) );
  OAI22D1BWP30P140 U19 ( .A1(n27), .A2(n15), .B1(n41), .B2(n82), .ZN(N305) );
  OAI22D1BWP30P140 U20 ( .A1(n33), .A2(n18), .B1(n31), .B2(n84), .ZN(N307) );
  OAI22D1BWP30P140 U21 ( .A1(n33), .A2(n19), .B1(n31), .B2(n85), .ZN(N308) );
  OAI22D1BWP30P140 U22 ( .A1(n33), .A2(n20), .B1(n31), .B2(n90), .ZN(N309) );
  OAI22D1BWP30P140 U23 ( .A1(n33), .A2(n21), .B1(n31), .B2(n74), .ZN(N310) );
  OAI22D1BWP30P140 U24 ( .A1(n33), .A2(n22), .B1(n31), .B2(n73), .ZN(N311) );
  OAI22D1BWP30P140 U25 ( .A1(n33), .A2(n23), .B1(n31), .B2(n72), .ZN(N312) );
  OAI22D1BWP30P140 U26 ( .A1(n33), .A2(n24), .B1(n31), .B2(n71), .ZN(N313) );
  OAI22D1BWP30P140 U27 ( .A1(n33), .A2(n30), .B1(n31), .B2(n70), .ZN(N314) );
  OAI22D1BWP30P140 U28 ( .A1(n33), .A2(n25), .B1(n31), .B2(n69), .ZN(N315) );
  OAI22D1BWP30P140 U29 ( .A1(n33), .A2(n32), .B1(n31), .B2(n68), .ZN(N316) );
  OAI22D1BWP30P140 U30 ( .A1(n33), .A2(n29), .B1(n31), .B2(n67), .ZN(N317) );
  OAI22D1BWP30P140 U31 ( .A1(n33), .A2(n28), .B1(n31), .B2(n66), .ZN(N318) );
  CKND2D2BWP30P140 U32 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U34 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U35 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U36 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U37 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U38 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U39 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U40 ( .I(n36), .ZN(n27) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[40]), .ZN(n7) );
  INR2D1BWP30P140 U42 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U43 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U44 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U45 ( .I(n34), .ZN(n41) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[8]), .ZN(n93) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[44]), .ZN(n8) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[12]), .ZN(n76) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[46]), .ZN(n9) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[14]), .ZN(n78) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[43]), .ZN(n10) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[11]), .ZN(n86) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[13]), .ZN(n77) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[47]), .ZN(n12) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[15]), .ZN(n79) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[48]), .ZN(n13) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[16]), .ZN(n80) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[49]), .ZN(n14) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[17]), .ZN(n81) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[50]), .ZN(n15) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[18]), .ZN(n82) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[41]), .ZN(n16) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[9]), .ZN(n88) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[42]), .ZN(n17) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[10]), .ZN(n87) );
  INVD2BWP30P140 U67 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[52]), .ZN(n18) );
  INVD2BWP30P140 U69 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[20]), .ZN(n84) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[53]), .ZN(n19) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[21]), .ZN(n85) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[54]), .ZN(n20) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[22]), .ZN(n90) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[55]), .ZN(n21) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[23]), .ZN(n74) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[56]), .ZN(n22) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[24]), .ZN(n73) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[57]), .ZN(n23) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[25]), .ZN(n72) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[58]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[26]), .ZN(n71) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[60]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[28]), .ZN(n69) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[51]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[19]), .ZN(n83) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[63]), .ZN(n28) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[31]), .ZN(n66) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[30]), .ZN(n67) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[59]), .ZN(n30) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[27]), .ZN(n70) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[61]), .ZN(n32) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[29]), .ZN(n68) );
  INVD1BWP30P140 U95 ( .I(n34), .ZN(n47) );
  OAI31D1BWP30P140 U96 ( .A1(n52), .A2(n53), .A3(n35), .B(n47), .ZN(N353) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[7]), .ZN(n58) );
  INVD2BWP30P140 U98 ( .I(n36), .ZN(n46) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[39]), .ZN(n37) );
  OAI22D1BWP30P140 U100 ( .A1(n41), .A2(n58), .B1(n46), .B2(n37), .ZN(N294) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[6]), .ZN(n59) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[38]), .ZN(n38) );
  OAI22D1BWP30P140 U103 ( .A1(n41), .A2(n59), .B1(n46), .B2(n38), .ZN(N293) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[5]), .ZN(n60) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[37]), .ZN(n39) );
  OAI22D1BWP30P140 U106 ( .A1(n41), .A2(n60), .B1(n46), .B2(n39), .ZN(N292) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[36]), .ZN(n40) );
  OAI22D1BWP30P140 U109 ( .A1(n41), .A2(n61), .B1(n46), .B2(n40), .ZN(N291) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[3]), .ZN(n62) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[35]), .ZN(n42) );
  OAI22D1BWP30P140 U112 ( .A1(n47), .A2(n62), .B1(n46), .B2(n42), .ZN(N290) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[2]), .ZN(n63) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[34]), .ZN(n43) );
  OAI22D1BWP30P140 U115 ( .A1(n47), .A2(n63), .B1(n46), .B2(n43), .ZN(N289) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[1]), .ZN(n65) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[33]), .ZN(n44) );
  OAI22D1BWP30P140 U118 ( .A1(n47), .A2(n65), .B1(n46), .B2(n44), .ZN(N288) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[32]), .ZN(n45) );
  OAI22D1BWP30P140 U121 ( .A1(n47), .A2(n64), .B1(n46), .B2(n45), .ZN(N287) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  INVD2BWP30P140 U136 ( .I(n75), .ZN(n89) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n89), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n89), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n89), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n89), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n89), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n89), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n89), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n89), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n89), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  INVD2BWP30P140 U146 ( .I(n75), .ZN(n92) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n92), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n92), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n92), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n92), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n92), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n92), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n92), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n92), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n89), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U156 ( .A1(n85), .A2(n89), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U157 ( .A1(n86), .A2(n92), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n87), .A2(n92), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n88), .A2(n92), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n89), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_93 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  ND2OPTIBD1BWP30P140 U3 ( .A1(n55), .A2(n54), .ZN(n56) );
  OAI22D1BWP30P140 U4 ( .A1(n29), .A2(n28), .B1(n30), .B2(n82), .ZN(N306) );
  INVD2BWP30P140 U5 ( .I(n56), .ZN(n69) );
  INVD3BWP30P140 U6 ( .I(n69), .ZN(n81) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  OAI22D1BWP30P140 U8 ( .A1(n32), .A2(n26), .B1(n30), .B2(n83), .ZN(N307) );
  OAI22D1BWP30P140 U9 ( .A1(n32), .A2(n25), .B1(n30), .B2(n84), .ZN(N308) );
  OAI22D1BWP30P140 U10 ( .A1(n32), .A2(n31), .B1(n30), .B2(n85), .ZN(N309) );
  OAI22D1BWP30P140 U11 ( .A1(n32), .A2(n21), .B1(n30), .B2(n86), .ZN(N310) );
  OAI22D1BWP30P140 U12 ( .A1(n32), .A2(n22), .B1(n30), .B2(n66), .ZN(N311) );
  OAI22D1BWP30P140 U13 ( .A1(n32), .A2(n20), .B1(n30), .B2(n65), .ZN(N312) );
  OAI22D1BWP30P140 U14 ( .A1(n32), .A2(n19), .B1(n30), .B2(n67), .ZN(N313) );
  OAI22D1BWP30P140 U15 ( .A1(n32), .A2(n18), .B1(n30), .B2(n68), .ZN(N314) );
  OAI22D1BWP30P140 U16 ( .A1(n32), .A2(n17), .B1(n30), .B2(n87), .ZN(N315) );
  OAI22D1BWP30P140 U17 ( .A1(n32), .A2(n24), .B1(n30), .B2(n88), .ZN(N316) );
  OAI22D1BWP30P140 U18 ( .A1(n32), .A2(n23), .B1(n30), .B2(n89), .ZN(N317) );
  OAI22D1BWP30P140 U19 ( .A1(n32), .A2(n27), .B1(n30), .B2(n92), .ZN(N318) );
  ND2D1BWP30P140 U20 ( .A1(n1), .A2(i_en), .ZN(n51) );
  INVD1BWP30P140 U21 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U22 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U23 ( .A1(n29), .A2(n16), .B1(n41), .B2(n77), .ZN(N295) );
  OAI22D1BWP30P140 U24 ( .A1(n29), .A2(n15), .B1(n41), .B2(n76), .ZN(N296) );
  OAI22D1BWP30P140 U25 ( .A1(n29), .A2(n14), .B1(n41), .B2(n70), .ZN(N297) );
  OAI22D1BWP30P140 U26 ( .A1(n29), .A2(n12), .B1(n41), .B2(n71), .ZN(N298) );
  OAI22D1BWP30P140 U27 ( .A1(n29), .A2(n10), .B1(n41), .B2(n72), .ZN(N299) );
  OAI22D1BWP30P140 U28 ( .A1(n29), .A2(n8), .B1(n41), .B2(n73), .ZN(N300) );
  OAI22D1BWP30P140 U29 ( .A1(n29), .A2(n7), .B1(n41), .B2(n74), .ZN(N301) );
  OAI22D1BWP30P140 U30 ( .A1(n29), .A2(n6), .B1(n41), .B2(n75), .ZN(N302) );
  OAI22D1BWP30P140 U31 ( .A1(n29), .A2(n9), .B1(n41), .B2(n78), .ZN(N303) );
  OAI22D1BWP30P140 U32 ( .A1(n29), .A2(n11), .B1(n41), .B2(n79), .ZN(N304) );
  OAI22D1BWP30P140 U33 ( .A1(n29), .A2(n13), .B1(n41), .B2(n80), .ZN(N305) );
  INVD1BWP30P140 U34 ( .I(rst), .ZN(n1) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD2BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n29) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[47]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n41) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[15]), .ZN(n75) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[46]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[14]), .ZN(n74) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[45]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[13]), .ZN(n73) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[48]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[16]), .ZN(n78) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[44]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[12]), .ZN(n72) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[49]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[17]), .ZN(n79) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[43]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[11]), .ZN(n71) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[50]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[18]), .ZN(n80) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[42]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[10]), .ZN(n70) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[41]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[9]), .ZN(n76) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[40]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[8]), .ZN(n77) );
  INVD2BWP30P140 U68 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[60]), .ZN(n17) );
  INVD2BWP30P140 U70 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[28]), .ZN(n87) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[59]), .ZN(n18) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[27]), .ZN(n68) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[58]), .ZN(n19) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[26]), .ZN(n67) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[57]), .ZN(n20) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[25]), .ZN(n65) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[55]), .ZN(n21) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[23]), .ZN(n86) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[56]), .ZN(n22) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[24]), .ZN(n66) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[62]), .ZN(n23) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[30]), .ZN(n89) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[61]), .ZN(n24) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[29]), .ZN(n88) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[53]), .ZN(n25) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[21]), .ZN(n84) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[52]), .ZN(n26) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[20]), .ZN(n83) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[63]), .ZN(n27) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[31]), .ZN(n92) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[51]), .ZN(n28) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[19]), .ZN(n82) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[54]), .ZN(n31) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[22]), .ZN(n85) );
  INVD1BWP30P140 U96 ( .I(n33), .ZN(n46) );
  OAI31D1BWP30P140 U97 ( .A1(n51), .A2(n52), .A3(n34), .B(n46), .ZN(N353) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD2BWP30P140 U99 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[32]), .ZN(n36) );
  OAI22D1BWP30P140 U101 ( .A1(n46), .A2(n57), .B1(n45), .B2(n36), .ZN(N287) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[39]), .ZN(n37) );
  OAI22D1BWP30P140 U104 ( .A1(n41), .A2(n64), .B1(n45), .B2(n37), .ZN(N294) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[38]), .ZN(n38) );
  OAI22D1BWP30P140 U107 ( .A1(n41), .A2(n63), .B1(n45), .B2(n38), .ZN(N293) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[37]), .ZN(n39) );
  OAI22D1BWP30P140 U110 ( .A1(n41), .A2(n62), .B1(n45), .B2(n39), .ZN(N292) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[36]), .ZN(n40) );
  OAI22D1BWP30P140 U113 ( .A1(n41), .A2(n61), .B1(n45), .B2(n40), .ZN(N291) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[35]), .ZN(n42) );
  OAI22D1BWP30P140 U116 ( .A1(n46), .A2(n60), .B1(n45), .B2(n42), .ZN(N290) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[34]), .ZN(n43) );
  OAI22D1BWP30P140 U119 ( .A1(n46), .A2(n59), .B1(n45), .B2(n43), .ZN(N289) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[33]), .ZN(n44) );
  OAI22D1BWP30P140 U122 ( .A1(n46), .A2(n58), .B1(n45), .B2(n44), .ZN(N288) );
  INVD1BWP30P140 U123 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U124 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U125 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U126 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MUX2NUD1BWP30P140 U127 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n81), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n81), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n81), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n81), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n81), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n81), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n81), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n81), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  INVD2BWP30P140 U136 ( .I(n69), .ZN(n91) );
  MOAI22D1BWP30P140 U137 ( .A1(n65), .A2(n91), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U138 ( .A1(n66), .A2(n91), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U139 ( .A1(n67), .A2(n91), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U140 ( .A1(n68), .A2(n91), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n81), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n81), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n81), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n81), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n81), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n81), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n81), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n81), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n81), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n81), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n81), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n81), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_94 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n33), .A2(n32), .B1(n31), .B2(n80), .ZN(N306) );
  INVD1BWP30P140 U4 ( .I(n57), .ZN(n79) );
  ND2D1BWP30P140 U5 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U6 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U7 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U8 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U9 ( .A1(n33), .A2(n16), .B1(n47), .B2(n93), .ZN(N295) );
  OAI22D1BWP30P140 U10 ( .A1(n33), .A2(n15), .B1(n47), .B2(n90), .ZN(N296) );
  OAI22D1BWP30P140 U11 ( .A1(n33), .A2(n14), .B1(n47), .B2(n89), .ZN(N297) );
  OAI22D1BWP30P140 U12 ( .A1(n33), .A2(n13), .B1(n47), .B2(n88), .ZN(N298) );
  OAI22D1BWP30P140 U13 ( .A1(n33), .A2(n12), .B1(n47), .B2(n87), .ZN(N299) );
  OAI22D1BWP30P140 U14 ( .A1(n33), .A2(n11), .B1(n47), .B2(n86), .ZN(N300) );
  OAI22D1BWP30P140 U15 ( .A1(n33), .A2(n10), .B1(n47), .B2(n85), .ZN(N301) );
  OAI22D1BWP30P140 U16 ( .A1(n33), .A2(n9), .B1(n47), .B2(n84), .ZN(N302) );
  OAI22D1BWP30P140 U17 ( .A1(n33), .A2(n8), .B1(n47), .B2(n83), .ZN(N303) );
  OAI22D1BWP30P140 U18 ( .A1(n33), .A2(n17), .B1(n47), .B2(n82), .ZN(N304) );
  OAI22D1BWP30P140 U19 ( .A1(n33), .A2(n7), .B1(n47), .B2(n81), .ZN(N305) );
  OAI22D1BWP30P140 U20 ( .A1(n30), .A2(n29), .B1(n31), .B2(n78), .ZN(N307) );
  OAI22D1BWP30P140 U21 ( .A1(n30), .A2(n28), .B1(n31), .B2(n76), .ZN(N308) );
  OAI22D1BWP30P140 U22 ( .A1(n30), .A2(n27), .B1(n31), .B2(n75), .ZN(N309) );
  OAI22D1BWP30P140 U23 ( .A1(n30), .A2(n26), .B1(n31), .B2(n74), .ZN(N310) );
  OAI22D1BWP30P140 U24 ( .A1(n30), .A2(n25), .B1(n31), .B2(n73), .ZN(N311) );
  OAI22D1BWP30P140 U25 ( .A1(n30), .A2(n24), .B1(n31), .B2(n72), .ZN(N312) );
  OAI22D1BWP30P140 U26 ( .A1(n30), .A2(n23), .B1(n31), .B2(n71), .ZN(N313) );
  OAI22D1BWP30P140 U27 ( .A1(n30), .A2(n22), .B1(n31), .B2(n70), .ZN(N314) );
  OAI22D1BWP30P140 U28 ( .A1(n30), .A2(n21), .B1(n31), .B2(n69), .ZN(N315) );
  OAI22D1BWP30P140 U29 ( .A1(n30), .A2(n20), .B1(n31), .B2(n68), .ZN(N316) );
  OAI22D1BWP30P140 U30 ( .A1(n30), .A2(n19), .B1(n31), .B2(n67), .ZN(N317) );
  OAI22D1BWP30P140 U31 ( .A1(n30), .A2(n18), .B1(n31), .B2(n66), .ZN(N318) );
  CKND2D2BWP30P140 U32 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U34 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U35 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U36 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U37 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U38 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U39 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U40 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[50]), .ZN(n7) );
  INR2D1BWP30P140 U42 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U43 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U44 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U45 ( .I(n34), .ZN(n47) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[18]), .ZN(n81) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[48]), .ZN(n8) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[16]), .ZN(n83) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[47]), .ZN(n9) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[15]), .ZN(n84) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[46]), .ZN(n10) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[14]), .ZN(n85) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[45]), .ZN(n11) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[13]), .ZN(n86) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n12) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n87) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[43]), .ZN(n13) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[11]), .ZN(n88) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[42]), .ZN(n14) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[10]), .ZN(n89) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[41]), .ZN(n15) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[9]), .ZN(n90) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[40]), .ZN(n16) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[8]), .ZN(n93) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n17) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n82) );
  INVD2BWP30P140 U67 ( .I(n36), .ZN(n30) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[63]), .ZN(n18) );
  INVD2BWP30P140 U69 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[31]), .ZN(n66) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[62]), .ZN(n19) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[30]), .ZN(n67) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[61]), .ZN(n20) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[29]), .ZN(n68) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[60]), .ZN(n21) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[28]), .ZN(n69) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[59]), .ZN(n22) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[27]), .ZN(n70) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[58]), .ZN(n23) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[26]), .ZN(n71) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[25]), .ZN(n72) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[56]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[24]), .ZN(n73) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[55]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[23]), .ZN(n74) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[54]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[22]), .ZN(n75) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[53]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[21]), .ZN(n76) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[52]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[20]), .ZN(n78) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[51]), .ZN(n32) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[19]), .ZN(n80) );
  INVD1BWP30P140 U95 ( .I(n34), .ZN(n41) );
  OAI31D1BWP30P140 U96 ( .A1(n52), .A2(n53), .A3(n35), .B(n41), .ZN(N353) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[0]), .ZN(n63) );
  INVD2BWP30P140 U98 ( .I(n36), .ZN(n46) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[32]), .ZN(n37) );
  OAI22D1BWP30P140 U100 ( .A1(n41), .A2(n63), .B1(n46), .B2(n37), .ZN(N287) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[1]), .ZN(n64) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[33]), .ZN(n38) );
  OAI22D1BWP30P140 U103 ( .A1(n41), .A2(n64), .B1(n46), .B2(n38), .ZN(N288) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[2]), .ZN(n65) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[34]), .ZN(n39) );
  OAI22D1BWP30P140 U106 ( .A1(n41), .A2(n65), .B1(n46), .B2(n39), .ZN(N289) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[3]), .ZN(n58) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[35]), .ZN(n40) );
  OAI22D1BWP30P140 U109 ( .A1(n41), .A2(n58), .B1(n46), .B2(n40), .ZN(N290) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[4]), .ZN(n59) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[36]), .ZN(n42) );
  OAI22D1BWP30P140 U112 ( .A1(n47), .A2(n59), .B1(n46), .B2(n42), .ZN(N291) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[5]), .ZN(n60) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[37]), .ZN(n43) );
  OAI22D1BWP30P140 U115 ( .A1(n47), .A2(n60), .B1(n46), .B2(n43), .ZN(N292) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[6]), .ZN(n61) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[38]), .ZN(n44) );
  OAI22D1BWP30P140 U118 ( .A1(n47), .A2(n61), .B1(n46), .B2(n44), .ZN(N293) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[7]), .ZN(n62) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[39]), .ZN(n45) );
  OAI22D1BWP30P140 U121 ( .A1(n47), .A2(n62), .B1(n46), .B2(n45), .ZN(N294) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  INVD2BWP30P140 U136 ( .I(n79), .ZN(n77) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n77), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n77), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n77), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n77), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n77), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n77), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n77), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n77), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n77), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n77), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n77), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n77), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  INVD2BWP30P140 U149 ( .I(n79), .ZN(n92) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n92), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_95 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  ND2OPTIBD1BWP30P140 U3 ( .A1(n55), .A2(n54), .ZN(n56) );
  OAI22D1BWP30P140 U4 ( .A1(n18), .A2(n17), .B1(n30), .B2(n79), .ZN(N306) );
  INVD2BWP30P140 U5 ( .I(n56), .ZN(n78) );
  INVD3BWP30P140 U6 ( .I(n78), .ZN(n91) );
  NR2D1BWP30P140 U7 ( .A1(n51), .A2(i_cmd[1]), .ZN(n55) );
  OAI22D1BWP30P140 U8 ( .A1(n32), .A2(n19), .B1(n30), .B2(n77), .ZN(N307) );
  OAI22D1BWP30P140 U9 ( .A1(n32), .A2(n20), .B1(n30), .B2(n75), .ZN(N308) );
  OAI22D1BWP30P140 U10 ( .A1(n32), .A2(n21), .B1(n30), .B2(n74), .ZN(N309) );
  OAI22D1BWP30P140 U11 ( .A1(n32), .A2(n22), .B1(n30), .B2(n73), .ZN(N310) );
  OAI22D1BWP30P140 U12 ( .A1(n32), .A2(n23), .B1(n30), .B2(n72), .ZN(N311) );
  OAI22D1BWP30P140 U13 ( .A1(n32), .A2(n24), .B1(n30), .B2(n71), .ZN(N312) );
  OAI22D1BWP30P140 U14 ( .A1(n32), .A2(n25), .B1(n30), .B2(n70), .ZN(N313) );
  OAI22D1BWP30P140 U15 ( .A1(n32), .A2(n26), .B1(n30), .B2(n69), .ZN(N314) );
  OAI22D1BWP30P140 U16 ( .A1(n32), .A2(n27), .B1(n30), .B2(n68), .ZN(N315) );
  OAI22D1BWP30P140 U17 ( .A1(n32), .A2(n28), .B1(n30), .B2(n67), .ZN(N316) );
  OAI22D1BWP30P140 U18 ( .A1(n32), .A2(n29), .B1(n30), .B2(n66), .ZN(N317) );
  OAI22D1BWP30P140 U19 ( .A1(n32), .A2(n31), .B1(n30), .B2(n65), .ZN(N318) );
  ND2D1BWP30P140 U20 ( .A1(n1), .A2(i_en), .ZN(n51) );
  INVD1BWP30P140 U21 ( .I(i_cmd[0]), .ZN(n34) );
  INVD1BWP30P140 U22 ( .I(n90), .ZN(n49) );
  OAI22D1BWP30P140 U23 ( .A1(n18), .A2(n16), .B1(n46), .B2(n92), .ZN(N295) );
  OAI22D1BWP30P140 U24 ( .A1(n18), .A2(n15), .B1(n46), .B2(n89), .ZN(N296) );
  OAI22D1BWP30P140 U25 ( .A1(n18), .A2(n14), .B1(n46), .B2(n88), .ZN(N297) );
  OAI22D1BWP30P140 U26 ( .A1(n18), .A2(n13), .B1(n46), .B2(n87), .ZN(N298) );
  OAI22D1BWP30P140 U27 ( .A1(n18), .A2(n6), .B1(n46), .B2(n86), .ZN(N299) );
  OAI22D1BWP30P140 U28 ( .A1(n18), .A2(n7), .B1(n46), .B2(n85), .ZN(N300) );
  OAI22D1BWP30P140 U29 ( .A1(n18), .A2(n8), .B1(n46), .B2(n84), .ZN(N301) );
  OAI22D1BWP30P140 U30 ( .A1(n18), .A2(n9), .B1(n46), .B2(n83), .ZN(N302) );
  OAI22D1BWP30P140 U31 ( .A1(n18), .A2(n10), .B1(n46), .B2(n82), .ZN(N303) );
  OAI22D1BWP30P140 U32 ( .A1(n18), .A2(n11), .B1(n46), .B2(n81), .ZN(N304) );
  OAI22D1BWP30P140 U33 ( .A1(n18), .A2(n12), .B1(n46), .B2(n80), .ZN(N305) );
  INVD1BWP30P140 U34 ( .I(rst), .ZN(n1) );
  NR2D1BWP30P140 U35 ( .A1(n51), .A2(n34), .ZN(n3) );
  INVD1BWP30P140 U36 ( .I(i_valid[0]), .ZN(n53) );
  INVD2BWP30P140 U37 ( .I(i_valid[1]), .ZN(n52) );
  MUX2NUD1BWP30P140 U38 ( .I0(n53), .I1(n52), .S(i_cmd[1]), .ZN(n2) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n3), .A2(n2), .ZN(n4) );
  INVD2BWP30P140 U40 ( .I(n4), .ZN(n35) );
  INVD2BWP30P140 U41 ( .I(n35), .ZN(n18) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[44]), .ZN(n6) );
  INR2D1BWP30P140 U43 ( .A1(i_valid[0]), .B1(n51), .ZN(n47) );
  CKND2D2BWP30P140 U44 ( .A1(n47), .A2(n34), .ZN(n5) );
  INVD2BWP30P140 U45 ( .I(n5), .ZN(n33) );
  INVD2BWP30P140 U46 ( .I(n33), .ZN(n46) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[12]), .ZN(n86) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[45]), .ZN(n7) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[13]), .ZN(n85) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[46]), .ZN(n8) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[14]), .ZN(n84) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[47]), .ZN(n9) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[15]), .ZN(n83) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[48]), .ZN(n10) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[16]), .ZN(n82) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[49]), .ZN(n11) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[17]), .ZN(n81) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[50]), .ZN(n12) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[18]), .ZN(n80) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[43]), .ZN(n13) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[11]), .ZN(n87) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[42]), .ZN(n14) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[10]), .ZN(n88) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[41]), .ZN(n15) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[9]), .ZN(n89) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[40]), .ZN(n16) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[8]), .ZN(n92) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[51]), .ZN(n17) );
  INVD2BWP30P140 U69 ( .I(n33), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[19]), .ZN(n79) );
  INVD2BWP30P140 U71 ( .I(n35), .ZN(n32) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[52]), .ZN(n19) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[21]), .ZN(n75) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[54]), .ZN(n21) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[23]), .ZN(n73) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[24]), .ZN(n72) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[25]), .ZN(n71) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[26]), .ZN(n70) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[27]), .ZN(n69) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[28]), .ZN(n68) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[29]), .ZN(n67) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[30]), .ZN(n66) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[31]), .ZN(n65) );
  INVD1BWP30P140 U96 ( .I(n33), .ZN(n41) );
  OAI31D1BWP30P140 U97 ( .A1(n51), .A2(n52), .A3(n34), .B(n41), .ZN(N353) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD2BWP30P140 U99 ( .I(n35), .ZN(n45) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[36]), .ZN(n36) );
  OAI22D1BWP30P140 U101 ( .A1(n46), .A2(n61), .B1(n45), .B2(n36), .ZN(N291) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[35]), .ZN(n37) );
  OAI22D1BWP30P140 U104 ( .A1(n41), .A2(n60), .B1(n45), .B2(n37), .ZN(N290) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[34]), .ZN(n38) );
  OAI22D1BWP30P140 U107 ( .A1(n41), .A2(n59), .B1(n45), .B2(n38), .ZN(N289) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[33]), .ZN(n39) );
  OAI22D1BWP30P140 U110 ( .A1(n41), .A2(n58), .B1(n45), .B2(n39), .ZN(N288) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[0]), .ZN(n57) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[32]), .ZN(n40) );
  OAI22D1BWP30P140 U113 ( .A1(n41), .A2(n57), .B1(n45), .B2(n40), .ZN(N287) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[37]), .ZN(n42) );
  OAI22D1BWP30P140 U116 ( .A1(n46), .A2(n62), .B1(n45), .B2(n42), .ZN(N292) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[38]), .ZN(n43) );
  OAI22D1BWP30P140 U119 ( .A1(n46), .A2(n63), .B1(n45), .B2(n43), .ZN(N293) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[39]), .ZN(n44) );
  OAI22D1BWP30P140 U122 ( .A1(n46), .A2(n64), .B1(n45), .B2(n44), .ZN(N294) );
  INVD1BWP30P140 U123 ( .I(n47), .ZN(n50) );
  INVD1BWP30P140 U124 ( .I(n51), .ZN(n48) );
  AN3D4BWP30P140 U125 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n48), .Z(n90) );
  OAI21D1BWP30P140 U126 ( .A1(n50), .A2(i_cmd[1]), .B(n49), .ZN(N354) );
  MUX2NUD1BWP30P140 U127 ( .I0(n53), .I1(n52), .S(i_cmd[0]), .ZN(n54) );
  MOAI22D1BWP30P140 U128 ( .A1(n57), .A2(n91), .B1(i_data_bus[32]), .B2(n90), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n91), .B1(i_data_bus[33]), .B2(n90), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n91), .B1(i_data_bus[34]), .B2(n90), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n91), .B1(i_data_bus[35]), .B2(n90), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n91), .B1(i_data_bus[36]), .B2(n90), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n91), .B1(i_data_bus[37]), .B2(n90), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n91), .B1(i_data_bus[38]), .B2(n90), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n91), .B1(i_data_bus[39]), .B2(n90), 
        .ZN(N326) );
  INVD2BWP30P140 U136 ( .I(n78), .ZN(n76) );
  MOAI22D1BWP30P140 U137 ( .A1(n65), .A2(n76), .B1(i_data_bus[63]), .B2(n90), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U138 ( .A1(n66), .A2(n76), .B1(i_data_bus[62]), .B2(n90), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U139 ( .A1(n67), .A2(n76), .B1(i_data_bus[61]), .B2(n90), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U140 ( .A1(n68), .A2(n76), .B1(i_data_bus[60]), .B2(n90), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U141 ( .A1(n69), .A2(n76), .B1(i_data_bus[59]), .B2(n90), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U142 ( .A1(n70), .A2(n76), .B1(i_data_bus[58]), .B2(n90), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U143 ( .A1(n71), .A2(n76), .B1(i_data_bus[57]), .B2(n90), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U144 ( .A1(n72), .A2(n76), .B1(i_data_bus[56]), .B2(n90), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U145 ( .A1(n73), .A2(n76), .B1(i_data_bus[55]), .B2(n90), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U146 ( .A1(n74), .A2(n76), .B1(i_data_bus[54]), .B2(n90), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U147 ( .A1(n75), .A2(n76), .B1(i_data_bus[53]), .B2(n90), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n76), .B1(i_data_bus[52]), .B2(n90), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U149 ( .A1(n79), .A2(n91), .B1(i_data_bus[51]), .B2(n90), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n91), .B1(i_data_bus[50]), .B2(n90), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n91), .B1(i_data_bus[49]), .B2(n90), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n91), .B1(i_data_bus[48]), .B2(n90), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n91), .B1(i_data_bus[47]), .B2(n90), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n91), .B1(i_data_bus[46]), .B2(n90), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n91), .B1(i_data_bus[45]), .B2(n90), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n91), .B1(i_data_bus[44]), .B2(n90), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n91), .B1(i_data_bus[43]), .B2(n90), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n91), .B1(i_data_bus[42]), .B2(n90), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n91), .B1(i_data_bus[41]), .B2(n90), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U160 ( .A1(n92), .A2(n91), .B1(i_data_bus[40]), .B2(n90), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_96 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  OAI22D1BWP30P140 U3 ( .A1(n33), .A2(n32), .B1(n31), .B2(n80), .ZN(N306) );
  INVD1BWP30P140 U4 ( .I(n57), .ZN(n79) );
  ND2D1BWP30P140 U5 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U6 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U7 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U8 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U9 ( .A1(n33), .A2(n17), .B1(n47), .B2(n93), .ZN(N295) );
  OAI22D1BWP30P140 U10 ( .A1(n33), .A2(n16), .B1(n47), .B2(n90), .ZN(N296) );
  OAI22D1BWP30P140 U11 ( .A1(n33), .A2(n15), .B1(n47), .B2(n89), .ZN(N297) );
  OAI22D1BWP30P140 U12 ( .A1(n33), .A2(n14), .B1(n47), .B2(n88), .ZN(N298) );
  OAI22D1BWP30P140 U13 ( .A1(n33), .A2(n13), .B1(n47), .B2(n87), .ZN(N299) );
  OAI22D1BWP30P140 U14 ( .A1(n33), .A2(n12), .B1(n47), .B2(n86), .ZN(N300) );
  OAI22D1BWP30P140 U15 ( .A1(n33), .A2(n11), .B1(n47), .B2(n85), .ZN(N301) );
  OAI22D1BWP30P140 U16 ( .A1(n33), .A2(n10), .B1(n47), .B2(n84), .ZN(N302) );
  OAI22D1BWP30P140 U17 ( .A1(n33), .A2(n9), .B1(n47), .B2(n83), .ZN(N303) );
  OAI22D1BWP30P140 U18 ( .A1(n33), .A2(n8), .B1(n47), .B2(n82), .ZN(N304) );
  OAI22D1BWP30P140 U19 ( .A1(n33), .A2(n7), .B1(n47), .B2(n81), .ZN(N305) );
  OAI22D1BWP30P140 U20 ( .A1(n30), .A2(n29), .B1(n31), .B2(n78), .ZN(N307) );
  OAI22D1BWP30P140 U21 ( .A1(n30), .A2(n28), .B1(n31), .B2(n76), .ZN(N308) );
  OAI22D1BWP30P140 U22 ( .A1(n30), .A2(n27), .B1(n31), .B2(n75), .ZN(N309) );
  OAI22D1BWP30P140 U23 ( .A1(n30), .A2(n26), .B1(n31), .B2(n74), .ZN(N310) );
  OAI22D1BWP30P140 U24 ( .A1(n30), .A2(n25), .B1(n31), .B2(n73), .ZN(N311) );
  OAI22D1BWP30P140 U25 ( .A1(n30), .A2(n24), .B1(n31), .B2(n72), .ZN(N312) );
  OAI22D1BWP30P140 U26 ( .A1(n30), .A2(n23), .B1(n31), .B2(n71), .ZN(N313) );
  OAI22D1BWP30P140 U27 ( .A1(n30), .A2(n22), .B1(n31), .B2(n70), .ZN(N314) );
  OAI22D1BWP30P140 U28 ( .A1(n30), .A2(n21), .B1(n31), .B2(n69), .ZN(N315) );
  OAI22D1BWP30P140 U29 ( .A1(n30), .A2(n20), .B1(n31), .B2(n68), .ZN(N316) );
  OAI22D1BWP30P140 U30 ( .A1(n30), .A2(n19), .B1(n31), .B2(n67), .ZN(N317) );
  OAI22D1BWP30P140 U31 ( .A1(n30), .A2(n18), .B1(n31), .B2(n66), .ZN(N318) );
  CKND2D2BWP30P140 U32 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U34 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U35 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U36 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U37 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U38 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U39 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U40 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[50]), .ZN(n7) );
  INR2D1BWP30P140 U42 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U43 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U44 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U45 ( .I(n34), .ZN(n47) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[18]), .ZN(n81) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[49]), .ZN(n8) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[17]), .ZN(n82) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[48]), .ZN(n9) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[16]), .ZN(n83) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[47]), .ZN(n10) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[15]), .ZN(n84) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[46]), .ZN(n11) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[14]), .ZN(n85) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[13]), .ZN(n86) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[44]), .ZN(n13) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[12]), .ZN(n87) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[43]), .ZN(n14) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[11]), .ZN(n88) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[42]), .ZN(n15) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[10]), .ZN(n89) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[41]), .ZN(n16) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[9]), .ZN(n90) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[40]), .ZN(n17) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[8]), .ZN(n93) );
  INVD2BWP30P140 U67 ( .I(n36), .ZN(n30) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[63]), .ZN(n18) );
  INVD2BWP30P140 U69 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[31]), .ZN(n66) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[62]), .ZN(n19) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[30]), .ZN(n67) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[61]), .ZN(n20) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[29]), .ZN(n68) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[60]), .ZN(n21) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[28]), .ZN(n69) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[59]), .ZN(n22) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[27]), .ZN(n70) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[58]), .ZN(n23) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[26]), .ZN(n71) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[25]), .ZN(n72) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[56]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[24]), .ZN(n73) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[55]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[23]), .ZN(n74) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[54]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[22]), .ZN(n75) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[53]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[21]), .ZN(n76) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[52]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[20]), .ZN(n78) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[51]), .ZN(n32) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[19]), .ZN(n80) );
  INVD1BWP30P140 U95 ( .I(n34), .ZN(n41) );
  OAI31D1BWP30P140 U96 ( .A1(n52), .A2(n53), .A3(n35), .B(n41), .ZN(N353) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[0]), .ZN(n61) );
  INVD2BWP30P140 U98 ( .I(n36), .ZN(n46) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[32]), .ZN(n37) );
  OAI22D1BWP30P140 U100 ( .A1(n41), .A2(n61), .B1(n46), .B2(n37), .ZN(N287) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[1]), .ZN(n62) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[33]), .ZN(n38) );
  OAI22D1BWP30P140 U103 ( .A1(n41), .A2(n62), .B1(n46), .B2(n38), .ZN(N288) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[2]), .ZN(n63) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[34]), .ZN(n39) );
  OAI22D1BWP30P140 U106 ( .A1(n41), .A2(n63), .B1(n46), .B2(n39), .ZN(N289) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[3]), .ZN(n64) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[35]), .ZN(n40) );
  OAI22D1BWP30P140 U109 ( .A1(n41), .A2(n64), .B1(n46), .B2(n40), .ZN(N290) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[4]), .ZN(n58) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[36]), .ZN(n42) );
  OAI22D1BWP30P140 U112 ( .A1(n47), .A2(n58), .B1(n46), .B2(n42), .ZN(N291) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[5]), .ZN(n60) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[37]), .ZN(n43) );
  OAI22D1BWP30P140 U115 ( .A1(n47), .A2(n60), .B1(n46), .B2(n43), .ZN(N292) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[7]), .ZN(n65) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[39]), .ZN(n44) );
  OAI22D1BWP30P140 U118 ( .A1(n47), .A2(n65), .B1(n46), .B2(n44), .ZN(N294) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[6]), .ZN(n59) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[38]), .ZN(n45) );
  OAI22D1BWP30P140 U121 ( .A1(n47), .A2(n59), .B1(n46), .B2(n45), .ZN(N293) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  INVD2BWP30P140 U136 ( .I(n79), .ZN(n77) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n77), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n77), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n77), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n77), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n77), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n77), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n77), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n77), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n77), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n77), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n77), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n77), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  INVD2BWP30P140 U149 ( .I(n79), .ZN(n92) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n92), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_97 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD2BWP30P140 U3 ( .I(n36), .ZN(n46) );
  OAI22D1BWP30P140 U4 ( .A1(n47), .A2(n60), .B1(n46), .B2(n45), .ZN(N287) );
  OAI22D1BWP30P140 U5 ( .A1(n23), .A2(n22), .B1(n31), .B2(n69), .ZN(N306) );
  INVD1BWP30P140 U6 ( .I(n57), .ZN(n71) );
  ND2D1BWP30P140 U7 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U9 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U10 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U11 ( .A1(n23), .A2(n17), .B1(n41), .B2(n76), .ZN(N295) );
  OAI22D1BWP30P140 U12 ( .A1(n23), .A2(n16), .B1(n41), .B2(n75), .ZN(N296) );
  OAI22D1BWP30P140 U13 ( .A1(n23), .A2(n15), .B1(n41), .B2(n74), .ZN(N297) );
  OAI22D1BWP30P140 U14 ( .A1(n23), .A2(n14), .B1(n41), .B2(n70), .ZN(N298) );
  OAI22D1BWP30P140 U15 ( .A1(n23), .A2(n13), .B1(n41), .B2(n67), .ZN(N299) );
  OAI22D1BWP30P140 U16 ( .A1(n23), .A2(n12), .B1(n41), .B2(n82), .ZN(N300) );
  OAI22D1BWP30P140 U17 ( .A1(n23), .A2(n11), .B1(n41), .B2(n80), .ZN(N301) );
  OAI22D1BWP30P140 U18 ( .A1(n23), .A2(n10), .B1(n41), .B2(n78), .ZN(N302) );
  OAI22D1BWP30P140 U19 ( .A1(n23), .A2(n9), .B1(n41), .B2(n79), .ZN(N303) );
  OAI22D1BWP30P140 U20 ( .A1(n23), .A2(n8), .B1(n41), .B2(n66), .ZN(N304) );
  OAI22D1BWP30P140 U21 ( .A1(n23), .A2(n7), .B1(n41), .B2(n68), .ZN(N305) );
  OAI22D1BWP30P140 U22 ( .A1(n33), .A2(n21), .B1(n31), .B2(n77), .ZN(N307) );
  OAI22D1BWP30P140 U23 ( .A1(n33), .A2(n20), .B1(n31), .B2(n72), .ZN(N308) );
  OAI22D1BWP30P140 U24 ( .A1(n33), .A2(n19), .B1(n31), .B2(n73), .ZN(N309) );
  OAI22D1BWP30P140 U25 ( .A1(n33), .A2(n18), .B1(n31), .B2(n83), .ZN(N310) );
  OAI22D1BWP30P140 U26 ( .A1(n33), .A2(n24), .B1(n31), .B2(n84), .ZN(N311) );
  OAI22D1BWP30P140 U27 ( .A1(n33), .A2(n25), .B1(n31), .B2(n93), .ZN(N312) );
  OAI22D1BWP30P140 U28 ( .A1(n33), .A2(n32), .B1(n31), .B2(n90), .ZN(N313) );
  OAI22D1BWP30P140 U29 ( .A1(n33), .A2(n27), .B1(n31), .B2(n89), .ZN(N314) );
  OAI22D1BWP30P140 U30 ( .A1(n33), .A2(n29), .B1(n31), .B2(n88), .ZN(N315) );
  OAI22D1BWP30P140 U31 ( .A1(n33), .A2(n30), .B1(n31), .B2(n87), .ZN(N316) );
  OAI22D1BWP30P140 U32 ( .A1(n33), .A2(n26), .B1(n31), .B2(n86), .ZN(N317) );
  OAI22D1BWP30P140 U33 ( .A1(n33), .A2(n28), .B1(n31), .B2(n85), .ZN(N318) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n23) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[50]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n41) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[18]), .ZN(n68) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[49]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[17]), .ZN(n66) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[48]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[16]), .ZN(n79) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[47]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[15]), .ZN(n78) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[46]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[14]), .ZN(n80) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n82) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[44]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[12]), .ZN(n67) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[43]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[11]), .ZN(n70) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[42]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[10]), .ZN(n74) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[41]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[9]), .ZN(n75) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[40]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[8]), .ZN(n76) );
  INVD2BWP30P140 U69 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[55]), .ZN(n18) );
  INVD2BWP30P140 U71 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[23]), .ZN(n83) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[54]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[22]), .ZN(n73) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n72) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[52]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[20]), .ZN(n77) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[51]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[19]), .ZN(n69) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n84) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n93) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[62]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[30]), .ZN(n86) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n89) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[63]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[31]), .ZN(n85) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[60]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[28]), .ZN(n88) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[61]), .ZN(n30) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[29]), .ZN(n87) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[58]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[26]), .ZN(n90) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n47) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n47), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n58) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[39]), .ZN(n37) );
  OAI22D1BWP30P140 U101 ( .A1(n41), .A2(n58), .B1(n46), .B2(n37), .ZN(N294) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[6]), .ZN(n59) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[38]), .ZN(n38) );
  OAI22D1BWP30P140 U104 ( .A1(n41), .A2(n59), .B1(n46), .B2(n38), .ZN(N293) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[5]), .ZN(n65) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[37]), .ZN(n39) );
  OAI22D1BWP30P140 U107 ( .A1(n41), .A2(n65), .B1(n46), .B2(n39), .ZN(N292) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[4]), .ZN(n64) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[36]), .ZN(n40) );
  OAI22D1BWP30P140 U110 ( .A1(n41), .A2(n64), .B1(n46), .B2(n40), .ZN(N291) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[3]), .ZN(n63) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[35]), .ZN(n42) );
  OAI22D1BWP30P140 U113 ( .A1(n47), .A2(n63), .B1(n46), .B2(n42), .ZN(N290) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[2]), .ZN(n62) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[34]), .ZN(n43) );
  OAI22D1BWP30P140 U116 ( .A1(n47), .A2(n62), .B1(n46), .B2(n43), .ZN(N289) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[1]), .ZN(n61) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[33]), .ZN(n44) );
  OAI22D1BWP30P140 U119 ( .A1(n47), .A2(n61), .B1(n46), .B2(n44), .ZN(N288) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[0]), .ZN(n60) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[32]), .ZN(n45) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  INVD2BWP30P140 U136 ( .I(n71), .ZN(n81) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n81), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n81), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n81), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n81), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n81), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  INVD2BWP30P140 U142 ( .I(n71), .ZN(n92) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n92), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n92), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n81), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n81), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n81), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n92), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n81), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n81), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n81), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n81), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_98 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD4BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n33), .A2(n32), .B1(n31), .B2(n80), .ZN(N306) );
  INVD1BWP30P140 U4 ( .I(n57), .ZN(n79) );
  ND2D1BWP30P140 U5 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U6 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U7 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U8 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U9 ( .A1(n33), .A2(n16), .B1(n41), .B2(n93), .ZN(N295) );
  OAI22D1BWP30P140 U10 ( .A1(n33), .A2(n15), .B1(n41), .B2(n90), .ZN(N296) );
  OAI22D1BWP30P140 U11 ( .A1(n33), .A2(n17), .B1(n41), .B2(n89), .ZN(N297) );
  OAI22D1BWP30P140 U12 ( .A1(n33), .A2(n14), .B1(n41), .B2(n88), .ZN(N298) );
  OAI22D1BWP30P140 U13 ( .A1(n33), .A2(n13), .B1(n41), .B2(n87), .ZN(N299) );
  OAI22D1BWP30P140 U14 ( .A1(n33), .A2(n12), .B1(n41), .B2(n86), .ZN(N300) );
  OAI22D1BWP30P140 U15 ( .A1(n33), .A2(n11), .B1(n41), .B2(n85), .ZN(N301) );
  OAI22D1BWP30P140 U16 ( .A1(n33), .A2(n10), .B1(n41), .B2(n84), .ZN(N302) );
  OAI22D1BWP30P140 U17 ( .A1(n33), .A2(n9), .B1(n41), .B2(n83), .ZN(N303) );
  OAI22D1BWP30P140 U18 ( .A1(n33), .A2(n8), .B1(n41), .B2(n82), .ZN(N304) );
  OAI22D1BWP30P140 U19 ( .A1(n33), .A2(n7), .B1(n41), .B2(n81), .ZN(N305) );
  OAI22D1BWP30P140 U20 ( .A1(n30), .A2(n29), .B1(n31), .B2(n78), .ZN(N307) );
  OAI22D1BWP30P140 U21 ( .A1(n30), .A2(n28), .B1(n31), .B2(n76), .ZN(N308) );
  OAI22D1BWP30P140 U22 ( .A1(n30), .A2(n27), .B1(n31), .B2(n75), .ZN(N309) );
  OAI22D1BWP30P140 U23 ( .A1(n30), .A2(n26), .B1(n31), .B2(n74), .ZN(N310) );
  OAI22D1BWP30P140 U24 ( .A1(n30), .A2(n25), .B1(n31), .B2(n73), .ZN(N311) );
  OAI22D1BWP30P140 U25 ( .A1(n30), .A2(n24), .B1(n31), .B2(n72), .ZN(N312) );
  OAI22D1BWP30P140 U26 ( .A1(n30), .A2(n23), .B1(n31), .B2(n71), .ZN(N313) );
  OAI22D1BWP30P140 U27 ( .A1(n30), .A2(n22), .B1(n31), .B2(n70), .ZN(N314) );
  OAI22D1BWP30P140 U28 ( .A1(n30), .A2(n21), .B1(n31), .B2(n69), .ZN(N315) );
  OAI22D1BWP30P140 U29 ( .A1(n30), .A2(n20), .B1(n31), .B2(n68), .ZN(N316) );
  OAI22D1BWP30P140 U30 ( .A1(n30), .A2(n19), .B1(n31), .B2(n67), .ZN(N317) );
  OAI22D1BWP30P140 U31 ( .A1(n30), .A2(n18), .B1(n31), .B2(n66), .ZN(N318) );
  CKND2D2BWP30P140 U32 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U34 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U35 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U36 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U37 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U38 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U39 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U40 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[50]), .ZN(n7) );
  INR2D1BWP30P140 U42 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U43 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U44 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U45 ( .I(n34), .ZN(n41) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[18]), .ZN(n81) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[49]), .ZN(n8) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[17]), .ZN(n82) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[48]), .ZN(n9) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[16]), .ZN(n83) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[47]), .ZN(n10) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[15]), .ZN(n84) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[46]), .ZN(n11) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[14]), .ZN(n85) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[13]), .ZN(n86) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[44]), .ZN(n13) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[12]), .ZN(n87) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[43]), .ZN(n14) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[11]), .ZN(n88) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[41]), .ZN(n15) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[9]), .ZN(n90) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[40]), .ZN(n16) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[8]), .ZN(n93) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[42]), .ZN(n17) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[10]), .ZN(n89) );
  INVD2BWP30P140 U67 ( .I(n36), .ZN(n30) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[63]), .ZN(n18) );
  INVD2BWP30P140 U69 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[31]), .ZN(n66) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[62]), .ZN(n19) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[30]), .ZN(n67) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[61]), .ZN(n20) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[29]), .ZN(n68) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[60]), .ZN(n21) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[28]), .ZN(n69) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[59]), .ZN(n22) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[27]), .ZN(n70) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[58]), .ZN(n23) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[26]), .ZN(n71) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[25]), .ZN(n72) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[56]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[24]), .ZN(n73) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[55]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[23]), .ZN(n74) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[54]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[22]), .ZN(n75) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[53]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[21]), .ZN(n76) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[52]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[20]), .ZN(n78) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[51]), .ZN(n32) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[19]), .ZN(n80) );
  INVD1BWP30P140 U95 ( .I(n34), .ZN(n47) );
  OAI31D1BWP30P140 U96 ( .A1(n52), .A2(n53), .A3(n35), .B(n47), .ZN(N353) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[6]), .ZN(n64) );
  INVD2BWP30P140 U98 ( .I(n36), .ZN(n46) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U100 ( .A1(n41), .A2(n64), .B1(n46), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[7]), .ZN(n65) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[39]), .ZN(n38) );
  OAI22D1BWP30P140 U103 ( .A1(n41), .A2(n65), .B1(n46), .B2(n38), .ZN(N294) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[5]), .ZN(n63) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[37]), .ZN(n39) );
  OAI22D1BWP30P140 U106 ( .A1(n41), .A2(n63), .B1(n46), .B2(n39), .ZN(N292) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[36]), .ZN(n40) );
  OAI22D1BWP30P140 U109 ( .A1(n41), .A2(n62), .B1(n46), .B2(n40), .ZN(N291) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[35]), .ZN(n42) );
  OAI22D1BWP30P140 U112 ( .A1(n47), .A2(n61), .B1(n46), .B2(n42), .ZN(N290) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[34]), .ZN(n43) );
  OAI22D1BWP30P140 U115 ( .A1(n47), .A2(n60), .B1(n46), .B2(n43), .ZN(N289) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[33]), .ZN(n44) );
  OAI22D1BWP30P140 U118 ( .A1(n47), .A2(n59), .B1(n46), .B2(n44), .ZN(N288) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[0]), .ZN(n58) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[32]), .ZN(n45) );
  OAI22D1BWP30P140 U121 ( .A1(n47), .A2(n58), .B1(n46), .B2(n45), .ZN(N287) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  INVD2BWP30P140 U136 ( .I(n79), .ZN(n77) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n77), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n77), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n77), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n77), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n77), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n77), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n77), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n77), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n77), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n77), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n77), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n77), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  INVD2BWP30P140 U149 ( .I(n79), .ZN(n92) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n92), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_99 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD1BWP30P140 U3 ( .I(n57), .ZN(n67) );
  OAI22D1BWP30P140 U4 ( .A1(n28), .A2(n27), .B1(n31), .B2(n81), .ZN(N306) );
  INVD2BWP30P140 U5 ( .I(n67), .ZN(n79) );
  NR2D1BWP30P140 U6 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  OAI22D1BWP30P140 U7 ( .A1(n33), .A2(n29), .B1(n31), .B2(n80), .ZN(N307) );
  OAI22D1BWP30P140 U8 ( .A1(n33), .A2(n30), .B1(n31), .B2(n78), .ZN(N308) );
  OAI22D1BWP30P140 U9 ( .A1(n33), .A2(n32), .B1(n31), .B2(n77), .ZN(N309) );
  OAI22D1BWP30P140 U10 ( .A1(n33), .A2(n21), .B1(n31), .B2(n76), .ZN(N310) );
  OAI22D1BWP30P140 U11 ( .A1(n33), .A2(n20), .B1(n31), .B2(n75), .ZN(N311) );
  OAI22D1BWP30P140 U12 ( .A1(n33), .A2(n19), .B1(n31), .B2(n74), .ZN(N312) );
  OAI22D1BWP30P140 U13 ( .A1(n33), .A2(n18), .B1(n31), .B2(n73), .ZN(N313) );
  OAI22D1BWP30P140 U14 ( .A1(n33), .A2(n26), .B1(n31), .B2(n72), .ZN(N314) );
  OAI22D1BWP30P140 U15 ( .A1(n33), .A2(n22), .B1(n31), .B2(n71), .ZN(N315) );
  OAI22D1BWP30P140 U16 ( .A1(n33), .A2(n25), .B1(n31), .B2(n70), .ZN(N316) );
  OAI22D1BWP30P140 U17 ( .A1(n33), .A2(n24), .B1(n31), .B2(n69), .ZN(N317) );
  OAI22D1BWP30P140 U18 ( .A1(n33), .A2(n23), .B1(n31), .B2(n68), .ZN(N318) );
  ND2D1BWP30P140 U19 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U20 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U21 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U22 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U23 ( .A1(n28), .A2(n10), .B1(n47), .B2(n66), .ZN(N295) );
  OAI22D1BWP30P140 U24 ( .A1(n28), .A2(n13), .B1(n47), .B2(n93), .ZN(N296) );
  OAI22D1BWP30P140 U25 ( .A1(n28), .A2(n7), .B1(n47), .B2(n90), .ZN(N297) );
  OAI22D1BWP30P140 U26 ( .A1(n28), .A2(n8), .B1(n47), .B2(n89), .ZN(N298) );
  OAI22D1BWP30P140 U27 ( .A1(n28), .A2(n11), .B1(n47), .B2(n88), .ZN(N299) );
  OAI22D1BWP30P140 U28 ( .A1(n28), .A2(n16), .B1(n47), .B2(n87), .ZN(N300) );
  OAI22D1BWP30P140 U29 ( .A1(n28), .A2(n12), .B1(n47), .B2(n86), .ZN(N301) );
  OAI22D1BWP30P140 U30 ( .A1(n28), .A2(n17), .B1(n47), .B2(n85), .ZN(N302) );
  OAI22D1BWP30P140 U31 ( .A1(n28), .A2(n14), .B1(n47), .B2(n84), .ZN(N303) );
  OAI22D1BWP30P140 U32 ( .A1(n28), .A2(n15), .B1(n47), .B2(n83), .ZN(N304) );
  OAI22D1BWP30P140 U33 ( .A1(n28), .A2(n9), .B1(n47), .B2(n82), .ZN(N305) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n28) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[42]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n47) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[10]), .ZN(n90) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[43]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[11]), .ZN(n89) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[50]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[18]), .ZN(n82) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[40]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n88) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[46]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[14]), .ZN(n86) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[41]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[9]), .ZN(n93) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[16]), .ZN(n84) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[17]), .ZN(n83) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[45]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[13]), .ZN(n87) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[47]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[15]), .ZN(n85) );
  INVD2BWP30P140 U69 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[58]), .ZN(n18) );
  INVD2BWP30P140 U71 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[26]), .ZN(n73) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[57]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[25]), .ZN(n74) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[56]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[24]), .ZN(n75) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[55]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[23]), .ZN(n76) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[60]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[28]), .ZN(n71) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[63]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[31]), .ZN(n68) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[62]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[30]), .ZN(n69) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[61]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[29]), .ZN(n70) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n72) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[51]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[19]), .ZN(n81) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[52]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[53]), .ZN(n30) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[21]), .ZN(n78) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[54]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[22]), .ZN(n77) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n41) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n41), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[0]), .ZN(n58) );
  INVD2BWP30P140 U100 ( .I(n36), .ZN(n46) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[32]), .ZN(n37) );
  OAI22D1BWP30P140 U102 ( .A1(n41), .A2(n58), .B1(n46), .B2(n37), .ZN(N287) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[33]), .ZN(n38) );
  OAI22D1BWP30P140 U105 ( .A1(n41), .A2(n59), .B1(n46), .B2(n38), .ZN(N288) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[34]), .ZN(n39) );
  OAI22D1BWP30P140 U108 ( .A1(n41), .A2(n60), .B1(n46), .B2(n39), .ZN(N289) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[35]), .ZN(n40) );
  OAI22D1BWP30P140 U111 ( .A1(n41), .A2(n61), .B1(n46), .B2(n40), .ZN(N290) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[36]), .ZN(n42) );
  OAI22D1BWP30P140 U114 ( .A1(n47), .A2(n62), .B1(n46), .B2(n42), .ZN(N291) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[5]), .ZN(n63) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[37]), .ZN(n43) );
  OAI22D1BWP30P140 U117 ( .A1(n47), .A2(n63), .B1(n46), .B2(n43), .ZN(N292) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[6]), .ZN(n64) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[38]), .ZN(n44) );
  OAI22D1BWP30P140 U120 ( .A1(n47), .A2(n64), .B1(n46), .B2(n44), .ZN(N293) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[7]), .ZN(n65) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[39]), .ZN(n45) );
  OAI22D1BWP30P140 U123 ( .A1(n47), .A2(n65), .B1(n46), .B2(n45), .ZN(N294) );
  INVD1BWP30P140 U124 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U125 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U127 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  MUX2NUD1BWP30P140 U128 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  INVD2BWP30P140 U137 ( .I(n67), .ZN(n92) );
  MOAI22D1BWP30P140 U138 ( .A1(n66), .A2(n92), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n79), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n79), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n79), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n79), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n79), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n79), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n79), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n79), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n79), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n79), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n79), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n79), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_100 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n33), .A2(n32), .B1(n31), .B2(n67), .ZN(N306) );
  INVD1BWP30P140 U4 ( .I(n57), .ZN(n70) );
  ND2D1BWP30P140 U5 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U6 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U7 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U8 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U9 ( .A1(n33), .A2(n17), .B1(n41), .B2(n87), .ZN(N295) );
  OAI22D1BWP30P140 U10 ( .A1(n33), .A2(n16), .B1(n41), .B2(n88), .ZN(N296) );
  OAI22D1BWP30P140 U11 ( .A1(n33), .A2(n15), .B1(n41), .B2(n89), .ZN(N297) );
  OAI22D1BWP30P140 U12 ( .A1(n33), .A2(n14), .B1(n41), .B2(n90), .ZN(N298) );
  OAI22D1BWP30P140 U13 ( .A1(n33), .A2(n13), .B1(n41), .B2(n93), .ZN(N299) );
  OAI22D1BWP30P140 U14 ( .A1(n33), .A2(n12), .B1(n41), .B2(n86), .ZN(N300) );
  OAI22D1BWP30P140 U15 ( .A1(n33), .A2(n11), .B1(n41), .B2(n85), .ZN(N301) );
  OAI22D1BWP30P140 U16 ( .A1(n33), .A2(n10), .B1(n41), .B2(n69), .ZN(N302) );
  OAI22D1BWP30P140 U17 ( .A1(n33), .A2(n9), .B1(n41), .B2(n68), .ZN(N303) );
  OAI22D1BWP30P140 U18 ( .A1(n33), .A2(n8), .B1(n41), .B2(n66), .ZN(N304) );
  OAI22D1BWP30P140 U19 ( .A1(n33), .A2(n7), .B1(n41), .B2(n73), .ZN(N305) );
  OAI22D1BWP30P140 U20 ( .A1(n30), .A2(n29), .B1(n31), .B2(n71), .ZN(N307) );
  OAI22D1BWP30P140 U21 ( .A1(n30), .A2(n28), .B1(n31), .B2(n72), .ZN(N308) );
  OAI22D1BWP30P140 U22 ( .A1(n30), .A2(n27), .B1(n31), .B2(n74), .ZN(N309) );
  OAI22D1BWP30P140 U23 ( .A1(n30), .A2(n26), .B1(n31), .B2(n75), .ZN(N310) );
  OAI22D1BWP30P140 U24 ( .A1(n30), .A2(n25), .B1(n31), .B2(n76), .ZN(N311) );
  OAI22D1BWP30P140 U25 ( .A1(n30), .A2(n24), .B1(n31), .B2(n77), .ZN(N312) );
  OAI22D1BWP30P140 U26 ( .A1(n30), .A2(n23), .B1(n31), .B2(n78), .ZN(N313) );
  OAI22D1BWP30P140 U27 ( .A1(n30), .A2(n22), .B1(n31), .B2(n79), .ZN(N314) );
  OAI22D1BWP30P140 U28 ( .A1(n30), .A2(n21), .B1(n31), .B2(n80), .ZN(N315) );
  OAI22D1BWP30P140 U29 ( .A1(n30), .A2(n20), .B1(n31), .B2(n81), .ZN(N316) );
  OAI22D1BWP30P140 U30 ( .A1(n30), .A2(n19), .B1(n31), .B2(n82), .ZN(N317) );
  OAI22D1BWP30P140 U31 ( .A1(n30), .A2(n18), .B1(n31), .B2(n84), .ZN(N318) );
  CKND2D2BWP30P140 U32 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U34 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U35 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U36 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U37 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U38 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U39 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U40 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[50]), .ZN(n7) );
  INR2D1BWP30P140 U42 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U43 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U44 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U45 ( .I(n34), .ZN(n41) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[18]), .ZN(n73) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[49]), .ZN(n8) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[17]), .ZN(n66) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[48]), .ZN(n9) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[16]), .ZN(n68) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[47]), .ZN(n10) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[15]), .ZN(n69) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[46]), .ZN(n11) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[14]), .ZN(n85) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[13]), .ZN(n86) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[44]), .ZN(n13) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[12]), .ZN(n93) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[43]), .ZN(n14) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[11]), .ZN(n90) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[42]), .ZN(n15) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[10]), .ZN(n89) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[41]), .ZN(n16) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[9]), .ZN(n88) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[40]), .ZN(n17) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[8]), .ZN(n87) );
  INVD2BWP30P140 U67 ( .I(n36), .ZN(n30) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[63]), .ZN(n18) );
  INVD2BWP30P140 U69 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[31]), .ZN(n84) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[62]), .ZN(n19) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[30]), .ZN(n82) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[61]), .ZN(n20) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[29]), .ZN(n81) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[60]), .ZN(n21) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[28]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[59]), .ZN(n22) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[27]), .ZN(n79) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[58]), .ZN(n23) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[26]), .ZN(n78) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[25]), .ZN(n77) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[56]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[24]), .ZN(n76) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[55]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[23]), .ZN(n75) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[54]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[22]), .ZN(n74) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[53]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[21]), .ZN(n72) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[52]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[20]), .ZN(n71) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[51]), .ZN(n32) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[19]), .ZN(n67) );
  INVD1BWP30P140 U95 ( .I(n34), .ZN(n47) );
  OAI31D1BWP30P140 U96 ( .A1(n52), .A2(n53), .A3(n35), .B(n47), .ZN(N353) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[7]), .ZN(n65) );
  INVD2BWP30P140 U98 ( .I(n36), .ZN(n46) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[39]), .ZN(n37) );
  OAI22D1BWP30P140 U100 ( .A1(n41), .A2(n65), .B1(n46), .B2(n37), .ZN(N294) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[6]), .ZN(n64) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[38]), .ZN(n38) );
  OAI22D1BWP30P140 U103 ( .A1(n41), .A2(n64), .B1(n46), .B2(n38), .ZN(N293) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[5]), .ZN(n63) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[37]), .ZN(n39) );
  OAI22D1BWP30P140 U106 ( .A1(n41), .A2(n63), .B1(n46), .B2(n39), .ZN(N292) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[36]), .ZN(n40) );
  OAI22D1BWP30P140 U109 ( .A1(n41), .A2(n62), .B1(n46), .B2(n40), .ZN(N291) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[33]), .ZN(n42) );
  OAI22D1BWP30P140 U112 ( .A1(n47), .A2(n59), .B1(n46), .B2(n42), .ZN(N288) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[35]), .ZN(n43) );
  OAI22D1BWP30P140 U115 ( .A1(n47), .A2(n61), .B1(n46), .B2(n43), .ZN(N290) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[0]), .ZN(n58) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U118 ( .A1(n47), .A2(n58), .B1(n46), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[34]), .ZN(n45) );
  OAI22D1BWP30P140 U121 ( .A1(n47), .A2(n60), .B1(n46), .B2(n45), .ZN(N289) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  INVD2BWP30P140 U136 ( .I(n70), .ZN(n92) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n92), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n92), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n92), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n92), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  INVD2BWP30P140 U141 ( .I(n70), .ZN(n83) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n83), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n83), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n92), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n83), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n83), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n83), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n83), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n83), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n83), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n83), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n83), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n83), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n83), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_101 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n33), .A2(n32), .B1(n31), .B2(n78), .ZN(N306) );
  INVD1BWP30P140 U4 ( .I(n57), .ZN(n79) );
  ND2D1BWP30P140 U5 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U6 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U7 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U8 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U9 ( .A1(n33), .A2(n17), .B1(n41), .B2(n66), .ZN(N295) );
  OAI22D1BWP30P140 U10 ( .A1(n33), .A2(n16), .B1(n41), .B2(n67), .ZN(N296) );
  OAI22D1BWP30P140 U11 ( .A1(n33), .A2(n15), .B1(n41), .B2(n68), .ZN(N297) );
  OAI22D1BWP30P140 U12 ( .A1(n33), .A2(n14), .B1(n41), .B2(n69), .ZN(N298) );
  OAI22D1BWP30P140 U13 ( .A1(n33), .A2(n13), .B1(n41), .B2(n70), .ZN(N299) );
  OAI22D1BWP30P140 U14 ( .A1(n33), .A2(n12), .B1(n41), .B2(n71), .ZN(N300) );
  OAI22D1BWP30P140 U15 ( .A1(n33), .A2(n11), .B1(n41), .B2(n72), .ZN(N301) );
  OAI22D1BWP30P140 U16 ( .A1(n33), .A2(n10), .B1(n41), .B2(n73), .ZN(N302) );
  OAI22D1BWP30P140 U17 ( .A1(n33), .A2(n9), .B1(n41), .B2(n74), .ZN(N303) );
  OAI22D1BWP30P140 U18 ( .A1(n33), .A2(n8), .B1(n41), .B2(n75), .ZN(N304) );
  OAI22D1BWP30P140 U19 ( .A1(n33), .A2(n7), .B1(n41), .B2(n76), .ZN(N305) );
  OAI22D1BWP30P140 U20 ( .A1(n30), .A2(n29), .B1(n31), .B2(n80), .ZN(N307) );
  OAI22D1BWP30P140 U21 ( .A1(n30), .A2(n28), .B1(n31), .B2(n81), .ZN(N308) );
  OAI22D1BWP30P140 U22 ( .A1(n30), .A2(n27), .B1(n31), .B2(n82), .ZN(N309) );
  OAI22D1BWP30P140 U23 ( .A1(n30), .A2(n26), .B1(n31), .B2(n83), .ZN(N310) );
  OAI22D1BWP30P140 U24 ( .A1(n30), .A2(n25), .B1(n31), .B2(n84), .ZN(N311) );
  OAI22D1BWP30P140 U25 ( .A1(n30), .A2(n24), .B1(n31), .B2(n85), .ZN(N312) );
  OAI22D1BWP30P140 U26 ( .A1(n30), .A2(n23), .B1(n31), .B2(n86), .ZN(N313) );
  OAI22D1BWP30P140 U27 ( .A1(n30), .A2(n22), .B1(n31), .B2(n87), .ZN(N314) );
  OAI22D1BWP30P140 U28 ( .A1(n30), .A2(n21), .B1(n31), .B2(n88), .ZN(N315) );
  OAI22D1BWP30P140 U29 ( .A1(n30), .A2(n20), .B1(n31), .B2(n89), .ZN(N316) );
  OAI22D1BWP30P140 U30 ( .A1(n30), .A2(n19), .B1(n31), .B2(n90), .ZN(N317) );
  OAI22D1BWP30P140 U31 ( .A1(n30), .A2(n18), .B1(n31), .B2(n93), .ZN(N318) );
  CKND2D2BWP30P140 U32 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U34 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U35 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U36 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U37 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U38 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U39 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U40 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[50]), .ZN(n7) );
  INR2D1BWP30P140 U42 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U43 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U44 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U45 ( .I(n34), .ZN(n41) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[18]), .ZN(n76) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[49]), .ZN(n8) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[17]), .ZN(n75) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[48]), .ZN(n9) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[16]), .ZN(n74) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[47]), .ZN(n10) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[15]), .ZN(n73) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[46]), .ZN(n11) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[14]), .ZN(n72) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[13]), .ZN(n71) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[44]), .ZN(n13) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[12]), .ZN(n70) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[43]), .ZN(n14) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[42]), .ZN(n15) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[10]), .ZN(n68) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[41]), .ZN(n16) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[9]), .ZN(n67) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[40]), .ZN(n17) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD2BWP30P140 U67 ( .I(n36), .ZN(n30) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[63]), .ZN(n18) );
  INVD2BWP30P140 U69 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[31]), .ZN(n93) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[62]), .ZN(n19) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[30]), .ZN(n90) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[61]), .ZN(n20) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[29]), .ZN(n89) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[60]), .ZN(n21) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[28]), .ZN(n88) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[59]), .ZN(n22) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[27]), .ZN(n87) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[58]), .ZN(n23) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[26]), .ZN(n86) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[25]), .ZN(n85) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[56]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[24]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[55]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[23]), .ZN(n83) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[54]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[22]), .ZN(n82) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[53]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[21]), .ZN(n81) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[52]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[51]), .ZN(n32) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD1BWP30P140 U95 ( .I(n34), .ZN(n47) );
  OAI31D1BWP30P140 U96 ( .A1(n52), .A2(n53), .A3(n35), .B(n47), .ZN(N353) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[7]), .ZN(n65) );
  INVD2BWP30P140 U98 ( .I(n36), .ZN(n46) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[39]), .ZN(n37) );
  OAI22D1BWP30P140 U100 ( .A1(n41), .A2(n65), .B1(n46), .B2(n37), .ZN(N294) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[6]), .ZN(n64) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[38]), .ZN(n38) );
  OAI22D1BWP30P140 U103 ( .A1(n41), .A2(n64), .B1(n46), .B2(n38), .ZN(N293) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[5]), .ZN(n63) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[37]), .ZN(n39) );
  OAI22D1BWP30P140 U106 ( .A1(n41), .A2(n63), .B1(n46), .B2(n39), .ZN(N292) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[36]), .ZN(n40) );
  OAI22D1BWP30P140 U109 ( .A1(n41), .A2(n62), .B1(n46), .B2(n40), .ZN(N291) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[35]), .ZN(n42) );
  OAI22D1BWP30P140 U112 ( .A1(n47), .A2(n61), .B1(n46), .B2(n42), .ZN(N290) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[34]), .ZN(n43) );
  OAI22D1BWP30P140 U115 ( .A1(n47), .A2(n60), .B1(n46), .B2(n43), .ZN(N289) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[33]), .ZN(n44) );
  OAI22D1BWP30P140 U118 ( .A1(n47), .A2(n59), .B1(n46), .B2(n44), .ZN(N288) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[0]), .ZN(n58) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[32]), .ZN(n45) );
  OAI22D1BWP30P140 U121 ( .A1(n47), .A2(n58), .B1(n46), .B2(n45), .ZN(N287) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  INVD2BWP30P140 U136 ( .I(n79), .ZN(n77) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n77), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n77), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n77), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n77), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n77), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n77), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n77), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n77), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n77), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n77), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n77), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n77), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  INVD2BWP30P140 U149 ( .I(n79), .ZN(n92) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n92), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_102 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  OAI22D1BWP30P140 U3 ( .A1(n33), .A2(n32), .B1(n31), .B2(n78), .ZN(N306) );
  INVD1BWP30P140 U4 ( .I(n57), .ZN(n79) );
  ND2D1BWP30P140 U5 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U6 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U7 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U8 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U9 ( .A1(n33), .A2(n17), .B1(n43), .B2(n66), .ZN(N295) );
  OAI22D1BWP30P140 U10 ( .A1(n33), .A2(n16), .B1(n43), .B2(n67), .ZN(N296) );
  OAI22D1BWP30P140 U11 ( .A1(n33), .A2(n15), .B1(n43), .B2(n68), .ZN(N297) );
  OAI22D1BWP30P140 U12 ( .A1(n33), .A2(n14), .B1(n43), .B2(n69), .ZN(N298) );
  OAI22D1BWP30P140 U13 ( .A1(n33), .A2(n13), .B1(n43), .B2(n70), .ZN(N299) );
  OAI22D1BWP30P140 U14 ( .A1(n33), .A2(n12), .B1(n43), .B2(n71), .ZN(N300) );
  OAI22D1BWP30P140 U15 ( .A1(n33), .A2(n11), .B1(n43), .B2(n72), .ZN(N301) );
  OAI22D1BWP30P140 U16 ( .A1(n33), .A2(n10), .B1(n43), .B2(n73), .ZN(N302) );
  OAI22D1BWP30P140 U17 ( .A1(n33), .A2(n9), .B1(n43), .B2(n74), .ZN(N303) );
  OAI22D1BWP30P140 U18 ( .A1(n33), .A2(n8), .B1(n43), .B2(n75), .ZN(N304) );
  OAI22D1BWP30P140 U19 ( .A1(n33), .A2(n7), .B1(n43), .B2(n76), .ZN(N305) );
  OAI22D1BWP30P140 U20 ( .A1(n30), .A2(n29), .B1(n31), .B2(n80), .ZN(N307) );
  OAI22D1BWP30P140 U21 ( .A1(n30), .A2(n28), .B1(n31), .B2(n81), .ZN(N308) );
  OAI22D1BWP30P140 U22 ( .A1(n30), .A2(n27), .B1(n31), .B2(n82), .ZN(N309) );
  OAI22D1BWP30P140 U23 ( .A1(n30), .A2(n26), .B1(n31), .B2(n83), .ZN(N310) );
  OAI22D1BWP30P140 U24 ( .A1(n30), .A2(n25), .B1(n31), .B2(n84), .ZN(N311) );
  OAI22D1BWP30P140 U25 ( .A1(n30), .A2(n24), .B1(n31), .B2(n85), .ZN(N312) );
  OAI22D1BWP30P140 U26 ( .A1(n30), .A2(n23), .B1(n31), .B2(n86), .ZN(N313) );
  OAI22D1BWP30P140 U27 ( .A1(n30), .A2(n22), .B1(n31), .B2(n87), .ZN(N314) );
  OAI22D1BWP30P140 U28 ( .A1(n30), .A2(n21), .B1(n31), .B2(n88), .ZN(N315) );
  OAI22D1BWP30P140 U29 ( .A1(n30), .A2(n20), .B1(n31), .B2(n89), .ZN(N316) );
  OAI22D1BWP30P140 U30 ( .A1(n30), .A2(n19), .B1(n31), .B2(n90), .ZN(N317) );
  OAI22D1BWP30P140 U31 ( .A1(n30), .A2(n18), .B1(n31), .B2(n93), .ZN(N318) );
  CKND2D2BWP30P140 U32 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U34 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U35 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U36 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U37 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U38 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U39 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U40 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[50]), .ZN(n7) );
  INR2D1BWP30P140 U42 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U43 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U44 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U45 ( .I(n34), .ZN(n43) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[18]), .ZN(n76) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[49]), .ZN(n8) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[17]), .ZN(n75) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[48]), .ZN(n9) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[16]), .ZN(n74) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[47]), .ZN(n10) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[15]), .ZN(n73) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[46]), .ZN(n11) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[14]), .ZN(n72) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[13]), .ZN(n71) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[44]), .ZN(n13) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[12]), .ZN(n70) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[43]), .ZN(n14) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[42]), .ZN(n15) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[10]), .ZN(n68) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[41]), .ZN(n16) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[9]), .ZN(n67) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[40]), .ZN(n17) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD2BWP30P140 U67 ( .I(n36), .ZN(n30) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[63]), .ZN(n18) );
  INVD2BWP30P140 U69 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[31]), .ZN(n93) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[62]), .ZN(n19) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[30]), .ZN(n90) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[61]), .ZN(n20) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[29]), .ZN(n89) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[60]), .ZN(n21) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[28]), .ZN(n88) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[59]), .ZN(n22) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[27]), .ZN(n87) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[58]), .ZN(n23) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[26]), .ZN(n86) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[25]), .ZN(n85) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[56]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[24]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[55]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[23]), .ZN(n83) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[54]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[22]), .ZN(n82) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[53]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[21]), .ZN(n81) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[52]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[51]), .ZN(n32) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD1BWP30P140 U95 ( .I(n34), .ZN(n47) );
  OAI31D1BWP30P140 U96 ( .A1(n52), .A2(n53), .A3(n35), .B(n47), .ZN(N353) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD2BWP30P140 U98 ( .I(n36), .ZN(n46) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[33]), .ZN(n37) );
  OAI22D1BWP30P140 U100 ( .A1(n47), .A2(n59), .B1(n46), .B2(n37), .ZN(N288) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[35]), .ZN(n38) );
  OAI22D1BWP30P140 U103 ( .A1(n47), .A2(n61), .B1(n46), .B2(n38), .ZN(N290) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U106 ( .A1(n43), .A2(n62), .B1(n46), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[5]), .ZN(n63) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[37]), .ZN(n40) );
  OAI22D1BWP30P140 U109 ( .A1(n43), .A2(n63), .B1(n46), .B2(n40), .ZN(N292) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[6]), .ZN(n64) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[38]), .ZN(n41) );
  OAI22D1BWP30P140 U112 ( .A1(n43), .A2(n64), .B1(n46), .B2(n41), .ZN(N293) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[7]), .ZN(n65) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[39]), .ZN(n42) );
  OAI22D1BWP30P140 U115 ( .A1(n43), .A2(n65), .B1(n46), .B2(n42), .ZN(N294) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[34]), .ZN(n44) );
  OAI22D1BWP30P140 U118 ( .A1(n47), .A2(n60), .B1(n46), .B2(n44), .ZN(N289) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[0]), .ZN(n58) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[32]), .ZN(n45) );
  OAI22D1BWP30P140 U121 ( .A1(n47), .A2(n58), .B1(n46), .B2(n45), .ZN(N287) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  INVD2BWP30P140 U136 ( .I(n79), .ZN(n77) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n77), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n77), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n77), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n77), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n77), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n77), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n77), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n77), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n77), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n77), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n77), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n77), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  INVD2BWP30P140 U149 ( .I(n79), .ZN(n92) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n92), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_103 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n33), .A2(n32), .B1(n31), .B2(n78), .ZN(N306) );
  INVD1BWP30P140 U4 ( .I(n57), .ZN(n79) );
  ND2D1BWP30P140 U5 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U6 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U7 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U8 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U9 ( .A1(n33), .A2(n17), .B1(n44), .B2(n66), .ZN(N295) );
  OAI22D1BWP30P140 U10 ( .A1(n33), .A2(n16), .B1(n44), .B2(n67), .ZN(N296) );
  OAI22D1BWP30P140 U11 ( .A1(n33), .A2(n15), .B1(n44), .B2(n68), .ZN(N297) );
  OAI22D1BWP30P140 U12 ( .A1(n33), .A2(n14), .B1(n44), .B2(n69), .ZN(N298) );
  OAI22D1BWP30P140 U13 ( .A1(n33), .A2(n13), .B1(n44), .B2(n70), .ZN(N299) );
  OAI22D1BWP30P140 U14 ( .A1(n33), .A2(n12), .B1(n44), .B2(n71), .ZN(N300) );
  OAI22D1BWP30P140 U15 ( .A1(n33), .A2(n11), .B1(n44), .B2(n72), .ZN(N301) );
  OAI22D1BWP30P140 U16 ( .A1(n33), .A2(n10), .B1(n44), .B2(n73), .ZN(N302) );
  OAI22D1BWP30P140 U17 ( .A1(n33), .A2(n9), .B1(n44), .B2(n74), .ZN(N303) );
  OAI22D1BWP30P140 U18 ( .A1(n33), .A2(n8), .B1(n44), .B2(n75), .ZN(N304) );
  OAI22D1BWP30P140 U19 ( .A1(n33), .A2(n7), .B1(n44), .B2(n76), .ZN(N305) );
  OAI22D1BWP30P140 U20 ( .A1(n30), .A2(n29), .B1(n31), .B2(n80), .ZN(N307) );
  OAI22D1BWP30P140 U21 ( .A1(n30), .A2(n28), .B1(n31), .B2(n81), .ZN(N308) );
  OAI22D1BWP30P140 U22 ( .A1(n30), .A2(n27), .B1(n31), .B2(n82), .ZN(N309) );
  OAI22D1BWP30P140 U23 ( .A1(n30), .A2(n26), .B1(n31), .B2(n83), .ZN(N310) );
  OAI22D1BWP30P140 U24 ( .A1(n30), .A2(n25), .B1(n31), .B2(n84), .ZN(N311) );
  OAI22D1BWP30P140 U25 ( .A1(n30), .A2(n24), .B1(n31), .B2(n85), .ZN(N312) );
  OAI22D1BWP30P140 U26 ( .A1(n30), .A2(n23), .B1(n31), .B2(n86), .ZN(N313) );
  OAI22D1BWP30P140 U27 ( .A1(n30), .A2(n22), .B1(n31), .B2(n87), .ZN(N314) );
  OAI22D1BWP30P140 U28 ( .A1(n30), .A2(n21), .B1(n31), .B2(n88), .ZN(N315) );
  OAI22D1BWP30P140 U29 ( .A1(n30), .A2(n20), .B1(n31), .B2(n89), .ZN(N316) );
  OAI22D1BWP30P140 U30 ( .A1(n30), .A2(n19), .B1(n31), .B2(n90), .ZN(N317) );
  OAI22D1BWP30P140 U31 ( .A1(n30), .A2(n18), .B1(n31), .B2(n93), .ZN(N318) );
  CKND2D2BWP30P140 U32 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U34 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U35 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U36 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U37 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U38 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U39 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U40 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U41 ( .I(i_data_bus[50]), .ZN(n7) );
  INR2D1BWP30P140 U42 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U43 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U44 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U45 ( .I(n34), .ZN(n44) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[18]), .ZN(n76) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[49]), .ZN(n8) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[17]), .ZN(n75) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[48]), .ZN(n9) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[16]), .ZN(n74) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[47]), .ZN(n10) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[15]), .ZN(n73) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[46]), .ZN(n11) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[14]), .ZN(n72) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[13]), .ZN(n71) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[44]), .ZN(n13) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[12]), .ZN(n70) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[43]), .ZN(n14) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[42]), .ZN(n15) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[10]), .ZN(n68) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[41]), .ZN(n16) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[9]), .ZN(n67) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[40]), .ZN(n17) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD2BWP30P140 U67 ( .I(n36), .ZN(n30) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[63]), .ZN(n18) );
  INVD2BWP30P140 U69 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[31]), .ZN(n93) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[62]), .ZN(n19) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[30]), .ZN(n90) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[61]), .ZN(n20) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[29]), .ZN(n89) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[60]), .ZN(n21) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[28]), .ZN(n88) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[59]), .ZN(n22) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[27]), .ZN(n87) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[58]), .ZN(n23) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[26]), .ZN(n86) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[25]), .ZN(n85) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[56]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[24]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[55]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[23]), .ZN(n83) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[54]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[22]), .ZN(n82) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[53]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[21]), .ZN(n81) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[52]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[51]), .ZN(n32) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD1BWP30P140 U95 ( .I(n34), .ZN(n47) );
  OAI31D1BWP30P140 U96 ( .A1(n52), .A2(n53), .A3(n35), .B(n47), .ZN(N353) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD2BWP30P140 U98 ( .I(n36), .ZN(n46) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[33]), .ZN(n37) );
  OAI22D1BWP30P140 U100 ( .A1(n47), .A2(n59), .B1(n46), .B2(n37), .ZN(N288) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[34]), .ZN(n38) );
  OAI22D1BWP30P140 U103 ( .A1(n47), .A2(n60), .B1(n46), .B2(n38), .ZN(N289) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[35]), .ZN(n39) );
  OAI22D1BWP30P140 U106 ( .A1(n47), .A2(n61), .B1(n46), .B2(n39), .ZN(N290) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[36]), .ZN(n40) );
  OAI22D1BWP30P140 U109 ( .A1(n44), .A2(n62), .B1(n46), .B2(n40), .ZN(N291) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[5]), .ZN(n63) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[37]), .ZN(n41) );
  OAI22D1BWP30P140 U112 ( .A1(n44), .A2(n63), .B1(n46), .B2(n41), .ZN(N292) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[6]), .ZN(n64) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[38]), .ZN(n42) );
  OAI22D1BWP30P140 U115 ( .A1(n44), .A2(n64), .B1(n46), .B2(n42), .ZN(N293) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[7]), .ZN(n65) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[39]), .ZN(n43) );
  OAI22D1BWP30P140 U118 ( .A1(n44), .A2(n65), .B1(n46), .B2(n43), .ZN(N294) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[0]), .ZN(n58) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[32]), .ZN(n45) );
  OAI22D1BWP30P140 U121 ( .A1(n47), .A2(n58), .B1(n46), .B2(n45), .ZN(N287) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  INVD2BWP30P140 U136 ( .I(n79), .ZN(n77) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n77), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n77), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n77), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n77), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n77), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n77), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n77), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n77), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n77), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n77), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n77), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n77), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  INVD2BWP30P140 U149 ( .I(n79), .ZN(n92) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n92), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_104 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n33), .A2(n32), .B1(n31), .B2(n78), .ZN(N306) );
  INVD2BWP30P140 U4 ( .I(n36), .ZN(n46) );
  OAI22D1BWP30P140 U5 ( .A1(n47), .A2(n58), .B1(n46), .B2(n45), .ZN(N287) );
  INVD1BWP30P140 U6 ( .I(n57), .ZN(n79) );
  ND2D1BWP30P140 U7 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U9 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U10 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U11 ( .A1(n33), .A2(n17), .B1(n41), .B2(n66), .ZN(N295) );
  OAI22D1BWP30P140 U12 ( .A1(n33), .A2(n16), .B1(n41), .B2(n67), .ZN(N296) );
  OAI22D1BWP30P140 U13 ( .A1(n33), .A2(n15), .B1(n41), .B2(n68), .ZN(N297) );
  OAI22D1BWP30P140 U14 ( .A1(n33), .A2(n14), .B1(n41), .B2(n69), .ZN(N298) );
  OAI22D1BWP30P140 U15 ( .A1(n33), .A2(n13), .B1(n41), .B2(n70), .ZN(N299) );
  OAI22D1BWP30P140 U16 ( .A1(n33), .A2(n12), .B1(n41), .B2(n71), .ZN(N300) );
  OAI22D1BWP30P140 U17 ( .A1(n33), .A2(n11), .B1(n41), .B2(n72), .ZN(N301) );
  OAI22D1BWP30P140 U18 ( .A1(n33), .A2(n10), .B1(n41), .B2(n73), .ZN(N302) );
  OAI22D1BWP30P140 U19 ( .A1(n33), .A2(n9), .B1(n41), .B2(n74), .ZN(N303) );
  OAI22D1BWP30P140 U20 ( .A1(n33), .A2(n8), .B1(n41), .B2(n75), .ZN(N304) );
  OAI22D1BWP30P140 U21 ( .A1(n33), .A2(n7), .B1(n41), .B2(n76), .ZN(N305) );
  OAI22D1BWP30P140 U22 ( .A1(n30), .A2(n29), .B1(n31), .B2(n80), .ZN(N307) );
  OAI22D1BWP30P140 U23 ( .A1(n30), .A2(n28), .B1(n31), .B2(n81), .ZN(N308) );
  OAI22D1BWP30P140 U24 ( .A1(n30), .A2(n27), .B1(n31), .B2(n82), .ZN(N309) );
  OAI22D1BWP30P140 U25 ( .A1(n30), .A2(n26), .B1(n31), .B2(n83), .ZN(N310) );
  OAI22D1BWP30P140 U26 ( .A1(n30), .A2(n25), .B1(n31), .B2(n84), .ZN(N311) );
  OAI22D1BWP30P140 U27 ( .A1(n30), .A2(n24), .B1(n31), .B2(n85), .ZN(N312) );
  OAI22D1BWP30P140 U28 ( .A1(n30), .A2(n23), .B1(n31), .B2(n86), .ZN(N313) );
  OAI22D1BWP30P140 U29 ( .A1(n30), .A2(n22), .B1(n31), .B2(n87), .ZN(N314) );
  OAI22D1BWP30P140 U30 ( .A1(n30), .A2(n21), .B1(n31), .B2(n88), .ZN(N315) );
  OAI22D1BWP30P140 U31 ( .A1(n30), .A2(n20), .B1(n31), .B2(n89), .ZN(N316) );
  OAI22D1BWP30P140 U32 ( .A1(n30), .A2(n19), .B1(n31), .B2(n90), .ZN(N317) );
  OAI22D1BWP30P140 U33 ( .A1(n30), .A2(n18), .B1(n31), .B2(n93), .ZN(N318) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[50]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n41) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[18]), .ZN(n76) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[49]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[17]), .ZN(n75) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[48]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[16]), .ZN(n74) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[47]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[15]), .ZN(n73) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[46]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[14]), .ZN(n72) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n71) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[44]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[12]), .ZN(n70) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[43]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[42]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[10]), .ZN(n68) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[41]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[9]), .ZN(n67) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[40]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD2BWP30P140 U69 ( .I(n36), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[63]), .ZN(n18) );
  INVD2BWP30P140 U71 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[31]), .ZN(n93) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[62]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[30]), .ZN(n90) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[61]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[29]), .ZN(n89) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[60]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[28]), .ZN(n88) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[59]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[27]), .ZN(n87) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[58]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[26]), .ZN(n86) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n85) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[56]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[24]), .ZN(n84) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[55]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[23]), .ZN(n83) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[54]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[22]), .ZN(n82) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[53]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[21]), .ZN(n81) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[52]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[51]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n47) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n47), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n65) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[39]), .ZN(n37) );
  OAI22D1BWP30P140 U101 ( .A1(n41), .A2(n65), .B1(n46), .B2(n37), .ZN(N294) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[6]), .ZN(n64) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[38]), .ZN(n38) );
  OAI22D1BWP30P140 U104 ( .A1(n41), .A2(n64), .B1(n46), .B2(n38), .ZN(N293) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[5]), .ZN(n63) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[37]), .ZN(n39) );
  OAI22D1BWP30P140 U107 ( .A1(n41), .A2(n63), .B1(n46), .B2(n39), .ZN(N292) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[36]), .ZN(n40) );
  OAI22D1BWP30P140 U110 ( .A1(n41), .A2(n62), .B1(n46), .B2(n40), .ZN(N291) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[35]), .ZN(n42) );
  OAI22D1BWP30P140 U113 ( .A1(n47), .A2(n61), .B1(n46), .B2(n42), .ZN(N290) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[34]), .ZN(n43) );
  OAI22D1BWP30P140 U116 ( .A1(n47), .A2(n60), .B1(n46), .B2(n43), .ZN(N289) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[33]), .ZN(n44) );
  OAI22D1BWP30P140 U119 ( .A1(n47), .A2(n59), .B1(n46), .B2(n44), .ZN(N288) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[0]), .ZN(n58) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[32]), .ZN(n45) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  INVD2BWP30P140 U136 ( .I(n79), .ZN(n77) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n77), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n77), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n77), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n77), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n77), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n77), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n77), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n77), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n77), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n77), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n77), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n77), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  INVD2BWP30P140 U149 ( .I(n79), .ZN(n92) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n92), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_105 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD1BWP30P140 U3 ( .I(n57), .ZN(n79) );
  OAI22D1BWP30P140 U4 ( .A1(n33), .A2(n32), .B1(n31), .B2(n78), .ZN(N306) );
  INVD2BWP30P140 U5 ( .I(n79), .ZN(n92) );
  NR2D1BWP30P140 U6 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  OAI22D1BWP30P140 U7 ( .A1(n33), .A2(n17), .B1(n42), .B2(n66), .ZN(N295) );
  OAI22D1BWP30P140 U8 ( .A1(n33), .A2(n16), .B1(n42), .B2(n67), .ZN(N296) );
  OAI22D1BWP30P140 U9 ( .A1(n33), .A2(n15), .B1(n42), .B2(n68), .ZN(N297) );
  OAI22D1BWP30P140 U10 ( .A1(n33), .A2(n14), .B1(n42), .B2(n69), .ZN(N298) );
  OAI22D1BWP30P140 U11 ( .A1(n33), .A2(n13), .B1(n42), .B2(n70), .ZN(N299) );
  OAI22D1BWP30P140 U12 ( .A1(n33), .A2(n12), .B1(n42), .B2(n71), .ZN(N300) );
  OAI22D1BWP30P140 U13 ( .A1(n33), .A2(n11), .B1(n42), .B2(n72), .ZN(N301) );
  OAI22D1BWP30P140 U14 ( .A1(n33), .A2(n10), .B1(n42), .B2(n73), .ZN(N302) );
  OAI22D1BWP30P140 U15 ( .A1(n33), .A2(n9), .B1(n42), .B2(n74), .ZN(N303) );
  OAI22D1BWP30P140 U16 ( .A1(n33), .A2(n8), .B1(n42), .B2(n75), .ZN(N304) );
  OAI22D1BWP30P140 U17 ( .A1(n33), .A2(n7), .B1(n42), .B2(n76), .ZN(N305) );
  ND2D1BWP30P140 U18 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U19 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U20 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U21 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U22 ( .A1(n30), .A2(n29), .B1(n31), .B2(n80), .ZN(N307) );
  OAI22D1BWP30P140 U23 ( .A1(n30), .A2(n28), .B1(n31), .B2(n81), .ZN(N308) );
  OAI22D1BWP30P140 U24 ( .A1(n30), .A2(n27), .B1(n31), .B2(n82), .ZN(N309) );
  OAI22D1BWP30P140 U25 ( .A1(n30), .A2(n26), .B1(n31), .B2(n83), .ZN(N310) );
  OAI22D1BWP30P140 U26 ( .A1(n30), .A2(n25), .B1(n31), .B2(n84), .ZN(N311) );
  OAI22D1BWP30P140 U27 ( .A1(n30), .A2(n24), .B1(n31), .B2(n85), .ZN(N312) );
  OAI22D1BWP30P140 U28 ( .A1(n30), .A2(n23), .B1(n31), .B2(n86), .ZN(N313) );
  OAI22D1BWP30P140 U29 ( .A1(n30), .A2(n22), .B1(n31), .B2(n87), .ZN(N314) );
  OAI22D1BWP30P140 U30 ( .A1(n30), .A2(n21), .B1(n31), .B2(n88), .ZN(N315) );
  OAI22D1BWP30P140 U31 ( .A1(n30), .A2(n20), .B1(n31), .B2(n89), .ZN(N316) );
  OAI22D1BWP30P140 U32 ( .A1(n30), .A2(n19), .B1(n31), .B2(n90), .ZN(N317) );
  OAI22D1BWP30P140 U33 ( .A1(n30), .A2(n18), .B1(n31), .B2(n93), .ZN(N318) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[50]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n42) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[18]), .ZN(n76) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[49]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[17]), .ZN(n75) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[48]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[16]), .ZN(n74) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[47]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[15]), .ZN(n73) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[46]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[14]), .ZN(n72) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n71) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[44]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[12]), .ZN(n70) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[43]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[42]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[10]), .ZN(n68) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[41]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[9]), .ZN(n67) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[40]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD2BWP30P140 U69 ( .I(n36), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[63]), .ZN(n18) );
  INVD2BWP30P140 U71 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[31]), .ZN(n93) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[62]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[30]), .ZN(n90) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[61]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[29]), .ZN(n89) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[60]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[28]), .ZN(n88) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[59]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[27]), .ZN(n87) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[58]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[26]), .ZN(n86) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n85) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[56]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[24]), .ZN(n84) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[55]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[23]), .ZN(n83) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[54]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[22]), .ZN(n82) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[53]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[21]), .ZN(n81) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[52]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[51]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n47) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n47), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD2BWP30P140 U100 ( .I(n36), .ZN(n46) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[35]), .ZN(n37) );
  OAI22D1BWP30P140 U102 ( .A1(n47), .A2(n61), .B1(n46), .B2(n37), .ZN(N290) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[39]), .ZN(n38) );
  OAI22D1BWP30P140 U105 ( .A1(n42), .A2(n64), .B1(n46), .B2(n38), .ZN(N294) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U108 ( .A1(n42), .A2(n62), .B1(n46), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[5]), .ZN(n65) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[37]), .ZN(n40) );
  OAI22D1BWP30P140 U111 ( .A1(n42), .A2(n65), .B1(n46), .B2(n40), .ZN(N292) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[38]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n42), .A2(n63), .B1(n46), .B2(n41), .ZN(N293) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U117 ( .A1(n47), .A2(n59), .B1(n46), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[34]), .ZN(n44) );
  OAI22D1BWP30P140 U120 ( .A1(n47), .A2(n60), .B1(n46), .B2(n44), .ZN(N289) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n58) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n45) );
  OAI22D1BWP30P140 U123 ( .A1(n47), .A2(n58), .B1(n46), .B2(n45), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U125 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U127 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  MUX2NUD1BWP30P140 U128 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  INVD2BWP30P140 U137 ( .I(n79), .ZN(n77) );
  MOAI22D1BWP30P140 U138 ( .A1(n66), .A2(n77), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U139 ( .A1(n67), .A2(n77), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U140 ( .A1(n68), .A2(n77), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U141 ( .A1(n69), .A2(n77), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U142 ( .A1(n70), .A2(n77), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U143 ( .A1(n71), .A2(n77), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U144 ( .A1(n72), .A2(n77), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U145 ( .A1(n73), .A2(n77), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U146 ( .A1(n74), .A2(n77), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U147 ( .A1(n75), .A2(n77), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U148 ( .A1(n76), .A2(n77), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n77), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n92), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_106 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n33), .A2(n32), .B1(n31), .B2(n78), .ZN(N306) );
  INVD2BWP30P140 U4 ( .I(n36), .ZN(n46) );
  OAI22D1BWP30P140 U5 ( .A1(n42), .A2(n61), .B1(n46), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U6 ( .I(n57), .ZN(n79) );
  ND2D1BWP30P140 U7 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U9 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U10 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U11 ( .A1(n33), .A2(n17), .B1(n47), .B2(n66), .ZN(N295) );
  OAI22D1BWP30P140 U12 ( .A1(n33), .A2(n16), .B1(n47), .B2(n67), .ZN(N296) );
  OAI22D1BWP30P140 U13 ( .A1(n33), .A2(n15), .B1(n47), .B2(n68), .ZN(N297) );
  OAI22D1BWP30P140 U14 ( .A1(n33), .A2(n14), .B1(n47), .B2(n69), .ZN(N298) );
  OAI22D1BWP30P140 U15 ( .A1(n33), .A2(n13), .B1(n47), .B2(n70), .ZN(N299) );
  OAI22D1BWP30P140 U16 ( .A1(n33), .A2(n12), .B1(n47), .B2(n71), .ZN(N300) );
  OAI22D1BWP30P140 U17 ( .A1(n33), .A2(n11), .B1(n47), .B2(n72), .ZN(N301) );
  OAI22D1BWP30P140 U18 ( .A1(n33), .A2(n10), .B1(n47), .B2(n73), .ZN(N302) );
  OAI22D1BWP30P140 U19 ( .A1(n33), .A2(n9), .B1(n47), .B2(n74), .ZN(N303) );
  OAI22D1BWP30P140 U20 ( .A1(n33), .A2(n8), .B1(n47), .B2(n75), .ZN(N304) );
  OAI22D1BWP30P140 U21 ( .A1(n33), .A2(n7), .B1(n47), .B2(n76), .ZN(N305) );
  OAI22D1BWP30P140 U22 ( .A1(n30), .A2(n29), .B1(n31), .B2(n80), .ZN(N307) );
  OAI22D1BWP30P140 U23 ( .A1(n30), .A2(n28), .B1(n31), .B2(n81), .ZN(N308) );
  OAI22D1BWP30P140 U24 ( .A1(n30), .A2(n27), .B1(n31), .B2(n82), .ZN(N309) );
  OAI22D1BWP30P140 U25 ( .A1(n30), .A2(n26), .B1(n31), .B2(n83), .ZN(N310) );
  OAI22D1BWP30P140 U26 ( .A1(n30), .A2(n25), .B1(n31), .B2(n84), .ZN(N311) );
  OAI22D1BWP30P140 U27 ( .A1(n30), .A2(n24), .B1(n31), .B2(n85), .ZN(N312) );
  OAI22D1BWP30P140 U28 ( .A1(n30), .A2(n23), .B1(n31), .B2(n86), .ZN(N313) );
  OAI22D1BWP30P140 U29 ( .A1(n30), .A2(n22), .B1(n31), .B2(n87), .ZN(N314) );
  OAI22D1BWP30P140 U30 ( .A1(n30), .A2(n21), .B1(n31), .B2(n88), .ZN(N315) );
  OAI22D1BWP30P140 U31 ( .A1(n30), .A2(n20), .B1(n31), .B2(n89), .ZN(N316) );
  OAI22D1BWP30P140 U32 ( .A1(n30), .A2(n19), .B1(n31), .B2(n90), .ZN(N317) );
  OAI22D1BWP30P140 U33 ( .A1(n30), .A2(n18), .B1(n31), .B2(n93), .ZN(N318) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[50]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n47) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[18]), .ZN(n76) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[49]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[17]), .ZN(n75) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[48]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[16]), .ZN(n74) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[47]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[15]), .ZN(n73) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[46]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[14]), .ZN(n72) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n71) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[44]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[12]), .ZN(n70) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[43]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[42]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[10]), .ZN(n68) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[41]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[9]), .ZN(n67) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[40]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD2BWP30P140 U69 ( .I(n36), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[63]), .ZN(n18) );
  INVD2BWP30P140 U71 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[31]), .ZN(n93) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[62]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[30]), .ZN(n90) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[61]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[29]), .ZN(n89) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[60]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[28]), .ZN(n88) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[59]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[27]), .ZN(n87) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[58]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[26]), .ZN(n86) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n85) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[56]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[24]), .ZN(n84) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[55]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[23]), .ZN(n83) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[54]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[22]), .ZN(n82) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[53]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[21]), .ZN(n81) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[52]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[51]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n42) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n42), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n65) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[39]), .ZN(n37) );
  OAI22D1BWP30P140 U101 ( .A1(n47), .A2(n65), .B1(n46), .B2(n37), .ZN(N294) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[0]), .ZN(n58) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[32]), .ZN(n38) );
  OAI22D1BWP30P140 U104 ( .A1(n42), .A2(n58), .B1(n46), .B2(n38), .ZN(N287) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[33]), .ZN(n39) );
  OAI22D1BWP30P140 U107 ( .A1(n42), .A2(n59), .B1(n46), .B2(n39), .ZN(N288) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[34]), .ZN(n40) );
  OAI22D1BWP30P140 U110 ( .A1(n42), .A2(n60), .B1(n46), .B2(n40), .ZN(N289) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[35]), .ZN(n41) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[36]), .ZN(n43) );
  OAI22D1BWP30P140 U115 ( .A1(n47), .A2(n62), .B1(n46), .B2(n43), .ZN(N291) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[5]), .ZN(n63) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[37]), .ZN(n44) );
  OAI22D1BWP30P140 U118 ( .A1(n47), .A2(n63), .B1(n46), .B2(n44), .ZN(N292) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[6]), .ZN(n64) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[38]), .ZN(n45) );
  OAI22D1BWP30P140 U121 ( .A1(n47), .A2(n64), .B1(n46), .B2(n45), .ZN(N293) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  INVD2BWP30P140 U136 ( .I(n79), .ZN(n77) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n77), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n77), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n77), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n77), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n77), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n77), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n77), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n77), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n77), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n77), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n77), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n77), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  INVD2BWP30P140 U149 ( .I(n79), .ZN(n92) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n92), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_107 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD1BWP30P140 U3 ( .I(n57), .ZN(n79) );
  INVD2BWP30P140 U4 ( .I(n79), .ZN(n92) );
  NR2D1BWP30P140 U5 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  OAI22D1BWP30P140 U6 ( .A1(n33), .A2(n17), .B1(n44), .B2(n66), .ZN(N295) );
  OAI22D1BWP30P140 U7 ( .A1(n33), .A2(n16), .B1(n44), .B2(n67), .ZN(N296) );
  OAI22D1BWP30P140 U8 ( .A1(n33), .A2(n15), .B1(n44), .B2(n68), .ZN(N297) );
  OAI22D1BWP30P140 U9 ( .A1(n33), .A2(n14), .B1(n44), .B2(n69), .ZN(N298) );
  OAI22D1BWP30P140 U10 ( .A1(n33), .A2(n13), .B1(n44), .B2(n70), .ZN(N299) );
  OAI22D1BWP30P140 U11 ( .A1(n33), .A2(n12), .B1(n44), .B2(n71), .ZN(N300) );
  OAI22D1BWP30P140 U12 ( .A1(n33), .A2(n11), .B1(n44), .B2(n72), .ZN(N301) );
  OAI22D1BWP30P140 U13 ( .A1(n33), .A2(n10), .B1(n44), .B2(n73), .ZN(N302) );
  OAI22D1BWP30P140 U14 ( .A1(n33), .A2(n9), .B1(n44), .B2(n74), .ZN(N303) );
  OAI22D1BWP30P140 U15 ( .A1(n33), .A2(n8), .B1(n44), .B2(n75), .ZN(N304) );
  OAI22D1BWP30P140 U16 ( .A1(n33), .A2(n7), .B1(n44), .B2(n76), .ZN(N305) );
  OAI22D1BWP30P140 U17 ( .A1(n30), .A2(n29), .B1(n31), .B2(n80), .ZN(N307) );
  OAI22D1BWP30P140 U18 ( .A1(n30), .A2(n28), .B1(n31), .B2(n81), .ZN(N308) );
  OAI22D1BWP30P140 U19 ( .A1(n30), .A2(n27), .B1(n31), .B2(n82), .ZN(N309) );
  OAI22D1BWP30P140 U20 ( .A1(n30), .A2(n26), .B1(n31), .B2(n83), .ZN(N310) );
  OAI22D1BWP30P140 U21 ( .A1(n30), .A2(n25), .B1(n31), .B2(n84), .ZN(N311) );
  OAI22D1BWP30P140 U22 ( .A1(n30), .A2(n24), .B1(n31), .B2(n85), .ZN(N312) );
  OAI22D1BWP30P140 U23 ( .A1(n30), .A2(n23), .B1(n31), .B2(n86), .ZN(N313) );
  OAI22D1BWP30P140 U24 ( .A1(n30), .A2(n22), .B1(n31), .B2(n87), .ZN(N314) );
  OAI22D1BWP30P140 U25 ( .A1(n30), .A2(n21), .B1(n31), .B2(n88), .ZN(N315) );
  OAI22D1BWP30P140 U26 ( .A1(n30), .A2(n20), .B1(n31), .B2(n89), .ZN(N316) );
  OAI22D1BWP30P140 U27 ( .A1(n30), .A2(n19), .B1(n31), .B2(n90), .ZN(N317) );
  OAI22D1BWP30P140 U28 ( .A1(n30), .A2(n18), .B1(n31), .B2(n93), .ZN(N318) );
  ND2D1BWP30P140 U29 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U30 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U31 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U32 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U33 ( .A1(n33), .A2(n32), .B1(n31), .B2(n78), .ZN(N306) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[50]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n44) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[18]), .ZN(n76) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[49]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[17]), .ZN(n75) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[48]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[16]), .ZN(n74) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[47]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[15]), .ZN(n73) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[46]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[14]), .ZN(n72) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n71) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[44]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[12]), .ZN(n70) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[43]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[42]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[10]), .ZN(n68) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[41]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[9]), .ZN(n67) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[40]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD2BWP30P140 U69 ( .I(n36), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[63]), .ZN(n18) );
  INVD2BWP30P140 U71 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[31]), .ZN(n93) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[62]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[30]), .ZN(n90) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[61]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[29]), .ZN(n89) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[60]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[28]), .ZN(n88) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[59]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[27]), .ZN(n87) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[58]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[26]), .ZN(n86) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n85) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[56]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[24]), .ZN(n84) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[55]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[23]), .ZN(n83) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[54]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[22]), .ZN(n82) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[53]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[21]), .ZN(n81) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[52]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[51]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n47) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n47), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD2BWP30P140 U100 ( .I(n36), .ZN(n46) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[33]), .ZN(n37) );
  OAI22D1BWP30P140 U102 ( .A1(n47), .A2(n59), .B1(n46), .B2(n37), .ZN(N288) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[34]), .ZN(n38) );
  OAI22D1BWP30P140 U105 ( .A1(n47), .A2(n60), .B1(n46), .B2(n38), .ZN(N289) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[0]), .ZN(n58) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[32]), .ZN(n39) );
  OAI22D1BWP30P140 U108 ( .A1(n47), .A2(n58), .B1(n46), .B2(n39), .ZN(N287) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n40) );
  OAI22D1BWP30P140 U111 ( .A1(n44), .A2(n62), .B1(n46), .B2(n40), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[5]), .ZN(n63) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[37]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n44), .A2(n63), .B1(n46), .B2(n41), .ZN(N292) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[6]), .ZN(n64) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[38]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n44), .A2(n64), .B1(n46), .B2(n42), .ZN(N293) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[7]), .ZN(n65) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[39]), .ZN(n43) );
  OAI22D1BWP30P140 U120 ( .A1(n44), .A2(n65), .B1(n46), .B2(n43), .ZN(N294) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[35]), .ZN(n45) );
  OAI22D1BWP30P140 U123 ( .A1(n47), .A2(n61), .B1(n46), .B2(n45), .ZN(N290) );
  INVD1BWP30P140 U124 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U125 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U127 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  MUX2NUD1BWP30P140 U128 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  INVD2BWP30P140 U137 ( .I(n79), .ZN(n77) );
  MOAI22D1BWP30P140 U138 ( .A1(n66), .A2(n77), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U139 ( .A1(n67), .A2(n77), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U140 ( .A1(n68), .A2(n77), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U141 ( .A1(n69), .A2(n77), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U142 ( .A1(n70), .A2(n77), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U143 ( .A1(n71), .A2(n77), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U144 ( .A1(n72), .A2(n77), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U145 ( .A1(n73), .A2(n77), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U146 ( .A1(n74), .A2(n77), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U147 ( .A1(n75), .A2(n77), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U148 ( .A1(n76), .A2(n77), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n77), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n92), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_108 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n21), .A2(n20), .B1(n31), .B2(n78), .ZN(N306) );
  INVD2BWP30P140 U4 ( .I(n36), .ZN(n46) );
  OAI22D1BWP30P140 U5 ( .A1(n44), .A2(n60), .B1(n46), .B2(n43), .ZN(N289) );
  INVD1BWP30P140 U6 ( .I(n57), .ZN(n79) );
  ND2D1BWP30P140 U7 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U9 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U10 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U11 ( .A1(n21), .A2(n7), .B1(n47), .B2(n66), .ZN(N295) );
  OAI22D1BWP30P140 U12 ( .A1(n21), .A2(n8), .B1(n47), .B2(n67), .ZN(N296) );
  OAI22D1BWP30P140 U13 ( .A1(n21), .A2(n9), .B1(n47), .B2(n68), .ZN(N297) );
  OAI22D1BWP30P140 U14 ( .A1(n21), .A2(n10), .B1(n47), .B2(n69), .ZN(N298) );
  OAI22D1BWP30P140 U15 ( .A1(n21), .A2(n11), .B1(n47), .B2(n70), .ZN(N299) );
  OAI22D1BWP30P140 U16 ( .A1(n21), .A2(n12), .B1(n47), .B2(n71), .ZN(N300) );
  OAI22D1BWP30P140 U17 ( .A1(n21), .A2(n13), .B1(n47), .B2(n72), .ZN(N301) );
  OAI22D1BWP30P140 U18 ( .A1(n21), .A2(n14), .B1(n47), .B2(n73), .ZN(N302) );
  OAI22D1BWP30P140 U19 ( .A1(n21), .A2(n15), .B1(n47), .B2(n74), .ZN(N303) );
  OAI22D1BWP30P140 U20 ( .A1(n21), .A2(n16), .B1(n47), .B2(n75), .ZN(N304) );
  OAI22D1BWP30P140 U21 ( .A1(n21), .A2(n17), .B1(n47), .B2(n76), .ZN(N305) );
  OAI22D1BWP30P140 U22 ( .A1(n33), .A2(n22), .B1(n31), .B2(n80), .ZN(N307) );
  OAI22D1BWP30P140 U23 ( .A1(n33), .A2(n23), .B1(n31), .B2(n81), .ZN(N308) );
  OAI22D1BWP30P140 U24 ( .A1(n33), .A2(n24), .B1(n31), .B2(n82), .ZN(N309) );
  OAI22D1BWP30P140 U25 ( .A1(n33), .A2(n25), .B1(n31), .B2(n83), .ZN(N310) );
  OAI22D1BWP30P140 U26 ( .A1(n33), .A2(n26), .B1(n31), .B2(n84), .ZN(N311) );
  OAI22D1BWP30P140 U27 ( .A1(n33), .A2(n27), .B1(n31), .B2(n85), .ZN(N312) );
  OAI22D1BWP30P140 U28 ( .A1(n33), .A2(n28), .B1(n31), .B2(n86), .ZN(N313) );
  OAI22D1BWP30P140 U29 ( .A1(n33), .A2(n29), .B1(n31), .B2(n87), .ZN(N314) );
  OAI22D1BWP30P140 U30 ( .A1(n33), .A2(n30), .B1(n31), .B2(n88), .ZN(N315) );
  OAI22D1BWP30P140 U31 ( .A1(n33), .A2(n32), .B1(n31), .B2(n89), .ZN(N316) );
  OAI22D1BWP30P140 U32 ( .A1(n33), .A2(n19), .B1(n31), .B2(n90), .ZN(N317) );
  OAI22D1BWP30P140 U33 ( .A1(n33), .A2(n18), .B1(n31), .B2(n93), .ZN(N318) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n21) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n47) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n67) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n68) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n70) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n71) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[14]), .ZN(n72) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[47]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[15]), .ZN(n73) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[48]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n74) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n75) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n76) );
  INVD2BWP30P140 U69 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[63]), .ZN(n18) );
  INVD2BWP30P140 U71 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[31]), .ZN(n93) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[62]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[30]), .ZN(n90) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[51]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[52]), .ZN(n22) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[53]), .ZN(n23) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[21]), .ZN(n81) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[54]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[22]), .ZN(n82) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[55]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[23]), .ZN(n83) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[56]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[24]), .ZN(n84) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[57]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[25]), .ZN(n85) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[58]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[26]), .ZN(n86) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[59]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[27]), .ZN(n87) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[60]), .ZN(n30) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[28]), .ZN(n88) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[61]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[29]), .ZN(n89) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n44) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n44), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[35]), .ZN(n37) );
  OAI22D1BWP30P140 U101 ( .A1(n44), .A2(n61), .B1(n46), .B2(n37), .ZN(N290) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[36]), .ZN(n38) );
  OAI22D1BWP30P140 U104 ( .A1(n47), .A2(n62), .B1(n46), .B2(n38), .ZN(N291) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[5]), .ZN(n63) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[37]), .ZN(n39) );
  OAI22D1BWP30P140 U107 ( .A1(n47), .A2(n63), .B1(n46), .B2(n39), .ZN(N292) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[6]), .ZN(n64) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[38]), .ZN(n40) );
  OAI22D1BWP30P140 U110 ( .A1(n47), .A2(n64), .B1(n46), .B2(n40), .ZN(N293) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[0]), .ZN(n58) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[32]), .ZN(n41) );
  OAI22D1BWP30P140 U113 ( .A1(n44), .A2(n58), .B1(n46), .B2(n41), .ZN(N287) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[33]), .ZN(n42) );
  OAI22D1BWP30P140 U116 ( .A1(n44), .A2(n59), .B1(n46), .B2(n42), .ZN(N288) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[34]), .ZN(n43) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[7]), .ZN(n65) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[39]), .ZN(n45) );
  OAI22D1BWP30P140 U121 ( .A1(n47), .A2(n65), .B1(n46), .B2(n45), .ZN(N294) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  INVD2BWP30P140 U136 ( .I(n79), .ZN(n77) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n77), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n77), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n77), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n77), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n77), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n77), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n77), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n77), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n77), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n77), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n77), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n77), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  INVD2BWP30P140 U149 ( .I(n79), .ZN(n92) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n92), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_109 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD1BWP30P140 U3 ( .I(n57), .ZN(n79) );
  OAI22D1BWP30P140 U4 ( .A1(n19), .A2(n18), .B1(n31), .B2(n78), .ZN(N306) );
  INVD2BWP30P140 U5 ( .I(n79), .ZN(n92) );
  NR2D1BWP30P140 U6 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  OAI22D1BWP30P140 U7 ( .A1(n19), .A2(n7), .B1(n47), .B2(n66), .ZN(N295) );
  OAI22D1BWP30P140 U8 ( .A1(n19), .A2(n8), .B1(n47), .B2(n67), .ZN(N296) );
  OAI22D1BWP30P140 U9 ( .A1(n19), .A2(n9), .B1(n47), .B2(n68), .ZN(N297) );
  OAI22D1BWP30P140 U10 ( .A1(n19), .A2(n10), .B1(n47), .B2(n69), .ZN(N298) );
  OAI22D1BWP30P140 U11 ( .A1(n19), .A2(n11), .B1(n47), .B2(n70), .ZN(N299) );
  OAI22D1BWP30P140 U12 ( .A1(n19), .A2(n12), .B1(n47), .B2(n71), .ZN(N300) );
  OAI22D1BWP30P140 U13 ( .A1(n19), .A2(n13), .B1(n47), .B2(n72), .ZN(N301) );
  OAI22D1BWP30P140 U14 ( .A1(n19), .A2(n14), .B1(n47), .B2(n73), .ZN(N302) );
  OAI22D1BWP30P140 U15 ( .A1(n19), .A2(n15), .B1(n47), .B2(n74), .ZN(N303) );
  OAI22D1BWP30P140 U16 ( .A1(n19), .A2(n16), .B1(n47), .B2(n75), .ZN(N304) );
  OAI22D1BWP30P140 U17 ( .A1(n19), .A2(n17), .B1(n47), .B2(n76), .ZN(N305) );
  ND2D1BWP30P140 U18 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U19 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U20 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U21 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U22 ( .A1(n33), .A2(n20), .B1(n31), .B2(n80), .ZN(N307) );
  OAI22D1BWP30P140 U23 ( .A1(n33), .A2(n21), .B1(n31), .B2(n81), .ZN(N308) );
  OAI22D1BWP30P140 U24 ( .A1(n33), .A2(n22), .B1(n31), .B2(n82), .ZN(N309) );
  OAI22D1BWP30P140 U25 ( .A1(n33), .A2(n23), .B1(n31), .B2(n83), .ZN(N310) );
  OAI22D1BWP30P140 U26 ( .A1(n33), .A2(n24), .B1(n31), .B2(n84), .ZN(N311) );
  OAI22D1BWP30P140 U27 ( .A1(n33), .A2(n25), .B1(n31), .B2(n85), .ZN(N312) );
  OAI22D1BWP30P140 U28 ( .A1(n33), .A2(n26), .B1(n31), .B2(n86), .ZN(N313) );
  OAI22D1BWP30P140 U29 ( .A1(n33), .A2(n27), .B1(n31), .B2(n87), .ZN(N314) );
  OAI22D1BWP30P140 U30 ( .A1(n33), .A2(n28), .B1(n31), .B2(n88), .ZN(N315) );
  OAI22D1BWP30P140 U31 ( .A1(n33), .A2(n29), .B1(n31), .B2(n89), .ZN(N316) );
  OAI22D1BWP30P140 U32 ( .A1(n33), .A2(n30), .B1(n31), .B2(n90), .ZN(N317) );
  OAI22D1BWP30P140 U33 ( .A1(n33), .A2(n32), .B1(n31), .B2(n93), .ZN(N318) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n19) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n47) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n67) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n68) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n70) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n71) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[14]), .ZN(n72) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[47]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[15]), .ZN(n73) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[48]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n74) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n75) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n76) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n18) );
  INVD2BWP30P140 U70 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD2BWP30P140 U72 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n20) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n21) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n81) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n22) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n82) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n23) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n83) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n84) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n85) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n86) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n87) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n88) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n89) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n30) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n90) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n93) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n41) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n41), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[0]), .ZN(n58) );
  INVD2BWP30P140 U100 ( .I(n36), .ZN(n46) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[32]), .ZN(n37) );
  OAI22D1BWP30P140 U102 ( .A1(n41), .A2(n58), .B1(n46), .B2(n37), .ZN(N287) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[33]), .ZN(n38) );
  OAI22D1BWP30P140 U105 ( .A1(n41), .A2(n59), .B1(n46), .B2(n38), .ZN(N288) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[34]), .ZN(n39) );
  OAI22D1BWP30P140 U108 ( .A1(n41), .A2(n60), .B1(n46), .B2(n39), .ZN(N289) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[35]), .ZN(n40) );
  OAI22D1BWP30P140 U111 ( .A1(n41), .A2(n61), .B1(n46), .B2(n40), .ZN(N290) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[36]), .ZN(n42) );
  OAI22D1BWP30P140 U114 ( .A1(n47), .A2(n62), .B1(n46), .B2(n42), .ZN(N291) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[5]), .ZN(n63) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[37]), .ZN(n43) );
  OAI22D1BWP30P140 U117 ( .A1(n47), .A2(n63), .B1(n46), .B2(n43), .ZN(N292) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[6]), .ZN(n64) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[38]), .ZN(n44) );
  OAI22D1BWP30P140 U120 ( .A1(n47), .A2(n64), .B1(n46), .B2(n44), .ZN(N293) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[7]), .ZN(n65) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[39]), .ZN(n45) );
  OAI22D1BWP30P140 U123 ( .A1(n47), .A2(n65), .B1(n46), .B2(n45), .ZN(N294) );
  INVD1BWP30P140 U124 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U125 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U127 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  MUX2NUD1BWP30P140 U128 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  INVD2BWP30P140 U137 ( .I(n79), .ZN(n77) );
  MOAI22D1BWP30P140 U138 ( .A1(n66), .A2(n77), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U139 ( .A1(n67), .A2(n77), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U140 ( .A1(n68), .A2(n77), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U141 ( .A1(n69), .A2(n77), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U142 ( .A1(n70), .A2(n77), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U143 ( .A1(n71), .A2(n77), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U144 ( .A1(n72), .A2(n77), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U145 ( .A1(n73), .A2(n77), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U146 ( .A1(n74), .A2(n77), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U147 ( .A1(n75), .A2(n77), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U148 ( .A1(n76), .A2(n77), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n77), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n92), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_110 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n19), .A2(n18), .B1(n31), .B2(n78), .ZN(N306) );
  INVD2BWP30P140 U4 ( .I(n36), .ZN(n46) );
  OAI22D1BWP30P140 U5 ( .A1(n41), .A2(n61), .B1(n46), .B2(n40), .ZN(N290) );
  INVD1BWP30P140 U6 ( .I(n57), .ZN(n79) );
  ND2D1BWP30P140 U7 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U9 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U10 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U11 ( .A1(n19), .A2(n13), .B1(n47), .B2(n66), .ZN(N295) );
  OAI22D1BWP30P140 U12 ( .A1(n19), .A2(n14), .B1(n47), .B2(n67), .ZN(N296) );
  OAI22D1BWP30P140 U13 ( .A1(n19), .A2(n15), .B1(n47), .B2(n68), .ZN(N297) );
  OAI22D1BWP30P140 U14 ( .A1(n19), .A2(n16), .B1(n47), .B2(n69), .ZN(N298) );
  OAI22D1BWP30P140 U15 ( .A1(n19), .A2(n17), .B1(n47), .B2(n70), .ZN(N299) );
  OAI22D1BWP30P140 U16 ( .A1(n19), .A2(n12), .B1(n47), .B2(n71), .ZN(N300) );
  OAI22D1BWP30P140 U17 ( .A1(n19), .A2(n11), .B1(n47), .B2(n72), .ZN(N301) );
  OAI22D1BWP30P140 U18 ( .A1(n19), .A2(n7), .B1(n47), .B2(n73), .ZN(N302) );
  OAI22D1BWP30P140 U19 ( .A1(n19), .A2(n8), .B1(n47), .B2(n74), .ZN(N303) );
  OAI22D1BWP30P140 U20 ( .A1(n19), .A2(n9), .B1(n47), .B2(n75), .ZN(N304) );
  OAI22D1BWP30P140 U21 ( .A1(n19), .A2(n10), .B1(n47), .B2(n76), .ZN(N305) );
  OAI22D1BWP30P140 U22 ( .A1(n33), .A2(n20), .B1(n31), .B2(n80), .ZN(N307) );
  OAI22D1BWP30P140 U23 ( .A1(n33), .A2(n21), .B1(n31), .B2(n81), .ZN(N308) );
  OAI22D1BWP30P140 U24 ( .A1(n33), .A2(n22), .B1(n31), .B2(n82), .ZN(N309) );
  OAI22D1BWP30P140 U25 ( .A1(n33), .A2(n23), .B1(n31), .B2(n83), .ZN(N310) );
  OAI22D1BWP30P140 U26 ( .A1(n33), .A2(n24), .B1(n31), .B2(n84), .ZN(N311) );
  OAI22D1BWP30P140 U27 ( .A1(n33), .A2(n25), .B1(n31), .B2(n85), .ZN(N312) );
  OAI22D1BWP30P140 U28 ( .A1(n33), .A2(n26), .B1(n31), .B2(n86), .ZN(N313) );
  OAI22D1BWP30P140 U29 ( .A1(n33), .A2(n27), .B1(n31), .B2(n87), .ZN(N314) );
  OAI22D1BWP30P140 U30 ( .A1(n33), .A2(n28), .B1(n31), .B2(n88), .ZN(N315) );
  OAI22D1BWP30P140 U31 ( .A1(n33), .A2(n29), .B1(n31), .B2(n89), .ZN(N316) );
  OAI22D1BWP30P140 U32 ( .A1(n33), .A2(n30), .B1(n31), .B2(n90), .ZN(N317) );
  OAI22D1BWP30P140 U33 ( .A1(n33), .A2(n32), .B1(n31), .B2(n93), .ZN(N318) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n19) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[47]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n47) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[15]), .ZN(n73) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[48]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[16]), .ZN(n74) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[49]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[17]), .ZN(n75) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[50]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[18]), .ZN(n76) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[46]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[14]), .ZN(n72) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n71) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[40]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[41]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[9]), .ZN(n67) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[42]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[10]), .ZN(n68) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[43]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[44]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[12]), .ZN(n70) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n18) );
  INVD2BWP30P140 U70 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD2BWP30P140 U72 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n20) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n21) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n81) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n22) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n82) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n23) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n83) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n84) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n85) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n86) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n87) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n88) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n89) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n30) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n90) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n93) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n41) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n41), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[0]), .ZN(n58) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[32]), .ZN(n37) );
  OAI22D1BWP30P140 U101 ( .A1(n41), .A2(n58), .B1(n46), .B2(n37), .ZN(N287) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[33]), .ZN(n38) );
  OAI22D1BWP30P140 U104 ( .A1(n41), .A2(n59), .B1(n46), .B2(n38), .ZN(N288) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[34]), .ZN(n39) );
  OAI22D1BWP30P140 U107 ( .A1(n41), .A2(n60), .B1(n46), .B2(n39), .ZN(N289) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[35]), .ZN(n40) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[36]), .ZN(n42) );
  OAI22D1BWP30P140 U112 ( .A1(n47), .A2(n62), .B1(n46), .B2(n42), .ZN(N291) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[5]), .ZN(n63) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[37]), .ZN(n43) );
  OAI22D1BWP30P140 U115 ( .A1(n47), .A2(n63), .B1(n46), .B2(n43), .ZN(N292) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[6]), .ZN(n64) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[38]), .ZN(n44) );
  OAI22D1BWP30P140 U118 ( .A1(n47), .A2(n64), .B1(n46), .B2(n44), .ZN(N293) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[7]), .ZN(n65) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[39]), .ZN(n45) );
  OAI22D1BWP30P140 U121 ( .A1(n47), .A2(n65), .B1(n46), .B2(n45), .ZN(N294) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  INVD2BWP30P140 U136 ( .I(n79), .ZN(n77) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n77), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n77), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n77), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n77), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n77), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n77), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n77), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n77), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n77), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n77), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n77), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n77), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  INVD2BWP30P140 U149 ( .I(n79), .ZN(n92) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n92), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_111 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD1BWP30P140 U3 ( .I(n57), .ZN(n79) );
  INVD2BWP30P140 U4 ( .I(n79), .ZN(n92) );
  NR2D1BWP30P140 U5 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  OAI22D1BWP30P140 U6 ( .A1(n19), .A2(n7), .B1(n41), .B2(n66), .ZN(N295) );
  OAI22D1BWP30P140 U7 ( .A1(n19), .A2(n8), .B1(n41), .B2(n67), .ZN(N296) );
  OAI22D1BWP30P140 U8 ( .A1(n19), .A2(n9), .B1(n41), .B2(n68), .ZN(N297) );
  OAI22D1BWP30P140 U9 ( .A1(n19), .A2(n10), .B1(n41), .B2(n69), .ZN(N298) );
  OAI22D1BWP30P140 U10 ( .A1(n19), .A2(n11), .B1(n41), .B2(n70), .ZN(N299) );
  OAI22D1BWP30P140 U11 ( .A1(n19), .A2(n12), .B1(n41), .B2(n71), .ZN(N300) );
  OAI22D1BWP30P140 U12 ( .A1(n19), .A2(n13), .B1(n41), .B2(n72), .ZN(N301) );
  OAI22D1BWP30P140 U13 ( .A1(n19), .A2(n14), .B1(n41), .B2(n73), .ZN(N302) );
  OAI22D1BWP30P140 U14 ( .A1(n19), .A2(n15), .B1(n41), .B2(n74), .ZN(N303) );
  OAI22D1BWP30P140 U15 ( .A1(n19), .A2(n16), .B1(n41), .B2(n75), .ZN(N304) );
  OAI22D1BWP30P140 U16 ( .A1(n19), .A2(n17), .B1(n41), .B2(n76), .ZN(N305) );
  OAI22D1BWP30P140 U17 ( .A1(n33), .A2(n20), .B1(n31), .B2(n80), .ZN(N307) );
  OAI22D1BWP30P140 U18 ( .A1(n33), .A2(n21), .B1(n31), .B2(n81), .ZN(N308) );
  OAI22D1BWP30P140 U19 ( .A1(n33), .A2(n22), .B1(n31), .B2(n82), .ZN(N309) );
  OAI22D1BWP30P140 U20 ( .A1(n33), .A2(n23), .B1(n31), .B2(n83), .ZN(N310) );
  OAI22D1BWP30P140 U21 ( .A1(n33), .A2(n24), .B1(n31), .B2(n84), .ZN(N311) );
  OAI22D1BWP30P140 U22 ( .A1(n33), .A2(n25), .B1(n31), .B2(n85), .ZN(N312) );
  OAI22D1BWP30P140 U23 ( .A1(n33), .A2(n26), .B1(n31), .B2(n86), .ZN(N313) );
  OAI22D1BWP30P140 U24 ( .A1(n33), .A2(n27), .B1(n31), .B2(n87), .ZN(N314) );
  OAI22D1BWP30P140 U25 ( .A1(n33), .A2(n28), .B1(n31), .B2(n88), .ZN(N315) );
  OAI22D1BWP30P140 U26 ( .A1(n33), .A2(n29), .B1(n31), .B2(n89), .ZN(N316) );
  OAI22D1BWP30P140 U27 ( .A1(n33), .A2(n30), .B1(n31), .B2(n90), .ZN(N317) );
  OAI22D1BWP30P140 U28 ( .A1(n33), .A2(n32), .B1(n31), .B2(n93), .ZN(N318) );
  ND2D1BWP30P140 U29 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U30 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U31 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U32 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U33 ( .A1(n19), .A2(n18), .B1(n31), .B2(n78), .ZN(N306) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n19) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n41) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n67) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n68) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n70) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n71) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[14]), .ZN(n72) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[47]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[15]), .ZN(n73) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[48]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n74) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n75) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n76) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n18) );
  INVD2BWP30P140 U70 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD2BWP30P140 U72 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n20) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n21) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n81) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n22) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n82) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n23) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n83) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n84) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n85) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n86) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n87) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n88) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n89) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n30) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n90) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n93) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n47) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n47), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n65) );
  INVD2BWP30P140 U100 ( .I(n36), .ZN(n46) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n37) );
  OAI22D1BWP30P140 U102 ( .A1(n41), .A2(n65), .B1(n46), .B2(n37), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n64) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n38) );
  OAI22D1BWP30P140 U105 ( .A1(n41), .A2(n64), .B1(n46), .B2(n38), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n63) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n39) );
  OAI22D1BWP30P140 U108 ( .A1(n41), .A2(n63), .B1(n46), .B2(n39), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n40) );
  OAI22D1BWP30P140 U111 ( .A1(n41), .A2(n62), .B1(n46), .B2(n40), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U114 ( .A1(n47), .A2(n60), .B1(n46), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U117 ( .A1(n47), .A2(n59), .B1(n46), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[0]), .ZN(n58) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U120 ( .A1(n47), .A2(n58), .B1(n46), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[35]), .ZN(n45) );
  OAI22D1BWP30P140 U123 ( .A1(n47), .A2(n61), .B1(n46), .B2(n45), .ZN(N290) );
  INVD1BWP30P140 U124 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U125 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U127 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  MUX2NUD1BWP30P140 U128 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  INVD2BWP30P140 U137 ( .I(n79), .ZN(n77) );
  MOAI22D1BWP30P140 U138 ( .A1(n66), .A2(n77), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U139 ( .A1(n67), .A2(n77), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U140 ( .A1(n68), .A2(n77), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U141 ( .A1(n69), .A2(n77), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U142 ( .A1(n70), .A2(n77), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U143 ( .A1(n71), .A2(n77), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U144 ( .A1(n72), .A2(n77), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U145 ( .A1(n73), .A2(n77), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U146 ( .A1(n74), .A2(n77), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U147 ( .A1(n75), .A2(n77), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U148 ( .A1(n76), .A2(n77), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n77), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n92), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_112 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n19), .A2(n18), .B1(n31), .B2(n78), .ZN(N306) );
  INVD2BWP30P140 U4 ( .I(n36), .ZN(n46) );
  OAI22D1BWP30P140 U5 ( .A1(n41), .A2(n60), .B1(n46), .B2(n40), .ZN(N290) );
  INVD1BWP30P140 U6 ( .I(n57), .ZN(n79) );
  ND2D1BWP30P140 U7 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U9 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U10 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U11 ( .A1(n19), .A2(n7), .B1(n47), .B2(n66), .ZN(N295) );
  OAI22D1BWP30P140 U12 ( .A1(n19), .A2(n8), .B1(n47), .B2(n67), .ZN(N296) );
  OAI22D1BWP30P140 U13 ( .A1(n19), .A2(n9), .B1(n47), .B2(n68), .ZN(N297) );
  OAI22D1BWP30P140 U14 ( .A1(n19), .A2(n10), .B1(n47), .B2(n69), .ZN(N298) );
  OAI22D1BWP30P140 U15 ( .A1(n19), .A2(n11), .B1(n47), .B2(n70), .ZN(N299) );
  OAI22D1BWP30P140 U16 ( .A1(n19), .A2(n12), .B1(n47), .B2(n71), .ZN(N300) );
  OAI22D1BWP30P140 U17 ( .A1(n19), .A2(n13), .B1(n47), .B2(n72), .ZN(N301) );
  OAI22D1BWP30P140 U18 ( .A1(n19), .A2(n14), .B1(n47), .B2(n73), .ZN(N302) );
  OAI22D1BWP30P140 U19 ( .A1(n19), .A2(n15), .B1(n47), .B2(n74), .ZN(N303) );
  OAI22D1BWP30P140 U20 ( .A1(n19), .A2(n16), .B1(n47), .B2(n75), .ZN(N304) );
  OAI22D1BWP30P140 U21 ( .A1(n19), .A2(n17), .B1(n47), .B2(n76), .ZN(N305) );
  OAI22D1BWP30P140 U22 ( .A1(n33), .A2(n20), .B1(n31), .B2(n80), .ZN(N307) );
  OAI22D1BWP30P140 U23 ( .A1(n33), .A2(n21), .B1(n31), .B2(n81), .ZN(N308) );
  OAI22D1BWP30P140 U24 ( .A1(n33), .A2(n22), .B1(n31), .B2(n82), .ZN(N309) );
  OAI22D1BWP30P140 U25 ( .A1(n33), .A2(n23), .B1(n31), .B2(n83), .ZN(N310) );
  OAI22D1BWP30P140 U26 ( .A1(n33), .A2(n24), .B1(n31), .B2(n84), .ZN(N311) );
  OAI22D1BWP30P140 U27 ( .A1(n33), .A2(n25), .B1(n31), .B2(n85), .ZN(N312) );
  OAI22D1BWP30P140 U28 ( .A1(n33), .A2(n26), .B1(n31), .B2(n86), .ZN(N313) );
  OAI22D1BWP30P140 U29 ( .A1(n33), .A2(n27), .B1(n31), .B2(n87), .ZN(N314) );
  OAI22D1BWP30P140 U30 ( .A1(n33), .A2(n28), .B1(n31), .B2(n88), .ZN(N315) );
  OAI22D1BWP30P140 U31 ( .A1(n33), .A2(n29), .B1(n31), .B2(n89), .ZN(N316) );
  OAI22D1BWP30P140 U32 ( .A1(n33), .A2(n30), .B1(n31), .B2(n90), .ZN(N317) );
  OAI22D1BWP30P140 U33 ( .A1(n33), .A2(n32), .B1(n31), .B2(n93), .ZN(N318) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n19) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n47) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n67) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n68) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n70) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n71) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[14]), .ZN(n72) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[47]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[15]), .ZN(n73) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[48]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n74) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n75) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n76) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n18) );
  INVD2BWP30P140 U70 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD2BWP30P140 U72 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n20) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n21) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n81) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n22) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n82) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n23) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n83) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n84) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n85) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n86) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n87) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n88) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n89) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n30) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n90) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n93) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n41) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n41), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[0]), .ZN(n58) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[32]), .ZN(n37) );
  OAI22D1BWP30P140 U101 ( .A1(n41), .A2(n58), .B1(n46), .B2(n37), .ZN(N287) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[1]), .ZN(n65) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[33]), .ZN(n38) );
  OAI22D1BWP30P140 U104 ( .A1(n41), .A2(n65), .B1(n46), .B2(n38), .ZN(N288) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[2]), .ZN(n59) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[34]), .ZN(n39) );
  OAI22D1BWP30P140 U107 ( .A1(n41), .A2(n59), .B1(n46), .B2(n39), .ZN(N289) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[3]), .ZN(n60) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[35]), .ZN(n40) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[36]), .ZN(n42) );
  OAI22D1BWP30P140 U112 ( .A1(n47), .A2(n61), .B1(n46), .B2(n42), .ZN(N291) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[37]), .ZN(n43) );
  OAI22D1BWP30P140 U115 ( .A1(n47), .A2(n62), .B1(n46), .B2(n43), .ZN(N292) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[6]), .ZN(n63) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[38]), .ZN(n44) );
  OAI22D1BWP30P140 U118 ( .A1(n47), .A2(n63), .B1(n46), .B2(n44), .ZN(N293) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[7]), .ZN(n64) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[39]), .ZN(n45) );
  OAI22D1BWP30P140 U121 ( .A1(n47), .A2(n64), .B1(n46), .B2(n45), .ZN(N294) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  INVD2BWP30P140 U136 ( .I(n79), .ZN(n77) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n77), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n77), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n77), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n77), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n77), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n77), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n77), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n77), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n77), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n77), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n77), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n77), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  INVD2BWP30P140 U149 ( .I(n79), .ZN(n92) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n92), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_113 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD1BWP30P140 U3 ( .I(n57), .ZN(n84) );
  INVD2BWP30P140 U4 ( .I(n84), .ZN(n80) );
  NR2D1BWP30P140 U5 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  OAI22D1BWP30P140 U6 ( .A1(n19), .A2(n7), .B1(n43), .B2(n58), .ZN(N295) );
  OAI22D1BWP30P140 U7 ( .A1(n19), .A2(n8), .B1(n43), .B2(n59), .ZN(N296) );
  OAI22D1BWP30P140 U8 ( .A1(n19), .A2(n9), .B1(n43), .B2(n60), .ZN(N297) );
  OAI22D1BWP30P140 U9 ( .A1(n19), .A2(n10), .B1(n43), .B2(n61), .ZN(N298) );
  OAI22D1BWP30P140 U10 ( .A1(n19), .A2(n11), .B1(n43), .B2(n62), .ZN(N299) );
  OAI22D1BWP30P140 U11 ( .A1(n19), .A2(n12), .B1(n43), .B2(n63), .ZN(N300) );
  OAI22D1BWP30P140 U12 ( .A1(n19), .A2(n13), .B1(n43), .B2(n83), .ZN(N301) );
  OAI22D1BWP30P140 U13 ( .A1(n19), .A2(n14), .B1(n43), .B2(n64), .ZN(N302) );
  OAI22D1BWP30P140 U14 ( .A1(n19), .A2(n15), .B1(n43), .B2(n65), .ZN(N303) );
  OAI22D1BWP30P140 U15 ( .A1(n19), .A2(n16), .B1(n43), .B2(n66), .ZN(N304) );
  OAI22D1BWP30P140 U16 ( .A1(n19), .A2(n17), .B1(n43), .B2(n67), .ZN(N305) );
  OAI22D1BWP30P140 U17 ( .A1(n33), .A2(n20), .B1(n31), .B2(n69), .ZN(N307) );
  OAI22D1BWP30P140 U18 ( .A1(n33), .A2(n21), .B1(n31), .B2(n70), .ZN(N308) );
  OAI22D1BWP30P140 U19 ( .A1(n33), .A2(n32), .B1(n31), .B2(n71), .ZN(N309) );
  OAI22D1BWP30P140 U20 ( .A1(n33), .A2(n22), .B1(n31), .B2(n72), .ZN(N310) );
  OAI22D1BWP30P140 U21 ( .A1(n33), .A2(n23), .B1(n31), .B2(n73), .ZN(N311) );
  OAI22D1BWP30P140 U22 ( .A1(n33), .A2(n24), .B1(n31), .B2(n74), .ZN(N312) );
  OAI22D1BWP30P140 U23 ( .A1(n33), .A2(n25), .B1(n31), .B2(n75), .ZN(N313) );
  OAI22D1BWP30P140 U24 ( .A1(n33), .A2(n26), .B1(n31), .B2(n76), .ZN(N314) );
  OAI22D1BWP30P140 U25 ( .A1(n33), .A2(n27), .B1(n31), .B2(n77), .ZN(N315) );
  OAI22D1BWP30P140 U26 ( .A1(n33), .A2(n28), .B1(n31), .B2(n78), .ZN(N316) );
  OAI22D1BWP30P140 U27 ( .A1(n33), .A2(n29), .B1(n31), .B2(n79), .ZN(N317) );
  OAI22D1BWP30P140 U28 ( .A1(n33), .A2(n30), .B1(n31), .B2(n81), .ZN(N318) );
  ND2D1BWP30P140 U29 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U30 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U31 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U32 ( .I(n92), .ZN(n50) );
  OAI22D1BWP30P140 U33 ( .A1(n19), .A2(n18), .B1(n31), .B2(n68), .ZN(N306) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n19) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n43) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n58) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n59) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n60) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n61) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n62) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n63) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[14]), .ZN(n83) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[47]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[15]), .ZN(n64) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[48]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n65) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n66) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n67) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n18) );
  INVD2BWP30P140 U70 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n68) );
  INVD2BWP30P140 U72 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n20) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n69) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n21) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n70) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[23]), .ZN(n72) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[56]), .ZN(n23) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[24]), .ZN(n73) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[25]), .ZN(n74) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[58]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[26]), .ZN(n75) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[27]), .ZN(n76) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[60]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[28]), .ZN(n77) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[61]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[29]), .ZN(n78) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[30]), .ZN(n79) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[63]), .ZN(n30) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[31]), .ZN(n81) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[54]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[22]), .ZN(n71) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n47) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n47), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[2]), .ZN(n87) );
  INVD2BWP30P140 U100 ( .I(n36), .ZN(n46) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[34]), .ZN(n37) );
  OAI22D1BWP30P140 U102 ( .A1(n47), .A2(n87), .B1(n46), .B2(n37), .ZN(N289) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[1]), .ZN(n86) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[33]), .ZN(n38) );
  OAI22D1BWP30P140 U105 ( .A1(n47), .A2(n86), .B1(n46), .B2(n38), .ZN(N288) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[4]), .ZN(n89) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U108 ( .A1(n43), .A2(n89), .B1(n46), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[5]), .ZN(n90) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[37]), .ZN(n40) );
  OAI22D1BWP30P140 U111 ( .A1(n43), .A2(n90), .B1(n46), .B2(n40), .ZN(N292) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[6]), .ZN(n91) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[38]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n43), .A2(n91), .B1(n46), .B2(n41), .ZN(N293) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[7]), .ZN(n93) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[39]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n43), .A2(n93), .B1(n46), .B2(n42), .ZN(N294) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[0]), .ZN(n85) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[32]), .ZN(n44) );
  OAI22D1BWP30P140 U120 ( .A1(n47), .A2(n85), .B1(n46), .B2(n44), .ZN(N287) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[3]), .ZN(n88) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[35]), .ZN(n45) );
  OAI22D1BWP30P140 U123 ( .A1(n47), .A2(n88), .B1(n46), .B2(n45), .ZN(N290) );
  INVD1BWP30P140 U124 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U125 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n92) );
  OAI21D1BWP30P140 U127 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  MUX2NUD1BWP30P140 U128 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  INVD2BWP30P140 U129 ( .I(n84), .ZN(n82) );
  MOAI22D1BWP30P140 U130 ( .A1(n58), .A2(n82), .B1(i_data_bus[40]), .B2(n92), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U131 ( .A1(n59), .A2(n82), .B1(i_data_bus[41]), .B2(n92), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U132 ( .A1(n60), .A2(n82), .B1(i_data_bus[42]), .B2(n92), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U133 ( .A1(n61), .A2(n82), .B1(i_data_bus[43]), .B2(n92), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U134 ( .A1(n62), .A2(n82), .B1(i_data_bus[44]), .B2(n92), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U135 ( .A1(n63), .A2(n82), .B1(i_data_bus[45]), .B2(n92), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U136 ( .A1(n64), .A2(n82), .B1(i_data_bus[47]), .B2(n92), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U137 ( .A1(n65), .A2(n82), .B1(i_data_bus[48]), .B2(n92), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U138 ( .A1(n66), .A2(n82), .B1(i_data_bus[49]), .B2(n92), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U139 ( .A1(n67), .A2(n82), .B1(i_data_bus[50]), .B2(n92), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U140 ( .A1(n68), .A2(n82), .B1(i_data_bus[51]), .B2(n92), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U141 ( .A1(n69), .A2(n80), .B1(i_data_bus[52]), .B2(n92), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U142 ( .A1(n70), .A2(n80), .B1(i_data_bus[53]), .B2(n92), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U143 ( .A1(n71), .A2(n80), .B1(i_data_bus[54]), .B2(n92), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U144 ( .A1(n72), .A2(n80), .B1(i_data_bus[55]), .B2(n92), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U145 ( .A1(n73), .A2(n80), .B1(i_data_bus[56]), .B2(n92), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U146 ( .A1(n74), .A2(n80), .B1(i_data_bus[57]), .B2(n92), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U147 ( .A1(n75), .A2(n80), .B1(i_data_bus[58]), .B2(n92), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U148 ( .A1(n76), .A2(n80), .B1(i_data_bus[59]), .B2(n92), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U149 ( .A1(n77), .A2(n80), .B1(i_data_bus[60]), .B2(n92), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U150 ( .A1(n78), .A2(n80), .B1(i_data_bus[61]), .B2(n92), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U151 ( .A1(n79), .A2(n80), .B1(i_data_bus[62]), .B2(n92), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n80), .B1(i_data_bus[63]), .B2(n92), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n82), .B1(i_data_bus[46]), .B2(n92), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U154 ( .A1(n85), .A2(n1), .B1(i_data_bus[32]), .B2(n92), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U155 ( .A1(n86), .A2(n1), .B1(i_data_bus[33]), .B2(n92), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U156 ( .A1(n87), .A2(n1), .B1(i_data_bus[34]), .B2(n92), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U157 ( .A1(n88), .A2(n1), .B1(i_data_bus[35]), .B2(n92), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U158 ( .A1(n89), .A2(n1), .B1(i_data_bus[36]), .B2(n92), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U159 ( .A1(n90), .A2(n1), .B1(i_data_bus[37]), .B2(n92), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U160 ( .A1(n91), .A2(n1), .B1(i_data_bus[38]), .B2(n92), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n1), .B1(i_data_bus[39]), .B2(n92), 
        .ZN(N326) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_114 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n19), .A2(n18), .B1(n31), .B2(n70), .ZN(N306) );
  INVD2BWP30P140 U4 ( .I(n36), .ZN(n46) );
  OAI22D1BWP30P140 U5 ( .A1(n47), .A2(n85), .B1(n46), .B2(n45), .ZN(N287) );
  INVD1BWP30P140 U6 ( .I(n57), .ZN(n84) );
  ND2D1BWP30P140 U7 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U9 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U10 ( .I(n92), .ZN(n50) );
  OAI22D1BWP30P140 U11 ( .A1(n19), .A2(n7), .B1(n41), .B2(n58), .ZN(N295) );
  OAI22D1BWP30P140 U12 ( .A1(n19), .A2(n8), .B1(n41), .B2(n59), .ZN(N296) );
  OAI22D1BWP30P140 U13 ( .A1(n19), .A2(n9), .B1(n41), .B2(n60), .ZN(N297) );
  OAI22D1BWP30P140 U14 ( .A1(n19), .A2(n10), .B1(n41), .B2(n61), .ZN(N298) );
  OAI22D1BWP30P140 U15 ( .A1(n19), .A2(n11), .B1(n41), .B2(n62), .ZN(N299) );
  OAI22D1BWP30P140 U16 ( .A1(n19), .A2(n12), .B1(n41), .B2(n63), .ZN(N300) );
  OAI22D1BWP30P140 U17 ( .A1(n19), .A2(n13), .B1(n41), .B2(n64), .ZN(N301) );
  OAI22D1BWP30P140 U18 ( .A1(n19), .A2(n14), .B1(n41), .B2(n65), .ZN(N302) );
  OAI22D1BWP30P140 U19 ( .A1(n19), .A2(n15), .B1(n41), .B2(n66), .ZN(N303) );
  OAI22D1BWP30P140 U20 ( .A1(n19), .A2(n16), .B1(n41), .B2(n67), .ZN(N304) );
  OAI22D1BWP30P140 U21 ( .A1(n19), .A2(n17), .B1(n41), .B2(n68), .ZN(N305) );
  OAI22D1BWP30P140 U22 ( .A1(n33), .A2(n20), .B1(n31), .B2(n71), .ZN(N307) );
  OAI22D1BWP30P140 U23 ( .A1(n33), .A2(n21), .B1(n31), .B2(n72), .ZN(N308) );
  OAI22D1BWP30P140 U24 ( .A1(n33), .A2(n22), .B1(n31), .B2(n73), .ZN(N309) );
  OAI22D1BWP30P140 U25 ( .A1(n33), .A2(n23), .B1(n31), .B2(n74), .ZN(N310) );
  OAI22D1BWP30P140 U26 ( .A1(n33), .A2(n24), .B1(n31), .B2(n75), .ZN(N311) );
  OAI22D1BWP30P140 U27 ( .A1(n33), .A2(n25), .B1(n31), .B2(n76), .ZN(N312) );
  OAI22D1BWP30P140 U28 ( .A1(n33), .A2(n26), .B1(n31), .B2(n77), .ZN(N313) );
  OAI22D1BWP30P140 U29 ( .A1(n33), .A2(n27), .B1(n31), .B2(n78), .ZN(N314) );
  OAI22D1BWP30P140 U30 ( .A1(n33), .A2(n28), .B1(n31), .B2(n79), .ZN(N315) );
  OAI22D1BWP30P140 U31 ( .A1(n33), .A2(n29), .B1(n31), .B2(n80), .ZN(N316) );
  OAI22D1BWP30P140 U32 ( .A1(n33), .A2(n30), .B1(n31), .B2(n81), .ZN(N317) );
  OAI22D1BWP30P140 U33 ( .A1(n33), .A2(n32), .B1(n31), .B2(n83), .ZN(N318) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n19) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n41) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n58) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n59) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n60) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n61) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n62) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n63) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[14]), .ZN(n64) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[47]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[15]), .ZN(n65) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[48]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n66) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n67) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n68) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n18) );
  INVD2BWP30P140 U70 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n70) );
  INVD2BWP30P140 U72 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n20) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n71) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n21) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n72) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n22) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n73) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n23) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n74) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n75) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n76) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n77) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n78) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n79) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n80) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n30) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n81) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n83) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n47) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n47), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n93) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[39]), .ZN(n37) );
  OAI22D1BWP30P140 U101 ( .A1(n41), .A2(n93), .B1(n46), .B2(n37), .ZN(N294) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[6]), .ZN(n91) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[38]), .ZN(n38) );
  OAI22D1BWP30P140 U104 ( .A1(n41), .A2(n91), .B1(n46), .B2(n38), .ZN(N293) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[5]), .ZN(n90) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[37]), .ZN(n39) );
  OAI22D1BWP30P140 U107 ( .A1(n41), .A2(n90), .B1(n46), .B2(n39), .ZN(N292) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[4]), .ZN(n89) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[36]), .ZN(n40) );
  OAI22D1BWP30P140 U110 ( .A1(n41), .A2(n89), .B1(n46), .B2(n40), .ZN(N291) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[3]), .ZN(n88) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[35]), .ZN(n42) );
  OAI22D1BWP30P140 U113 ( .A1(n47), .A2(n88), .B1(n46), .B2(n42), .ZN(N290) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[2]), .ZN(n87) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[34]), .ZN(n43) );
  OAI22D1BWP30P140 U116 ( .A1(n47), .A2(n87), .B1(n46), .B2(n43), .ZN(N289) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[1]), .ZN(n86) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[33]), .ZN(n44) );
  OAI22D1BWP30P140 U119 ( .A1(n47), .A2(n86), .B1(n46), .B2(n44), .ZN(N288) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[0]), .ZN(n85) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[32]), .ZN(n45) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n92) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  INVD2BWP30P140 U128 ( .I(n84), .ZN(n69) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n69), .B1(i_data_bus[40]), .B2(n92), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n69), .B1(i_data_bus[41]), .B2(n92), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n69), .B1(i_data_bus[42]), .B2(n92), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n69), .B1(i_data_bus[43]), .B2(n92), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n69), .B1(i_data_bus[44]), .B2(n92), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n69), .B1(i_data_bus[45]), .B2(n92), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n69), .B1(i_data_bus[46]), .B2(n92), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n69), .B1(i_data_bus[47]), .B2(n92), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n69), .B1(i_data_bus[48]), .B2(n92), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n69), .B1(i_data_bus[49]), .B2(n92), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n69), .B1(i_data_bus[50]), .B2(n92), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U140 ( .A1(n70), .A2(n69), .B1(i_data_bus[51]), .B2(n92), 
        .ZN(N338) );
  INVD2BWP30P140 U141 ( .I(n84), .ZN(n82) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n82), .B1(i_data_bus[52]), .B2(n92), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n82), .B1(i_data_bus[53]), .B2(n92), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n82), .B1(i_data_bus[54]), .B2(n92), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n82), .B1(i_data_bus[55]), .B2(n92), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n82), .B1(i_data_bus[56]), .B2(n92), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n82), .B1(i_data_bus[57]), .B2(n92), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n82), .B1(i_data_bus[58]), .B2(n92), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n82), .B1(i_data_bus[59]), .B2(n92), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n82), .B1(i_data_bus[60]), .B2(n92), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n82), .B1(i_data_bus[61]), .B2(n92), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n82), .B1(i_data_bus[62]), .B2(n92), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n82), .B1(i_data_bus[63]), .B2(n92), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U154 ( .A1(n85), .A2(n1), .B1(i_data_bus[32]), .B2(n92), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U155 ( .A1(n86), .A2(n1), .B1(i_data_bus[33]), .B2(n92), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U156 ( .A1(n87), .A2(n1), .B1(i_data_bus[34]), .B2(n92), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U157 ( .A1(n88), .A2(n1), .B1(i_data_bus[35]), .B2(n92), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U158 ( .A1(n89), .A2(n1), .B1(i_data_bus[36]), .B2(n92), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U159 ( .A1(n90), .A2(n1), .B1(i_data_bus[37]), .B2(n92), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U160 ( .A1(n91), .A2(n1), .B1(i_data_bus[38]), .B2(n92), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n1), .B1(i_data_bus[39]), .B2(n92), 
        .ZN(N326) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_115 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD1BWP30P140 U3 ( .I(n57), .ZN(n84) );
  INVD2BWP30P140 U4 ( .I(n84), .ZN(n82) );
  NR2D1BWP30P140 U5 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  OAI22D1BWP30P140 U6 ( .A1(n19), .A2(n7), .B1(n41), .B2(n58), .ZN(N295) );
  OAI22D1BWP30P140 U7 ( .A1(n19), .A2(n8), .B1(n41), .B2(n59), .ZN(N296) );
  OAI22D1BWP30P140 U8 ( .A1(n19), .A2(n9), .B1(n41), .B2(n60), .ZN(N297) );
  OAI22D1BWP30P140 U9 ( .A1(n19), .A2(n10), .B1(n41), .B2(n61), .ZN(N298) );
  OAI22D1BWP30P140 U10 ( .A1(n19), .A2(n11), .B1(n41), .B2(n62), .ZN(N299) );
  OAI22D1BWP30P140 U11 ( .A1(n19), .A2(n12), .B1(n41), .B2(n63), .ZN(N300) );
  OAI22D1BWP30P140 U12 ( .A1(n19), .A2(n13), .B1(n41), .B2(n64), .ZN(N301) );
  OAI22D1BWP30P140 U13 ( .A1(n19), .A2(n14), .B1(n41), .B2(n65), .ZN(N302) );
  OAI22D1BWP30P140 U14 ( .A1(n19), .A2(n15), .B1(n41), .B2(n66), .ZN(N303) );
  OAI22D1BWP30P140 U15 ( .A1(n19), .A2(n16), .B1(n41), .B2(n67), .ZN(N304) );
  OAI22D1BWP30P140 U16 ( .A1(n19), .A2(n17), .B1(n41), .B2(n68), .ZN(N305) );
  OAI22D1BWP30P140 U17 ( .A1(n33), .A2(n20), .B1(n31), .B2(n71), .ZN(N307) );
  OAI22D1BWP30P140 U18 ( .A1(n33), .A2(n21), .B1(n31), .B2(n72), .ZN(N308) );
  OAI22D1BWP30P140 U19 ( .A1(n33), .A2(n22), .B1(n31), .B2(n73), .ZN(N309) );
  OAI22D1BWP30P140 U20 ( .A1(n33), .A2(n23), .B1(n31), .B2(n74), .ZN(N310) );
  OAI22D1BWP30P140 U21 ( .A1(n33), .A2(n24), .B1(n31), .B2(n75), .ZN(N311) );
  OAI22D1BWP30P140 U22 ( .A1(n33), .A2(n25), .B1(n31), .B2(n76), .ZN(N312) );
  OAI22D1BWP30P140 U23 ( .A1(n33), .A2(n26), .B1(n31), .B2(n77), .ZN(N313) );
  OAI22D1BWP30P140 U24 ( .A1(n33), .A2(n27), .B1(n31), .B2(n78), .ZN(N314) );
  OAI22D1BWP30P140 U25 ( .A1(n33), .A2(n28), .B1(n31), .B2(n79), .ZN(N315) );
  OAI22D1BWP30P140 U26 ( .A1(n33), .A2(n29), .B1(n31), .B2(n80), .ZN(N316) );
  OAI22D1BWP30P140 U27 ( .A1(n33), .A2(n30), .B1(n31), .B2(n81), .ZN(N317) );
  OAI22D1BWP30P140 U28 ( .A1(n33), .A2(n32), .B1(n31), .B2(n83), .ZN(N318) );
  ND2D1BWP30P140 U29 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U30 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U31 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U32 ( .I(n92), .ZN(n50) );
  OAI22D1BWP30P140 U33 ( .A1(n19), .A2(n18), .B1(n31), .B2(n70), .ZN(N306) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n19) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n41) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n58) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n59) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n60) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n61) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n62) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n63) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[14]), .ZN(n64) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[47]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[15]), .ZN(n65) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[48]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n66) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n67) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n68) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n18) );
  INVD2BWP30P140 U70 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n70) );
  INVD2BWP30P140 U72 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n20) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n71) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n21) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n72) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n22) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n73) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n23) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n74) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n75) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n76) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n77) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n78) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n79) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n80) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n30) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n81) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n83) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n47) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n47), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n93) );
  INVD2BWP30P140 U100 ( .I(n36), .ZN(n46) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n37) );
  OAI22D1BWP30P140 U102 ( .A1(n41), .A2(n93), .B1(n46), .B2(n37), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[6]), .ZN(n91) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[38]), .ZN(n38) );
  OAI22D1BWP30P140 U105 ( .A1(n41), .A2(n91), .B1(n46), .B2(n38), .ZN(N293) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[5]), .ZN(n90) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[37]), .ZN(n39) );
  OAI22D1BWP30P140 U108 ( .A1(n41), .A2(n90), .B1(n46), .B2(n39), .ZN(N292) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n89) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n40) );
  OAI22D1BWP30P140 U111 ( .A1(n41), .A2(n89), .B1(n46), .B2(n40), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n88) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n42) );
  OAI22D1BWP30P140 U114 ( .A1(n47), .A2(n88), .B1(n46), .B2(n42), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n87) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n43) );
  OAI22D1BWP30P140 U117 ( .A1(n47), .A2(n87), .B1(n46), .B2(n43), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n86) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n44) );
  OAI22D1BWP30P140 U120 ( .A1(n47), .A2(n86), .B1(n46), .B2(n44), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n85) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n45) );
  OAI22D1BWP30P140 U123 ( .A1(n47), .A2(n85), .B1(n46), .B2(n45), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U125 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n92) );
  OAI21D1BWP30P140 U127 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  MUX2NUD1BWP30P140 U128 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  INVD2BWP30P140 U129 ( .I(n84), .ZN(n69) );
  MOAI22D1BWP30P140 U130 ( .A1(n58), .A2(n69), .B1(i_data_bus[40]), .B2(n92), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U131 ( .A1(n59), .A2(n69), .B1(i_data_bus[41]), .B2(n92), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U132 ( .A1(n60), .A2(n69), .B1(i_data_bus[42]), .B2(n92), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U133 ( .A1(n61), .A2(n69), .B1(i_data_bus[43]), .B2(n92), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U134 ( .A1(n62), .A2(n69), .B1(i_data_bus[44]), .B2(n92), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U135 ( .A1(n63), .A2(n69), .B1(i_data_bus[45]), .B2(n92), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U136 ( .A1(n64), .A2(n69), .B1(i_data_bus[46]), .B2(n92), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U137 ( .A1(n65), .A2(n69), .B1(i_data_bus[47]), .B2(n92), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U138 ( .A1(n66), .A2(n69), .B1(i_data_bus[48]), .B2(n92), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U139 ( .A1(n67), .A2(n69), .B1(i_data_bus[49]), .B2(n92), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U140 ( .A1(n68), .A2(n69), .B1(i_data_bus[50]), .B2(n92), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n69), .B1(i_data_bus[51]), .B2(n92), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n82), .B1(i_data_bus[52]), .B2(n92), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n82), .B1(i_data_bus[53]), .B2(n92), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n82), .B1(i_data_bus[54]), .B2(n92), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n82), .B1(i_data_bus[55]), .B2(n92), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n82), .B1(i_data_bus[56]), .B2(n92), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n82), .B1(i_data_bus[57]), .B2(n92), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n82), .B1(i_data_bus[58]), .B2(n92), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n82), .B1(i_data_bus[59]), .B2(n92), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n82), .B1(i_data_bus[60]), .B2(n92), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n82), .B1(i_data_bus[61]), .B2(n92), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n82), .B1(i_data_bus[62]), .B2(n92), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n82), .B1(i_data_bus[63]), .B2(n92), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U154 ( .A1(n85), .A2(n1), .B1(i_data_bus[32]), .B2(n92), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U155 ( .A1(n86), .A2(n1), .B1(i_data_bus[33]), .B2(n92), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U156 ( .A1(n87), .A2(n1), .B1(i_data_bus[34]), .B2(n92), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U157 ( .A1(n88), .A2(n1), .B1(i_data_bus[35]), .B2(n92), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U158 ( .A1(n89), .A2(n1), .B1(i_data_bus[36]), .B2(n92), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U159 ( .A1(n90), .A2(n1), .B1(i_data_bus[37]), .B2(n92), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U160 ( .A1(n91), .A2(n1), .B1(i_data_bus[38]), .B2(n92), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n1), .B1(i_data_bus[39]), .B2(n92), 
        .ZN(N326) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_116 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n22), .A2(n21), .B1(n31), .B2(n63), .ZN(N306) );
  INVD2BWP30P140 U4 ( .I(n36), .ZN(n46) );
  OAI22D1BWP30P140 U5 ( .A1(n47), .A2(n85), .B1(n46), .B2(n45), .ZN(N287) );
  INVD1BWP30P140 U6 ( .I(n57), .ZN(n84) );
  ND2D1BWP30P140 U7 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U9 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U10 ( .I(n92), .ZN(n50) );
  OAI22D1BWP30P140 U11 ( .A1(n22), .A2(n7), .B1(n41), .B2(n83), .ZN(N295) );
  OAI22D1BWP30P140 U12 ( .A1(n22), .A2(n8), .B1(n41), .B2(n75), .ZN(N296) );
  OAI22D1BWP30P140 U13 ( .A1(n22), .A2(n9), .B1(n41), .B2(n74), .ZN(N297) );
  OAI22D1BWP30P140 U14 ( .A1(n22), .A2(n10), .B1(n41), .B2(n73), .ZN(N298) );
  OAI22D1BWP30P140 U15 ( .A1(n22), .A2(n11), .B1(n41), .B2(n72), .ZN(N299) );
  OAI22D1BWP30P140 U16 ( .A1(n22), .A2(n12), .B1(n41), .B2(n66), .ZN(N300) );
  OAI22D1BWP30P140 U17 ( .A1(n22), .A2(n13), .B1(n41), .B2(n67), .ZN(N301) );
  OAI22D1BWP30P140 U18 ( .A1(n22), .A2(n14), .B1(n41), .B2(n68), .ZN(N302) );
  OAI22D1BWP30P140 U19 ( .A1(n22), .A2(n15), .B1(n41), .B2(n76), .ZN(N303) );
  OAI22D1BWP30P140 U20 ( .A1(n22), .A2(n16), .B1(n41), .B2(n58), .ZN(N304) );
  OAI22D1BWP30P140 U21 ( .A1(n22), .A2(n17), .B1(n41), .B2(n59), .ZN(N305) );
  OAI22D1BWP30P140 U22 ( .A1(n33), .A2(n23), .B1(n31), .B2(n61), .ZN(N307) );
  OAI22D1BWP30P140 U23 ( .A1(n33), .A2(n24), .B1(n31), .B2(n62), .ZN(N308) );
  OAI22D1BWP30P140 U24 ( .A1(n33), .A2(n25), .B1(n31), .B2(n81), .ZN(N309) );
  OAI22D1BWP30P140 U25 ( .A1(n33), .A2(n26), .B1(n31), .B2(n64), .ZN(N310) );
  OAI22D1BWP30P140 U26 ( .A1(n33), .A2(n27), .B1(n31), .B2(n60), .ZN(N311) );
  OAI22D1BWP30P140 U27 ( .A1(n33), .A2(n28), .B1(n31), .B2(n69), .ZN(N312) );
  OAI22D1BWP30P140 U28 ( .A1(n33), .A2(n29), .B1(n31), .B2(n70), .ZN(N313) );
  OAI22D1BWP30P140 U29 ( .A1(n33), .A2(n30), .B1(n31), .B2(n71), .ZN(N314) );
  OAI22D1BWP30P140 U30 ( .A1(n33), .A2(n32), .B1(n31), .B2(n65), .ZN(N315) );
  OAI22D1BWP30P140 U31 ( .A1(n33), .A2(n20), .B1(n31), .B2(n77), .ZN(N316) );
  OAI22D1BWP30P140 U32 ( .A1(n33), .A2(n19), .B1(n31), .B2(n78), .ZN(N317) );
  OAI22D1BWP30P140 U33 ( .A1(n33), .A2(n18), .B1(n31), .B2(n79), .ZN(N318) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n22) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n41) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n83) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n75) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n74) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n73) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n72) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n66) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[14]), .ZN(n67) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[47]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[15]), .ZN(n68) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[48]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n76) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n58) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n59) );
  INVD2BWP30P140 U69 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[63]), .ZN(n18) );
  INVD2BWP30P140 U71 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[31]), .ZN(n79) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[62]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[30]), .ZN(n78) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[61]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[29]), .ZN(n77) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[51]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[19]), .ZN(n63) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[52]), .ZN(n23) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[20]), .ZN(n61) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[53]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[21]), .ZN(n62) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[54]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[22]), .ZN(n81) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[55]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[23]), .ZN(n64) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[56]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[24]), .ZN(n60) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[57]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[25]), .ZN(n69) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[58]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[26]), .ZN(n70) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[59]), .ZN(n30) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[27]), .ZN(n71) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[60]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[28]), .ZN(n65) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n47) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n47), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n93) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[39]), .ZN(n37) );
  OAI22D1BWP30P140 U101 ( .A1(n41), .A2(n93), .B1(n46), .B2(n37), .ZN(N294) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[6]), .ZN(n91) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[38]), .ZN(n38) );
  OAI22D1BWP30P140 U104 ( .A1(n41), .A2(n91), .B1(n46), .B2(n38), .ZN(N293) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[5]), .ZN(n90) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[37]), .ZN(n39) );
  OAI22D1BWP30P140 U107 ( .A1(n41), .A2(n90), .B1(n46), .B2(n39), .ZN(N292) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[4]), .ZN(n89) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[36]), .ZN(n40) );
  OAI22D1BWP30P140 U110 ( .A1(n41), .A2(n89), .B1(n46), .B2(n40), .ZN(N291) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[3]), .ZN(n88) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[35]), .ZN(n42) );
  OAI22D1BWP30P140 U113 ( .A1(n47), .A2(n88), .B1(n46), .B2(n42), .ZN(N290) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[2]), .ZN(n87) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[34]), .ZN(n43) );
  OAI22D1BWP30P140 U116 ( .A1(n47), .A2(n87), .B1(n46), .B2(n43), .ZN(N289) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[1]), .ZN(n86) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[33]), .ZN(n44) );
  OAI22D1BWP30P140 U119 ( .A1(n47), .A2(n86), .B1(n46), .B2(n44), .ZN(N288) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[0]), .ZN(n85) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[32]), .ZN(n45) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n92) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  INVD2BWP30P140 U128 ( .I(n84), .ZN(n82) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n82), .B1(i_data_bus[49]), .B2(n92), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n82), .B1(i_data_bus[50]), .B2(n92), 
        .ZN(N337) );
  INVD2BWP30P140 U131 ( .I(n84), .ZN(n80) );
  MOAI22D1BWP30P140 U132 ( .A1(n60), .A2(n80), .B1(i_data_bus[56]), .B2(n92), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U133 ( .A1(n61), .A2(n80), .B1(i_data_bus[52]), .B2(n92), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U134 ( .A1(n62), .A2(n80), .B1(i_data_bus[53]), .B2(n92), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U135 ( .A1(n63), .A2(n82), .B1(i_data_bus[51]), .B2(n92), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U136 ( .A1(n64), .A2(n80), .B1(i_data_bus[55]), .B2(n92), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U137 ( .A1(n65), .A2(n80), .B1(i_data_bus[60]), .B2(n92), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U138 ( .A1(n66), .A2(n82), .B1(i_data_bus[45]), .B2(n92), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U139 ( .A1(n67), .A2(n82), .B1(i_data_bus[46]), .B2(n92), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U140 ( .A1(n68), .A2(n82), .B1(i_data_bus[47]), .B2(n92), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U141 ( .A1(n69), .A2(n80), .B1(i_data_bus[57]), .B2(n92), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U142 ( .A1(n70), .A2(n80), .B1(i_data_bus[58]), .B2(n92), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U143 ( .A1(n71), .A2(n80), .B1(i_data_bus[59]), .B2(n92), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U144 ( .A1(n72), .A2(n82), .B1(i_data_bus[44]), .B2(n92), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U145 ( .A1(n73), .A2(n82), .B1(i_data_bus[43]), .B2(n92), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U146 ( .A1(n74), .A2(n82), .B1(i_data_bus[42]), .B2(n92), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U147 ( .A1(n75), .A2(n82), .B1(i_data_bus[41]), .B2(n92), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U148 ( .A1(n76), .A2(n82), .B1(i_data_bus[48]), .B2(n92), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U149 ( .A1(n77), .A2(n80), .B1(i_data_bus[61]), .B2(n92), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U150 ( .A1(n78), .A2(n80), .B1(i_data_bus[62]), .B2(n92), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U151 ( .A1(n79), .A2(n80), .B1(i_data_bus[63]), .B2(n92), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n80), .B1(i_data_bus[54]), .B2(n92), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n82), .B1(i_data_bus[40]), .B2(n92), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U154 ( .A1(n85), .A2(n1), .B1(i_data_bus[32]), .B2(n92), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U155 ( .A1(n86), .A2(n1), .B1(i_data_bus[33]), .B2(n92), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U156 ( .A1(n87), .A2(n1), .B1(i_data_bus[34]), .B2(n92), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U157 ( .A1(n88), .A2(n1), .B1(i_data_bus[35]), .B2(n92), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U158 ( .A1(n89), .A2(n1), .B1(i_data_bus[36]), .B2(n92), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U159 ( .A1(n90), .A2(n1), .B1(i_data_bus[37]), .B2(n92), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U160 ( .A1(n91), .A2(n1), .B1(i_data_bus[38]), .B2(n92), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n1), .B1(i_data_bus[39]), .B2(n92), 
        .ZN(N326) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_117 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD1BWP30P140 U3 ( .I(n57), .ZN(n84) );
  INVD2BWP30P140 U4 ( .I(n84), .ZN(n82) );
  NR2D1BWP30P140 U5 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  OAI22D1BWP30P140 U6 ( .A1(n19), .A2(n7), .B1(n47), .B2(n83), .ZN(N295) );
  OAI22D1BWP30P140 U7 ( .A1(n19), .A2(n8), .B1(n47), .B2(n81), .ZN(N296) );
  OAI22D1BWP30P140 U8 ( .A1(n19), .A2(n9), .B1(n47), .B2(n80), .ZN(N297) );
  OAI22D1BWP30P140 U9 ( .A1(n19), .A2(n10), .B1(n47), .B2(n79), .ZN(N298) );
  OAI22D1BWP30P140 U10 ( .A1(n19), .A2(n11), .B1(n47), .B2(n78), .ZN(N299) );
  OAI22D1BWP30P140 U11 ( .A1(n19), .A2(n12), .B1(n47), .B2(n77), .ZN(N300) );
  OAI22D1BWP30P140 U12 ( .A1(n19), .A2(n13), .B1(n47), .B2(n76), .ZN(N301) );
  OAI22D1BWP30P140 U13 ( .A1(n19), .A2(n14), .B1(n47), .B2(n75), .ZN(N302) );
  OAI22D1BWP30P140 U14 ( .A1(n19), .A2(n15), .B1(n47), .B2(n74), .ZN(N303) );
  OAI22D1BWP30P140 U15 ( .A1(n19), .A2(n16), .B1(n47), .B2(n73), .ZN(N304) );
  OAI22D1BWP30P140 U16 ( .A1(n19), .A2(n17), .B1(n47), .B2(n72), .ZN(N305) );
  OAI22D1BWP30P140 U17 ( .A1(n33), .A2(n20), .B1(n31), .B2(n70), .ZN(N307) );
  OAI22D1BWP30P140 U18 ( .A1(n33), .A2(n21), .B1(n31), .B2(n68), .ZN(N308) );
  OAI22D1BWP30P140 U19 ( .A1(n33), .A2(n22), .B1(n31), .B2(n67), .ZN(N309) );
  OAI22D1BWP30P140 U20 ( .A1(n33), .A2(n23), .B1(n31), .B2(n66), .ZN(N310) );
  OAI22D1BWP30P140 U21 ( .A1(n33), .A2(n24), .B1(n31), .B2(n65), .ZN(N311) );
  OAI22D1BWP30P140 U22 ( .A1(n33), .A2(n25), .B1(n31), .B2(n64), .ZN(N312) );
  OAI22D1BWP30P140 U23 ( .A1(n33), .A2(n26), .B1(n31), .B2(n63), .ZN(N313) );
  OAI22D1BWP30P140 U24 ( .A1(n33), .A2(n27), .B1(n31), .B2(n62), .ZN(N314) );
  OAI22D1BWP30P140 U25 ( .A1(n33), .A2(n28), .B1(n31), .B2(n61), .ZN(N315) );
  OAI22D1BWP30P140 U26 ( .A1(n33), .A2(n29), .B1(n31), .B2(n60), .ZN(N316) );
  OAI22D1BWP30P140 U27 ( .A1(n33), .A2(n30), .B1(n31), .B2(n59), .ZN(N317) );
  OAI22D1BWP30P140 U28 ( .A1(n33), .A2(n32), .B1(n31), .B2(n58), .ZN(N318) );
  ND2D1BWP30P140 U29 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U30 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U31 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U32 ( .I(n92), .ZN(n50) );
  OAI22D1BWP30P140 U33 ( .A1(n19), .A2(n18), .B1(n31), .B2(n71), .ZN(N306) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n19) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n47) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n83) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n81) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n80) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n79) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n78) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n77) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[14]), .ZN(n76) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[47]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[15]), .ZN(n75) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[48]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n74) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n73) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n72) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n18) );
  INVD2BWP30P140 U70 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n71) );
  INVD2BWP30P140 U72 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n20) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n70) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n21) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n68) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n22) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n67) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n23) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n66) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n65) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n64) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n63) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n62) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n61) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n60) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n30) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n59) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n58) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n43) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n43), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[1]), .ZN(n86) );
  INVD2BWP30P140 U100 ( .I(n36), .ZN(n46) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[33]), .ZN(n37) );
  OAI22D1BWP30P140 U102 ( .A1(n43), .A2(n86), .B1(n46), .B2(n37), .ZN(N288) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[0]), .ZN(n85) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[32]), .ZN(n38) );
  OAI22D1BWP30P140 U105 ( .A1(n43), .A2(n85), .B1(n46), .B2(n38), .ZN(N287) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[6]), .ZN(n91) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[38]), .ZN(n39) );
  OAI22D1BWP30P140 U108 ( .A1(n47), .A2(n91), .B1(n46), .B2(n39), .ZN(N293) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[7]), .ZN(n93) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[39]), .ZN(n40) );
  OAI22D1BWP30P140 U111 ( .A1(n47), .A2(n93), .B1(n46), .B2(n40), .ZN(N294) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n88) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n43), .A2(n88), .B1(n46), .B2(n41), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n87) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n43), .A2(n87), .B1(n46), .B2(n42), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[4]), .ZN(n89) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[36]), .ZN(n44) );
  OAI22D1BWP30P140 U120 ( .A1(n47), .A2(n89), .B1(n46), .B2(n44), .ZN(N291) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[5]), .ZN(n90) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[37]), .ZN(n45) );
  OAI22D1BWP30P140 U123 ( .A1(n47), .A2(n90), .B1(n46), .B2(n45), .ZN(N292) );
  INVD1BWP30P140 U124 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U125 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n92) );
  OAI21D1BWP30P140 U127 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  MUX2NUD1BWP30P140 U128 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  INVD2BWP30P140 U129 ( .I(n84), .ZN(n69) );
  MOAI22D1BWP30P140 U130 ( .A1(n58), .A2(n69), .B1(i_data_bus[63]), .B2(n92), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U131 ( .A1(n59), .A2(n69), .B1(i_data_bus[62]), .B2(n92), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U132 ( .A1(n60), .A2(n69), .B1(i_data_bus[61]), .B2(n92), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U133 ( .A1(n61), .A2(n69), .B1(i_data_bus[60]), .B2(n92), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U134 ( .A1(n62), .A2(n69), .B1(i_data_bus[59]), .B2(n92), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U135 ( .A1(n63), .A2(n69), .B1(i_data_bus[58]), .B2(n92), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U136 ( .A1(n64), .A2(n69), .B1(i_data_bus[57]), .B2(n92), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U137 ( .A1(n65), .A2(n69), .B1(i_data_bus[56]), .B2(n92), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U138 ( .A1(n66), .A2(n69), .B1(i_data_bus[55]), .B2(n92), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U139 ( .A1(n67), .A2(n69), .B1(i_data_bus[54]), .B2(n92), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U140 ( .A1(n68), .A2(n69), .B1(i_data_bus[53]), .B2(n92), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n69), .B1(i_data_bus[52]), .B2(n92), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n82), .B1(i_data_bus[51]), .B2(n92), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n82), .B1(i_data_bus[50]), .B2(n92), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n82), .B1(i_data_bus[49]), .B2(n92), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n82), .B1(i_data_bus[48]), .B2(n92), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n82), .B1(i_data_bus[47]), .B2(n92), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n82), .B1(i_data_bus[46]), .B2(n92), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n82), .B1(i_data_bus[45]), .B2(n92), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n82), .B1(i_data_bus[44]), .B2(n92), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n82), .B1(i_data_bus[43]), .B2(n92), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n82), .B1(i_data_bus[42]), .B2(n92), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n82), .B1(i_data_bus[41]), .B2(n92), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n82), .B1(i_data_bus[40]), .B2(n92), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U154 ( .A1(n85), .A2(n1), .B1(i_data_bus[32]), .B2(n92), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U155 ( .A1(n86), .A2(n1), .B1(i_data_bus[33]), .B2(n92), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U156 ( .A1(n87), .A2(n1), .B1(i_data_bus[34]), .B2(n92), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U157 ( .A1(n88), .A2(n1), .B1(i_data_bus[35]), .B2(n92), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U158 ( .A1(n89), .A2(n1), .B1(i_data_bus[36]), .B2(n92), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U159 ( .A1(n90), .A2(n1), .B1(i_data_bus[37]), .B2(n92), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U160 ( .A1(n91), .A2(n1), .B1(i_data_bus[38]), .B2(n92), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n1), .B1(i_data_bus[39]), .B2(n92), 
        .ZN(N326) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_118 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n19), .A2(n18), .B1(n31), .B2(n71), .ZN(N306) );
  INVD2BWP30P140 U4 ( .I(n36), .ZN(n46) );
  OAI22D1BWP30P140 U5 ( .A1(n44), .A2(n88), .B1(n46), .B2(n43), .ZN(N290) );
  INVD1BWP30P140 U6 ( .I(n57), .ZN(n84) );
  ND2D1BWP30P140 U7 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U9 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U10 ( .I(n92), .ZN(n50) );
  OAI22D1BWP30P140 U11 ( .A1(n19), .A2(n17), .B1(n47), .B2(n83), .ZN(N295) );
  OAI22D1BWP30P140 U12 ( .A1(n19), .A2(n16), .B1(n47), .B2(n81), .ZN(N296) );
  OAI22D1BWP30P140 U13 ( .A1(n19), .A2(n15), .B1(n47), .B2(n80), .ZN(N297) );
  OAI22D1BWP30P140 U14 ( .A1(n19), .A2(n14), .B1(n47), .B2(n79), .ZN(N298) );
  OAI22D1BWP30P140 U15 ( .A1(n19), .A2(n13), .B1(n47), .B2(n78), .ZN(N299) );
  OAI22D1BWP30P140 U16 ( .A1(n19), .A2(n12), .B1(n47), .B2(n77), .ZN(N300) );
  OAI22D1BWP30P140 U17 ( .A1(n19), .A2(n11), .B1(n47), .B2(n76), .ZN(N301) );
  OAI22D1BWP30P140 U18 ( .A1(n19), .A2(n7), .B1(n47), .B2(n75), .ZN(N302) );
  OAI22D1BWP30P140 U19 ( .A1(n19), .A2(n8), .B1(n47), .B2(n74), .ZN(N303) );
  OAI22D1BWP30P140 U20 ( .A1(n19), .A2(n9), .B1(n47), .B2(n73), .ZN(N304) );
  OAI22D1BWP30P140 U21 ( .A1(n19), .A2(n10), .B1(n47), .B2(n72), .ZN(N305) );
  OAI22D1BWP30P140 U22 ( .A1(n33), .A2(n20), .B1(n31), .B2(n70), .ZN(N307) );
  OAI22D1BWP30P140 U23 ( .A1(n33), .A2(n21), .B1(n31), .B2(n68), .ZN(N308) );
  OAI22D1BWP30P140 U24 ( .A1(n33), .A2(n22), .B1(n31), .B2(n67), .ZN(N309) );
  OAI22D1BWP30P140 U25 ( .A1(n33), .A2(n23), .B1(n31), .B2(n66), .ZN(N310) );
  OAI22D1BWP30P140 U26 ( .A1(n33), .A2(n24), .B1(n31), .B2(n65), .ZN(N311) );
  OAI22D1BWP30P140 U27 ( .A1(n33), .A2(n25), .B1(n31), .B2(n64), .ZN(N312) );
  OAI22D1BWP30P140 U28 ( .A1(n33), .A2(n26), .B1(n31), .B2(n63), .ZN(N313) );
  OAI22D1BWP30P140 U29 ( .A1(n33), .A2(n27), .B1(n31), .B2(n62), .ZN(N314) );
  OAI22D1BWP30P140 U30 ( .A1(n33), .A2(n28), .B1(n31), .B2(n61), .ZN(N315) );
  OAI22D1BWP30P140 U31 ( .A1(n33), .A2(n29), .B1(n31), .B2(n60), .ZN(N316) );
  OAI22D1BWP30P140 U32 ( .A1(n33), .A2(n30), .B1(n31), .B2(n59), .ZN(N317) );
  OAI22D1BWP30P140 U33 ( .A1(n33), .A2(n32), .B1(n31), .B2(n58), .ZN(N318) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n19) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[47]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n47) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[15]), .ZN(n75) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[48]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[16]), .ZN(n74) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[49]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[17]), .ZN(n73) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[50]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[18]), .ZN(n72) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[46]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[14]), .ZN(n76) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n77) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[44]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[12]), .ZN(n78) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[43]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[11]), .ZN(n79) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[42]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[10]), .ZN(n80) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[41]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[9]), .ZN(n81) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[40]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[8]), .ZN(n83) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n18) );
  INVD2BWP30P140 U70 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n71) );
  INVD2BWP30P140 U72 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n20) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n70) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n21) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n68) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n22) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n67) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n23) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n66) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n65) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n64) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n63) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n62) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n61) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n60) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n30) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n59) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n58) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n44) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n44), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[2]), .ZN(n87) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[34]), .ZN(n37) );
  OAI22D1BWP30P140 U101 ( .A1(n44), .A2(n87), .B1(n46), .B2(n37), .ZN(N289) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[0]), .ZN(n85) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[32]), .ZN(n38) );
  OAI22D1BWP30P140 U104 ( .A1(n44), .A2(n85), .B1(n46), .B2(n38), .ZN(N287) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[6]), .ZN(n91) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[38]), .ZN(n39) );
  OAI22D1BWP30P140 U107 ( .A1(n47), .A2(n91), .B1(n46), .B2(n39), .ZN(N293) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[1]), .ZN(n86) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[33]), .ZN(n40) );
  OAI22D1BWP30P140 U110 ( .A1(n44), .A2(n86), .B1(n46), .B2(n40), .ZN(N288) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[5]), .ZN(n90) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[37]), .ZN(n41) );
  OAI22D1BWP30P140 U113 ( .A1(n47), .A2(n90), .B1(n46), .B2(n41), .ZN(N292) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[7]), .ZN(n93) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[39]), .ZN(n42) );
  OAI22D1BWP30P140 U116 ( .A1(n47), .A2(n93), .B1(n46), .B2(n42), .ZN(N294) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[3]), .ZN(n88) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[35]), .ZN(n43) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[4]), .ZN(n89) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[36]), .ZN(n45) );
  OAI22D1BWP30P140 U121 ( .A1(n47), .A2(n89), .B1(n46), .B2(n45), .ZN(N291) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n92) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  INVD2BWP30P140 U128 ( .I(n84), .ZN(n69) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n69), .B1(i_data_bus[63]), .B2(n92), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n69), .B1(i_data_bus[62]), .B2(n92), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n69), .B1(i_data_bus[61]), .B2(n92), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n69), .B1(i_data_bus[60]), .B2(n92), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n69), .B1(i_data_bus[59]), .B2(n92), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n69), .B1(i_data_bus[58]), .B2(n92), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n69), .B1(i_data_bus[57]), .B2(n92), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n69), .B1(i_data_bus[56]), .B2(n92), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n69), .B1(i_data_bus[55]), .B2(n92), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n69), .B1(i_data_bus[54]), .B2(n92), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n69), .B1(i_data_bus[53]), .B2(n92), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U140 ( .A1(n70), .A2(n69), .B1(i_data_bus[52]), .B2(n92), 
        .ZN(N339) );
  INVD2BWP30P140 U141 ( .I(n84), .ZN(n82) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n82), .B1(i_data_bus[51]), .B2(n92), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n82), .B1(i_data_bus[50]), .B2(n92), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n82), .B1(i_data_bus[49]), .B2(n92), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n82), .B1(i_data_bus[48]), .B2(n92), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n82), .B1(i_data_bus[47]), .B2(n92), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n82), .B1(i_data_bus[46]), .B2(n92), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n82), .B1(i_data_bus[45]), .B2(n92), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n82), .B1(i_data_bus[44]), .B2(n92), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n82), .B1(i_data_bus[43]), .B2(n92), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n82), .B1(i_data_bus[42]), .B2(n92), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n82), .B1(i_data_bus[41]), .B2(n92), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n82), .B1(i_data_bus[40]), .B2(n92), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U154 ( .A1(n85), .A2(n1), .B1(i_data_bus[32]), .B2(n92), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U155 ( .A1(n86), .A2(n1), .B1(i_data_bus[33]), .B2(n92), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U156 ( .A1(n87), .A2(n1), .B1(i_data_bus[34]), .B2(n92), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U157 ( .A1(n88), .A2(n1), .B1(i_data_bus[35]), .B2(n92), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U158 ( .A1(n89), .A2(n1), .B1(i_data_bus[36]), .B2(n92), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U159 ( .A1(n90), .A2(n1), .B1(i_data_bus[37]), .B2(n92), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U160 ( .A1(n91), .A2(n1), .B1(i_data_bus[38]), .B2(n92), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n1), .B1(i_data_bus[39]), .B2(n92), 
        .ZN(N326) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_119 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD1BWP30P140 U3 ( .I(n57), .ZN(n84) );
  INVD2BWP30P140 U4 ( .I(n84), .ZN(n82) );
  NR2D1BWP30P140 U5 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  OAI22D1BWP30P140 U6 ( .A1(n19), .A2(n7), .B1(n47), .B2(n83), .ZN(N295) );
  OAI22D1BWP30P140 U7 ( .A1(n19), .A2(n8), .B1(n47), .B2(n81), .ZN(N296) );
  OAI22D1BWP30P140 U8 ( .A1(n19), .A2(n9), .B1(n47), .B2(n80), .ZN(N297) );
  OAI22D1BWP30P140 U9 ( .A1(n19), .A2(n10), .B1(n47), .B2(n79), .ZN(N298) );
  OAI22D1BWP30P140 U10 ( .A1(n19), .A2(n11), .B1(n47), .B2(n78), .ZN(N299) );
  OAI22D1BWP30P140 U11 ( .A1(n19), .A2(n12), .B1(n47), .B2(n77), .ZN(N300) );
  OAI22D1BWP30P140 U12 ( .A1(n19), .A2(n13), .B1(n47), .B2(n76), .ZN(N301) );
  OAI22D1BWP30P140 U13 ( .A1(n19), .A2(n14), .B1(n47), .B2(n75), .ZN(N302) );
  OAI22D1BWP30P140 U14 ( .A1(n19), .A2(n15), .B1(n47), .B2(n74), .ZN(N303) );
  OAI22D1BWP30P140 U15 ( .A1(n19), .A2(n16), .B1(n47), .B2(n73), .ZN(N304) );
  OAI22D1BWP30P140 U16 ( .A1(n19), .A2(n17), .B1(n47), .B2(n72), .ZN(N305) );
  OAI22D1BWP30P140 U17 ( .A1(n33), .A2(n20), .B1(n31), .B2(n70), .ZN(N307) );
  OAI22D1BWP30P140 U18 ( .A1(n33), .A2(n21), .B1(n31), .B2(n68), .ZN(N308) );
  OAI22D1BWP30P140 U19 ( .A1(n33), .A2(n22), .B1(n31), .B2(n67), .ZN(N309) );
  OAI22D1BWP30P140 U20 ( .A1(n33), .A2(n23), .B1(n31), .B2(n66), .ZN(N310) );
  OAI22D1BWP30P140 U21 ( .A1(n33), .A2(n24), .B1(n31), .B2(n65), .ZN(N311) );
  OAI22D1BWP30P140 U22 ( .A1(n33), .A2(n25), .B1(n31), .B2(n64), .ZN(N312) );
  OAI22D1BWP30P140 U23 ( .A1(n33), .A2(n26), .B1(n31), .B2(n63), .ZN(N313) );
  OAI22D1BWP30P140 U24 ( .A1(n33), .A2(n27), .B1(n31), .B2(n62), .ZN(N314) );
  OAI22D1BWP30P140 U25 ( .A1(n33), .A2(n28), .B1(n31), .B2(n61), .ZN(N315) );
  OAI22D1BWP30P140 U26 ( .A1(n33), .A2(n29), .B1(n31), .B2(n60), .ZN(N316) );
  OAI22D1BWP30P140 U27 ( .A1(n33), .A2(n30), .B1(n31), .B2(n59), .ZN(N317) );
  OAI22D1BWP30P140 U28 ( .A1(n33), .A2(n32), .B1(n31), .B2(n58), .ZN(N318) );
  ND2D1BWP30P140 U29 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U30 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U31 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U32 ( .I(n92), .ZN(n50) );
  OAI22D1BWP30P140 U33 ( .A1(n19), .A2(n18), .B1(n31), .B2(n71), .ZN(N306) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n19) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n47) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n83) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n81) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n80) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n79) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n78) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n77) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[14]), .ZN(n76) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[47]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[15]), .ZN(n75) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[48]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n74) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n73) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n72) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n18) );
  INVD2BWP30P140 U70 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n71) );
  INVD2BWP30P140 U72 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n20) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n70) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n21) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n68) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n22) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n67) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n23) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n66) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n65) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n64) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n63) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n62) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n61) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n60) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n30) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n59) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n58) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n41) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n41), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[0]), .ZN(n85) );
  INVD2BWP30P140 U100 ( .I(n36), .ZN(n46) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[32]), .ZN(n37) );
  OAI22D1BWP30P140 U102 ( .A1(n41), .A2(n85), .B1(n46), .B2(n37), .ZN(N287) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[1]), .ZN(n86) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[33]), .ZN(n38) );
  OAI22D1BWP30P140 U105 ( .A1(n41), .A2(n86), .B1(n46), .B2(n38), .ZN(N288) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[2]), .ZN(n87) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[34]), .ZN(n39) );
  OAI22D1BWP30P140 U108 ( .A1(n41), .A2(n87), .B1(n46), .B2(n39), .ZN(N289) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[3]), .ZN(n88) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[35]), .ZN(n40) );
  OAI22D1BWP30P140 U111 ( .A1(n41), .A2(n88), .B1(n46), .B2(n40), .ZN(N290) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[4]), .ZN(n89) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[36]), .ZN(n42) );
  OAI22D1BWP30P140 U114 ( .A1(n47), .A2(n89), .B1(n46), .B2(n42), .ZN(N291) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[5]), .ZN(n90) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[37]), .ZN(n43) );
  OAI22D1BWP30P140 U117 ( .A1(n47), .A2(n90), .B1(n46), .B2(n43), .ZN(N292) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[6]), .ZN(n91) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[38]), .ZN(n44) );
  OAI22D1BWP30P140 U120 ( .A1(n47), .A2(n91), .B1(n46), .B2(n44), .ZN(N293) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[7]), .ZN(n93) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[39]), .ZN(n45) );
  OAI22D1BWP30P140 U123 ( .A1(n47), .A2(n93), .B1(n46), .B2(n45), .ZN(N294) );
  INVD1BWP30P140 U124 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U125 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n92) );
  OAI21D1BWP30P140 U127 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  MUX2NUD1BWP30P140 U128 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  INVD2BWP30P140 U129 ( .I(n84), .ZN(n69) );
  MOAI22D1BWP30P140 U130 ( .A1(n58), .A2(n69), .B1(i_data_bus[63]), .B2(n92), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U131 ( .A1(n59), .A2(n69), .B1(i_data_bus[62]), .B2(n92), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U132 ( .A1(n60), .A2(n69), .B1(i_data_bus[61]), .B2(n92), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U133 ( .A1(n61), .A2(n69), .B1(i_data_bus[60]), .B2(n92), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U134 ( .A1(n62), .A2(n69), .B1(i_data_bus[59]), .B2(n92), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U135 ( .A1(n63), .A2(n69), .B1(i_data_bus[58]), .B2(n92), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U136 ( .A1(n64), .A2(n69), .B1(i_data_bus[57]), .B2(n92), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U137 ( .A1(n65), .A2(n69), .B1(i_data_bus[56]), .B2(n92), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U138 ( .A1(n66), .A2(n69), .B1(i_data_bus[55]), .B2(n92), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U139 ( .A1(n67), .A2(n69), .B1(i_data_bus[54]), .B2(n92), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U140 ( .A1(n68), .A2(n69), .B1(i_data_bus[53]), .B2(n92), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n69), .B1(i_data_bus[52]), .B2(n92), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n82), .B1(i_data_bus[51]), .B2(n92), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n82), .B1(i_data_bus[50]), .B2(n92), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n82), .B1(i_data_bus[49]), .B2(n92), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n82), .B1(i_data_bus[48]), .B2(n92), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n82), .B1(i_data_bus[47]), .B2(n92), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n82), .B1(i_data_bus[46]), .B2(n92), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n82), .B1(i_data_bus[45]), .B2(n92), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n82), .B1(i_data_bus[44]), .B2(n92), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n82), .B1(i_data_bus[43]), .B2(n92), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n82), .B1(i_data_bus[42]), .B2(n92), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n82), .B1(i_data_bus[41]), .B2(n92), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n82), .B1(i_data_bus[40]), .B2(n92), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U154 ( .A1(n85), .A2(n1), .B1(i_data_bus[32]), .B2(n92), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U155 ( .A1(n86), .A2(n1), .B1(i_data_bus[33]), .B2(n92), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U156 ( .A1(n87), .A2(n1), .B1(i_data_bus[34]), .B2(n92), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U157 ( .A1(n88), .A2(n1), .B1(i_data_bus[35]), .B2(n92), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U158 ( .A1(n89), .A2(n1), .B1(i_data_bus[36]), .B2(n92), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U159 ( .A1(n90), .A2(n1), .B1(i_data_bus[37]), .B2(n92), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U160 ( .A1(n91), .A2(n1), .B1(i_data_bus[38]), .B2(n92), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n1), .B1(i_data_bus[39]), .B2(n92), 
        .ZN(N326) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_120 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n33), .A2(n32), .B1(n31), .B2(n63), .ZN(N306) );
  INVD2BWP30P140 U4 ( .I(n36), .ZN(n46) );
  OAI22D1BWP30P140 U5 ( .A1(n41), .A2(n88), .B1(n46), .B2(n40), .ZN(N290) );
  INVD1BWP30P140 U6 ( .I(n57), .ZN(n84) );
  ND2D1BWP30P140 U7 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U9 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U10 ( .I(n92), .ZN(n50) );
  OAI22D1BWP30P140 U11 ( .A1(n33), .A2(n10), .B1(n47), .B2(n66), .ZN(N295) );
  OAI22D1BWP30P140 U12 ( .A1(n33), .A2(n11), .B1(n47), .B2(n67), .ZN(N296) );
  OAI22D1BWP30P140 U13 ( .A1(n33), .A2(n12), .B1(n47), .B2(n68), .ZN(N297) );
  OAI22D1BWP30P140 U14 ( .A1(n33), .A2(n13), .B1(n47), .B2(n69), .ZN(N298) );
  OAI22D1BWP30P140 U15 ( .A1(n33), .A2(n15), .B1(n47), .B2(n70), .ZN(N299) );
  OAI22D1BWP30P140 U16 ( .A1(n33), .A2(n17), .B1(n47), .B2(n71), .ZN(N300) );
  OAI22D1BWP30P140 U17 ( .A1(n33), .A2(n9), .B1(n47), .B2(n72), .ZN(N301) );
  OAI22D1BWP30P140 U18 ( .A1(n33), .A2(n8), .B1(n47), .B2(n73), .ZN(N302) );
  OAI22D1BWP30P140 U19 ( .A1(n33), .A2(n16), .B1(n47), .B2(n75), .ZN(N303) );
  OAI22D1BWP30P140 U20 ( .A1(n33), .A2(n14), .B1(n47), .B2(n65), .ZN(N304) );
  OAI22D1BWP30P140 U21 ( .A1(n33), .A2(n7), .B1(n47), .B2(n64), .ZN(N305) );
  OAI22D1BWP30P140 U22 ( .A1(n30), .A2(n29), .B1(n31), .B2(n62), .ZN(N307) );
  OAI22D1BWP30P140 U23 ( .A1(n30), .A2(n28), .B1(n31), .B2(n61), .ZN(N308) );
  OAI22D1BWP30P140 U24 ( .A1(n30), .A2(n27), .B1(n31), .B2(n60), .ZN(N309) );
  OAI22D1BWP30P140 U25 ( .A1(n30), .A2(n26), .B1(n31), .B2(n59), .ZN(N310) );
  OAI22D1BWP30P140 U26 ( .A1(n30), .A2(n25), .B1(n31), .B2(n58), .ZN(N311) );
  OAI22D1BWP30P140 U27 ( .A1(n30), .A2(n24), .B1(n31), .B2(n83), .ZN(N312) );
  OAI22D1BWP30P140 U28 ( .A1(n30), .A2(n23), .B1(n31), .B2(n81), .ZN(N313) );
  OAI22D1BWP30P140 U29 ( .A1(n30), .A2(n22), .B1(n31), .B2(n80), .ZN(N314) );
  OAI22D1BWP30P140 U30 ( .A1(n30), .A2(n21), .B1(n31), .B2(n79), .ZN(N315) );
  OAI22D1BWP30P140 U31 ( .A1(n30), .A2(n18), .B1(n31), .B2(n78), .ZN(N316) );
  OAI22D1BWP30P140 U32 ( .A1(n30), .A2(n19), .B1(n31), .B2(n77), .ZN(N317) );
  OAI22D1BWP30P140 U33 ( .A1(n30), .A2(n20), .B1(n31), .B2(n76), .ZN(N318) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[50]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n47) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[18]), .ZN(n64) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[47]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[15]), .ZN(n73) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[46]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[14]), .ZN(n72) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[40]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[41]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[9]), .ZN(n67) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[42]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[10]), .ZN(n68) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[43]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[49]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[17]), .ZN(n65) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[44]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[12]), .ZN(n70) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[48]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[16]), .ZN(n75) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[45]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[13]), .ZN(n71) );
  INVD2BWP30P140 U69 ( .I(n36), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[61]), .ZN(n18) );
  INVD2BWP30P140 U71 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[29]), .ZN(n78) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[62]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[30]), .ZN(n77) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[63]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[31]), .ZN(n76) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[60]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[28]), .ZN(n79) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[59]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[27]), .ZN(n80) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[58]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[26]), .ZN(n81) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n83) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[56]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[24]), .ZN(n58) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[55]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[23]), .ZN(n59) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[54]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[22]), .ZN(n60) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[53]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[21]), .ZN(n61) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[52]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[20]), .ZN(n62) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[51]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[19]), .ZN(n63) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n41) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n41), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[1]), .ZN(n86) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[33]), .ZN(n37) );
  OAI22D1BWP30P140 U101 ( .A1(n41), .A2(n86), .B1(n46), .B2(n37), .ZN(N288) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[0]), .ZN(n85) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[32]), .ZN(n38) );
  OAI22D1BWP30P140 U104 ( .A1(n41), .A2(n85), .B1(n46), .B2(n38), .ZN(N287) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[2]), .ZN(n87) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[34]), .ZN(n39) );
  OAI22D1BWP30P140 U107 ( .A1(n41), .A2(n87), .B1(n46), .B2(n39), .ZN(N289) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[3]), .ZN(n88) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[35]), .ZN(n40) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[4]), .ZN(n89) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[36]), .ZN(n42) );
  OAI22D1BWP30P140 U112 ( .A1(n47), .A2(n89), .B1(n46), .B2(n42), .ZN(N291) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[5]), .ZN(n90) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[37]), .ZN(n43) );
  OAI22D1BWP30P140 U115 ( .A1(n47), .A2(n90), .B1(n46), .B2(n43), .ZN(N292) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[6]), .ZN(n91) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[38]), .ZN(n44) );
  OAI22D1BWP30P140 U118 ( .A1(n47), .A2(n91), .B1(n46), .B2(n44), .ZN(N293) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[7]), .ZN(n93) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[39]), .ZN(n45) );
  OAI22D1BWP30P140 U121 ( .A1(n47), .A2(n93), .B1(n46), .B2(n45), .ZN(N294) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n92) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  INVD2BWP30P140 U128 ( .I(n84), .ZN(n82) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n82), .B1(i_data_bus[56]), .B2(n92), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n82), .B1(i_data_bus[55]), .B2(n92), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n82), .B1(i_data_bus[54]), .B2(n92), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n82), .B1(i_data_bus[53]), .B2(n92), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n82), .B1(i_data_bus[52]), .B2(n92), 
        .ZN(N339) );
  INVD2BWP30P140 U134 ( .I(n84), .ZN(n74) );
  MOAI22D1BWP30P140 U135 ( .A1(n63), .A2(n74), .B1(i_data_bus[51]), .B2(n92), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U136 ( .A1(n64), .A2(n74), .B1(i_data_bus[50]), .B2(n92), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U137 ( .A1(n65), .A2(n74), .B1(i_data_bus[49]), .B2(n92), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U138 ( .A1(n66), .A2(n74), .B1(i_data_bus[40]), .B2(n92), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U139 ( .A1(n67), .A2(n74), .B1(i_data_bus[41]), .B2(n92), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U140 ( .A1(n68), .A2(n74), .B1(i_data_bus[42]), .B2(n92), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U141 ( .A1(n69), .A2(n74), .B1(i_data_bus[43]), .B2(n92), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U142 ( .A1(n70), .A2(n74), .B1(i_data_bus[44]), .B2(n92), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U143 ( .A1(n71), .A2(n74), .B1(i_data_bus[45]), .B2(n92), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U144 ( .A1(n72), .A2(n74), .B1(i_data_bus[46]), .B2(n92), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U145 ( .A1(n73), .A2(n74), .B1(i_data_bus[47]), .B2(n92), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n74), .B1(i_data_bus[48]), .B2(n92), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n82), .B1(i_data_bus[63]), .B2(n92), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U148 ( .A1(n77), .A2(n82), .B1(i_data_bus[62]), .B2(n92), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n82), .B1(i_data_bus[61]), .B2(n92), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n82), .B1(i_data_bus[60]), .B2(n92), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n82), .B1(i_data_bus[59]), .B2(n92), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n82), .B1(i_data_bus[58]), .B2(n92), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n82), .B1(i_data_bus[57]), .B2(n92), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U154 ( .A1(n85), .A2(n1), .B1(i_data_bus[32]), .B2(n92), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U155 ( .A1(n86), .A2(n1), .B1(i_data_bus[33]), .B2(n92), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U156 ( .A1(n87), .A2(n1), .B1(i_data_bus[34]), .B2(n92), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U157 ( .A1(n88), .A2(n1), .B1(i_data_bus[35]), .B2(n92), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U158 ( .A1(n89), .A2(n1), .B1(i_data_bus[36]), .B2(n92), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U159 ( .A1(n90), .A2(n1), .B1(i_data_bus[37]), .B2(n92), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U160 ( .A1(n91), .A2(n1), .B1(i_data_bus[38]), .B2(n92), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n1), .B1(i_data_bus[39]), .B2(n92), 
        .ZN(N326) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_121 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD1BWP30P140 U3 ( .I(i_cmd[0]), .ZN(n35) );
  OAI22D1BWP30P140 U4 ( .A1(n19), .A2(n15), .B1(n47), .B2(n66), .ZN(N295) );
  INVD2BWP30P140 U5 ( .I(n36), .ZN(n46) );
  OAI22D1BWP30P140 U6 ( .A1(n44), .A2(n62), .B1(n46), .B2(n43), .ZN(N290) );
  OAI22D1BWP30P140 U7 ( .A1(n33), .A2(n20), .B1(n31), .B2(n80), .ZN(N307) );
  OAI22D1BWP30P140 U8 ( .A1(n33), .A2(n21), .B1(n31), .B2(n81), .ZN(N308) );
  OAI22D1BWP30P140 U9 ( .A1(n33), .A2(n32), .B1(n31), .B2(n82), .ZN(N309) );
  OAI22D1BWP30P140 U10 ( .A1(n33), .A2(n22), .B1(n31), .B2(n83), .ZN(N310) );
  OAI22D1BWP30P140 U11 ( .A1(n33), .A2(n28), .B1(n31), .B2(n84), .ZN(N311) );
  OAI22D1BWP30P140 U12 ( .A1(n33), .A2(n23), .B1(n31), .B2(n85), .ZN(N312) );
  OAI22D1BWP30P140 U13 ( .A1(n33), .A2(n27), .B1(n31), .B2(n86), .ZN(N313) );
  OAI22D1BWP30P140 U14 ( .A1(n33), .A2(n30), .B1(n31), .B2(n87), .ZN(N314) );
  OAI22D1BWP30P140 U15 ( .A1(n33), .A2(n24), .B1(n31), .B2(n88), .ZN(N315) );
  OAI22D1BWP30P140 U16 ( .A1(n33), .A2(n26), .B1(n31), .B2(n89), .ZN(N316) );
  OAI22D1BWP30P140 U17 ( .A1(n33), .A2(n25), .B1(n31), .B2(n90), .ZN(N317) );
  OAI22D1BWP30P140 U18 ( .A1(n33), .A2(n29), .B1(n31), .B2(n93), .ZN(N318) );
  INVD1BWP30P140 U19 ( .I(n57), .ZN(n79) );
  ND2D1BWP30P140 U20 ( .A1(n2), .A2(i_en), .ZN(n52) );
  CKBD1BWP30P140 U21 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U22 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U23 ( .A1(n19), .A2(n14), .B1(n47), .B2(n67), .ZN(N296) );
  OAI22D1BWP30P140 U24 ( .A1(n19), .A2(n13), .B1(n47), .B2(n68), .ZN(N297) );
  OAI22D1BWP30P140 U25 ( .A1(n19), .A2(n12), .B1(n47), .B2(n69), .ZN(N298) );
  OAI22D1BWP30P140 U26 ( .A1(n19), .A2(n17), .B1(n47), .B2(n70), .ZN(N299) );
  OAI22D1BWP30P140 U27 ( .A1(n19), .A2(n16), .B1(n47), .B2(n71), .ZN(N300) );
  OAI22D1BWP30P140 U28 ( .A1(n19), .A2(n11), .B1(n47), .B2(n72), .ZN(N301) );
  OAI22D1BWP30P140 U29 ( .A1(n19), .A2(n10), .B1(n47), .B2(n73), .ZN(N302) );
  OAI22D1BWP30P140 U30 ( .A1(n19), .A2(n9), .B1(n47), .B2(n74), .ZN(N303) );
  OAI22D1BWP30P140 U31 ( .A1(n19), .A2(n8), .B1(n47), .B2(n75), .ZN(N304) );
  OAI22D1BWP30P140 U32 ( .A1(n19), .A2(n7), .B1(n47), .B2(n76), .ZN(N305) );
  OAI22D1BWP30P140 U33 ( .A1(n19), .A2(n18), .B1(n31), .B2(n78), .ZN(N306) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n19) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[50]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n47) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[18]), .ZN(n76) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[49]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[17]), .ZN(n75) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[48]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[16]), .ZN(n74) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[47]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[15]), .ZN(n73) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[46]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[14]), .ZN(n72) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[43]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[42]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[10]), .ZN(n68) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[41]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[9]), .ZN(n67) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[40]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[45]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[13]), .ZN(n71) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[44]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[12]), .ZN(n70) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n18) );
  INVD2BWP30P140 U70 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD2BWP30P140 U72 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n20) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n21) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n81) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[55]), .ZN(n22) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[23]), .ZN(n83) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[57]), .ZN(n23) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[25]), .ZN(n85) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[60]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[28]), .ZN(n88) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[62]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[30]), .ZN(n90) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[61]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[29]), .ZN(n89) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[58]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[26]), .ZN(n86) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[56]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[24]), .ZN(n84) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[63]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[31]), .ZN(n93) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[59]), .ZN(n30) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[27]), .ZN(n87) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[54]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[22]), .ZN(n82) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n44) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n44), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[2]), .ZN(n63) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[34]), .ZN(n37) );
  OAI22D1BWP30P140 U101 ( .A1(n44), .A2(n63), .B1(n46), .B2(n37), .ZN(N289) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[0]), .ZN(n65) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[32]), .ZN(n38) );
  OAI22D1BWP30P140 U104 ( .A1(n44), .A2(n65), .B1(n46), .B2(n38), .ZN(N287) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U107 ( .A1(n47), .A2(n61), .B1(n46), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[1]), .ZN(n64) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[33]), .ZN(n40) );
  OAI22D1BWP30P140 U110 ( .A1(n44), .A2(n64), .B1(n46), .B2(n40), .ZN(N288) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[7]), .ZN(n58) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[39]), .ZN(n41) );
  OAI22D1BWP30P140 U113 ( .A1(n47), .A2(n58), .B1(n46), .B2(n41), .ZN(N294) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[5]), .ZN(n60) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[37]), .ZN(n42) );
  OAI22D1BWP30P140 U116 ( .A1(n47), .A2(n60), .B1(n46), .B2(n42), .ZN(N292) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[3]), .ZN(n62) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[35]), .ZN(n43) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[6]), .ZN(n59) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[38]), .ZN(n45) );
  OAI22D1BWP30P140 U121 ( .A1(n47), .A2(n59), .B1(n46), .B2(n45), .ZN(N293) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  INVD2BWP30P140 U136 ( .I(n79), .ZN(n77) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n77), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n77), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n77), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n77), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n77), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n77), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n77), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n77), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n77), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n77), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n77), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n77), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  INVD2BWP30P140 U149 ( .I(n79), .ZN(n92) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n92), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_122 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n19), .A2(n18), .B1(n31), .B2(n78), .ZN(N306) );
  INVD2BWP30P140 U4 ( .I(n36), .ZN(n46) );
  OAI22D1BWP30P140 U5 ( .A1(n47), .A2(n65), .B1(n46), .B2(n45), .ZN(N287) );
  INVD1BWP30P140 U6 ( .I(n57), .ZN(n79) );
  ND2D1BWP30P140 U7 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U9 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U10 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U11 ( .A1(n19), .A2(n7), .B1(n41), .B2(n66), .ZN(N295) );
  OAI22D1BWP30P140 U12 ( .A1(n19), .A2(n8), .B1(n41), .B2(n67), .ZN(N296) );
  OAI22D1BWP30P140 U13 ( .A1(n19), .A2(n9), .B1(n41), .B2(n68), .ZN(N297) );
  OAI22D1BWP30P140 U14 ( .A1(n19), .A2(n10), .B1(n41), .B2(n69), .ZN(N298) );
  OAI22D1BWP30P140 U15 ( .A1(n19), .A2(n11), .B1(n41), .B2(n70), .ZN(N299) );
  OAI22D1BWP30P140 U16 ( .A1(n19), .A2(n12), .B1(n41), .B2(n71), .ZN(N300) );
  OAI22D1BWP30P140 U17 ( .A1(n19), .A2(n13), .B1(n41), .B2(n72), .ZN(N301) );
  OAI22D1BWP30P140 U18 ( .A1(n19), .A2(n14), .B1(n41), .B2(n73), .ZN(N302) );
  OAI22D1BWP30P140 U19 ( .A1(n19), .A2(n15), .B1(n41), .B2(n74), .ZN(N303) );
  OAI22D1BWP30P140 U20 ( .A1(n19), .A2(n16), .B1(n41), .B2(n75), .ZN(N304) );
  OAI22D1BWP30P140 U21 ( .A1(n19), .A2(n17), .B1(n41), .B2(n76), .ZN(N305) );
  OAI22D1BWP30P140 U22 ( .A1(n33), .A2(n20), .B1(n31), .B2(n80), .ZN(N307) );
  OAI22D1BWP30P140 U23 ( .A1(n33), .A2(n21), .B1(n31), .B2(n81), .ZN(N308) );
  OAI22D1BWP30P140 U24 ( .A1(n33), .A2(n22), .B1(n31), .B2(n82), .ZN(N309) );
  OAI22D1BWP30P140 U25 ( .A1(n33), .A2(n23), .B1(n31), .B2(n83), .ZN(N310) );
  OAI22D1BWP30P140 U26 ( .A1(n33), .A2(n24), .B1(n31), .B2(n84), .ZN(N311) );
  OAI22D1BWP30P140 U27 ( .A1(n33), .A2(n25), .B1(n31), .B2(n85), .ZN(N312) );
  OAI22D1BWP30P140 U28 ( .A1(n33), .A2(n26), .B1(n31), .B2(n86), .ZN(N313) );
  OAI22D1BWP30P140 U29 ( .A1(n33), .A2(n27), .B1(n31), .B2(n87), .ZN(N314) );
  OAI22D1BWP30P140 U30 ( .A1(n33), .A2(n28), .B1(n31), .B2(n88), .ZN(N315) );
  OAI22D1BWP30P140 U31 ( .A1(n33), .A2(n29), .B1(n31), .B2(n89), .ZN(N316) );
  OAI22D1BWP30P140 U32 ( .A1(n33), .A2(n30), .B1(n31), .B2(n90), .ZN(N317) );
  OAI22D1BWP30P140 U33 ( .A1(n33), .A2(n32), .B1(n31), .B2(n93), .ZN(N318) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n19) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n41) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n67) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n68) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n70) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n71) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[14]), .ZN(n72) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[47]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[15]), .ZN(n73) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[48]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n74) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n75) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n76) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[51]), .ZN(n18) );
  INVD2BWP30P140 U70 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD2BWP30P140 U72 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[52]), .ZN(n20) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[53]), .ZN(n21) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[21]), .ZN(n81) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[54]), .ZN(n22) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[22]), .ZN(n82) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[55]), .ZN(n23) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[23]), .ZN(n83) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[56]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n84) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n85) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[58]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[26]), .ZN(n86) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[59]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[27]), .ZN(n87) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[60]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[28]), .ZN(n88) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[61]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[29]), .ZN(n89) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[62]), .ZN(n30) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[30]), .ZN(n90) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[63]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[31]), .ZN(n93) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n47) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n47), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n58) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[39]), .ZN(n37) );
  OAI22D1BWP30P140 U101 ( .A1(n41), .A2(n58), .B1(n46), .B2(n37), .ZN(N294) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[6]), .ZN(n59) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[38]), .ZN(n38) );
  OAI22D1BWP30P140 U104 ( .A1(n41), .A2(n59), .B1(n46), .B2(n38), .ZN(N293) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[5]), .ZN(n60) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[37]), .ZN(n39) );
  OAI22D1BWP30P140 U107 ( .A1(n41), .A2(n60), .B1(n46), .B2(n39), .ZN(N292) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[4]), .ZN(n61) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[36]), .ZN(n40) );
  OAI22D1BWP30P140 U110 ( .A1(n41), .A2(n61), .B1(n46), .B2(n40), .ZN(N291) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[3]), .ZN(n62) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[35]), .ZN(n42) );
  OAI22D1BWP30P140 U113 ( .A1(n47), .A2(n62), .B1(n46), .B2(n42), .ZN(N290) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[2]), .ZN(n63) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[34]), .ZN(n43) );
  OAI22D1BWP30P140 U116 ( .A1(n47), .A2(n63), .B1(n46), .B2(n43), .ZN(N289) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[1]), .ZN(n64) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[33]), .ZN(n44) );
  OAI22D1BWP30P140 U119 ( .A1(n47), .A2(n64), .B1(n46), .B2(n44), .ZN(N288) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[0]), .ZN(n65) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[32]), .ZN(n45) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  INVD2BWP30P140 U136 ( .I(n79), .ZN(n77) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n77), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n77), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n77), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n77), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n77), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n77), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n77), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n77), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n77), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n77), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n77), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n77), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  INVD2BWP30P140 U149 ( .I(n79), .ZN(n92) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n92), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_123 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD1BWP30P140 U3 ( .I(n57), .ZN(n77) );
  INVD2BWP30P140 U4 ( .I(n77), .ZN(n89) );
  NR2D1BWP30P140 U5 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  OAI22D1BWP30P140 U6 ( .A1(n23), .A2(n14), .B1(n41), .B2(n93), .ZN(N295) );
  OAI22D1BWP30P140 U7 ( .A1(n23), .A2(n17), .B1(n41), .B2(n66), .ZN(N296) );
  OAI22D1BWP30P140 U8 ( .A1(n23), .A2(n13), .B1(n41), .B2(n67), .ZN(N297) );
  OAI22D1BWP30P140 U9 ( .A1(n23), .A2(n16), .B1(n41), .B2(n68), .ZN(N298) );
  OAI22D1BWP30P140 U10 ( .A1(n23), .A2(n8), .B1(n41), .B2(n69), .ZN(N299) );
  OAI22D1BWP30P140 U11 ( .A1(n23), .A2(n12), .B1(n41), .B2(n70), .ZN(N300) );
  OAI22D1BWP30P140 U12 ( .A1(n23), .A2(n11), .B1(n41), .B2(n71), .ZN(N301) );
  OAI22D1BWP30P140 U13 ( .A1(n23), .A2(n7), .B1(n41), .B2(n72), .ZN(N302) );
  OAI22D1BWP30P140 U14 ( .A1(n23), .A2(n10), .B1(n41), .B2(n73), .ZN(N303) );
  OAI22D1BWP30P140 U15 ( .A1(n23), .A2(n9), .B1(n41), .B2(n74), .ZN(N304) );
  OAI22D1BWP30P140 U16 ( .A1(n23), .A2(n15), .B1(n41), .B2(n75), .ZN(N305) );
  OAI22D1BWP30P140 U17 ( .A1(n33), .A2(n20), .B1(n31), .B2(n78), .ZN(N307) );
  OAI22D1BWP30P140 U18 ( .A1(n33), .A2(n32), .B1(n31), .B2(n79), .ZN(N308) );
  OAI22D1BWP30P140 U19 ( .A1(n33), .A2(n24), .B1(n31), .B2(n80), .ZN(N309) );
  OAI22D1BWP30P140 U20 ( .A1(n33), .A2(n30), .B1(n31), .B2(n81), .ZN(N310) );
  OAI22D1BWP30P140 U21 ( .A1(n33), .A2(n29), .B1(n31), .B2(n82), .ZN(N311) );
  OAI22D1BWP30P140 U22 ( .A1(n33), .A2(n28), .B1(n31), .B2(n83), .ZN(N312) );
  OAI22D1BWP30P140 U23 ( .A1(n33), .A2(n27), .B1(n31), .B2(n84), .ZN(N313) );
  OAI22D1BWP30P140 U24 ( .A1(n33), .A2(n26), .B1(n31), .B2(n85), .ZN(N314) );
  OAI22D1BWP30P140 U25 ( .A1(n33), .A2(n25), .B1(n31), .B2(n86), .ZN(N315) );
  OAI22D1BWP30P140 U26 ( .A1(n33), .A2(n21), .B1(n31), .B2(n87), .ZN(N316) );
  OAI22D1BWP30P140 U27 ( .A1(n33), .A2(n19), .B1(n31), .B2(n88), .ZN(N317) );
  OAI22D1BWP30P140 U28 ( .A1(n33), .A2(n18), .B1(n31), .B2(n90), .ZN(N318) );
  ND2D1BWP30P140 U29 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U30 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U31 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U32 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U33 ( .A1(n23), .A2(n22), .B1(n31), .B2(n76), .ZN(N306) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n23) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[47]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n41) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[15]), .ZN(n72) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[44]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[12]), .ZN(n69) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[49]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[17]), .ZN(n74) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[48]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[46]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[14]), .ZN(n71) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n70) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[42]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[10]), .ZN(n67) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[40]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[8]), .ZN(n93) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[50]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[18]), .ZN(n75) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[43]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[11]), .ZN(n68) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[41]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[9]), .ZN(n66) );
  INVD2BWP30P140 U69 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[63]), .ZN(n18) );
  INVD2BWP30P140 U71 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[31]), .ZN(n90) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[62]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[30]), .ZN(n88) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[52]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[20]), .ZN(n78) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[61]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[29]), .ZN(n87) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[51]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[19]), .ZN(n76) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[54]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[22]), .ZN(n80) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[60]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[28]), .ZN(n86) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[59]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[27]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[58]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[26]), .ZN(n84) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[57]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[25]), .ZN(n83) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[56]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[24]), .ZN(n82) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[55]), .ZN(n30) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[23]), .ZN(n81) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[53]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[21]), .ZN(n79) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n47) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n47), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n60) );
  INVD2BWP30P140 U100 ( .I(n36), .ZN(n46) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[39]), .ZN(n37) );
  OAI22D1BWP30P140 U102 ( .A1(n41), .A2(n60), .B1(n46), .B2(n37), .ZN(N294) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[5]), .ZN(n62) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U105 ( .A1(n41), .A2(n62), .B1(n46), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[6]), .ZN(n61) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[38]), .ZN(n39) );
  OAI22D1BWP30P140 U108 ( .A1(n41), .A2(n61), .B1(n46), .B2(n39), .ZN(N293) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[4]), .ZN(n63) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[36]), .ZN(n40) );
  OAI22D1BWP30P140 U111 ( .A1(n41), .A2(n63), .B1(n46), .B2(n40), .ZN(N291) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[3]), .ZN(n64) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[35]), .ZN(n42) );
  OAI22D1BWP30P140 U114 ( .A1(n47), .A2(n64), .B1(n46), .B2(n42), .ZN(N290) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[2]), .ZN(n65) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[34]), .ZN(n43) );
  OAI22D1BWP30P140 U117 ( .A1(n47), .A2(n65), .B1(n46), .B2(n43), .ZN(N289) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[1]), .ZN(n58) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[33]), .ZN(n44) );
  OAI22D1BWP30P140 U120 ( .A1(n47), .A2(n58), .B1(n46), .B2(n44), .ZN(N288) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[0]), .ZN(n59) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[32]), .ZN(n45) );
  OAI22D1BWP30P140 U123 ( .A1(n47), .A2(n59), .B1(n46), .B2(n45), .ZN(N287) );
  INVD1BWP30P140 U124 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U125 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U127 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  MUX2NUD1BWP30P140 U128 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  INVD2BWP30P140 U137 ( .I(n77), .ZN(n92) );
  MOAI22D1BWP30P140 U138 ( .A1(n66), .A2(n92), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U139 ( .A1(n67), .A2(n92), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U140 ( .A1(n68), .A2(n92), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U141 ( .A1(n69), .A2(n92), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U142 ( .A1(n70), .A2(n92), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U143 ( .A1(n71), .A2(n92), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U144 ( .A1(n72), .A2(n92), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U145 ( .A1(n73), .A2(n92), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U146 ( .A1(n74), .A2(n92), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U147 ( .A1(n75), .A2(n92), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U148 ( .A1(n76), .A2(n92), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n89), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U150 ( .A1(n79), .A2(n89), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U151 ( .A1(n80), .A2(n89), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U152 ( .A1(n81), .A2(n89), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U153 ( .A1(n82), .A2(n89), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U154 ( .A1(n83), .A2(n89), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U155 ( .A1(n84), .A2(n89), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U156 ( .A1(n85), .A2(n89), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U157 ( .A1(n86), .A2(n89), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U158 ( .A1(n87), .A2(n89), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U159 ( .A1(n88), .A2(n89), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n89), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_124 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n33), .A2(n32), .B1(n31), .B2(n78), .ZN(N306) );
  INVD2BWP30P140 U4 ( .I(n36), .ZN(n46) );
  OAI22D1BWP30P140 U5 ( .A1(n47), .A2(n58), .B1(n46), .B2(n45), .ZN(N287) );
  INVD1BWP30P140 U6 ( .I(n57), .ZN(n79) );
  ND2D1BWP30P140 U7 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U9 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U10 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U11 ( .A1(n33), .A2(n16), .B1(n44), .B2(n66), .ZN(N295) );
  OAI22D1BWP30P140 U12 ( .A1(n33), .A2(n17), .B1(n44), .B2(n67), .ZN(N296) );
  OAI22D1BWP30P140 U13 ( .A1(n33), .A2(n15), .B1(n44), .B2(n68), .ZN(N297) );
  OAI22D1BWP30P140 U14 ( .A1(n33), .A2(n14), .B1(n44), .B2(n69), .ZN(N298) );
  OAI22D1BWP30P140 U15 ( .A1(n33), .A2(n13), .B1(n44), .B2(n70), .ZN(N299) );
  OAI22D1BWP30P140 U16 ( .A1(n33), .A2(n12), .B1(n44), .B2(n71), .ZN(N300) );
  OAI22D1BWP30P140 U17 ( .A1(n33), .A2(n11), .B1(n44), .B2(n72), .ZN(N301) );
  OAI22D1BWP30P140 U18 ( .A1(n33), .A2(n10), .B1(n44), .B2(n73), .ZN(N302) );
  OAI22D1BWP30P140 U19 ( .A1(n33), .A2(n9), .B1(n44), .B2(n74), .ZN(N303) );
  OAI22D1BWP30P140 U20 ( .A1(n33), .A2(n8), .B1(n44), .B2(n75), .ZN(N304) );
  OAI22D1BWP30P140 U21 ( .A1(n33), .A2(n7), .B1(n44), .B2(n76), .ZN(N305) );
  OAI22D1BWP30P140 U22 ( .A1(n30), .A2(n29), .B1(n31), .B2(n80), .ZN(N307) );
  OAI22D1BWP30P140 U23 ( .A1(n30), .A2(n28), .B1(n31), .B2(n81), .ZN(N308) );
  OAI22D1BWP30P140 U24 ( .A1(n30), .A2(n27), .B1(n31), .B2(n82), .ZN(N309) );
  OAI22D1BWP30P140 U25 ( .A1(n30), .A2(n26), .B1(n31), .B2(n83), .ZN(N310) );
  OAI22D1BWP30P140 U26 ( .A1(n30), .A2(n25), .B1(n31), .B2(n84), .ZN(N311) );
  OAI22D1BWP30P140 U27 ( .A1(n30), .A2(n24), .B1(n31), .B2(n85), .ZN(N312) );
  OAI22D1BWP30P140 U28 ( .A1(n30), .A2(n23), .B1(n31), .B2(n86), .ZN(N313) );
  OAI22D1BWP30P140 U29 ( .A1(n30), .A2(n22), .B1(n31), .B2(n87), .ZN(N314) );
  OAI22D1BWP30P140 U30 ( .A1(n30), .A2(n21), .B1(n31), .B2(n88), .ZN(N315) );
  OAI22D1BWP30P140 U31 ( .A1(n30), .A2(n20), .B1(n31), .B2(n89), .ZN(N316) );
  OAI22D1BWP30P140 U32 ( .A1(n30), .A2(n19), .B1(n31), .B2(n90), .ZN(N317) );
  OAI22D1BWP30P140 U33 ( .A1(n30), .A2(n18), .B1(n31), .B2(n93), .ZN(N318) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[50]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n44) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[18]), .ZN(n76) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[49]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[17]), .ZN(n75) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[48]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[16]), .ZN(n74) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[47]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[15]), .ZN(n73) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[46]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[14]), .ZN(n72) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n71) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[44]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[12]), .ZN(n70) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[43]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[42]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[10]), .ZN(n68) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[40]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[41]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[9]), .ZN(n67) );
  INVD2BWP30P140 U69 ( .I(n36), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[63]), .ZN(n18) );
  INVD2BWP30P140 U71 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[31]), .ZN(n93) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[62]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[30]), .ZN(n90) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[61]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[29]), .ZN(n89) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[60]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[28]), .ZN(n88) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[59]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[27]), .ZN(n87) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[58]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[26]), .ZN(n86) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n85) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[56]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[24]), .ZN(n84) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[55]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[23]), .ZN(n83) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[54]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[22]), .ZN(n82) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[53]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[21]), .ZN(n81) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[52]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[51]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n47) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n47), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[35]), .ZN(n37) );
  OAI22D1BWP30P140 U101 ( .A1(n47), .A2(n61), .B1(n46), .B2(n37), .ZN(N290) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[34]), .ZN(n38) );
  OAI22D1BWP30P140 U104 ( .A1(n47), .A2(n60), .B1(n46), .B2(n38), .ZN(N289) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[33]), .ZN(n39) );
  OAI22D1BWP30P140 U107 ( .A1(n47), .A2(n59), .B1(n46), .B2(n39), .ZN(N288) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[7]), .ZN(n65) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[39]), .ZN(n40) );
  OAI22D1BWP30P140 U110 ( .A1(n44), .A2(n65), .B1(n46), .B2(n40), .ZN(N294) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[6]), .ZN(n64) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[38]), .ZN(n41) );
  OAI22D1BWP30P140 U113 ( .A1(n44), .A2(n64), .B1(n46), .B2(n41), .ZN(N293) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[5]), .ZN(n63) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[37]), .ZN(n42) );
  OAI22D1BWP30P140 U116 ( .A1(n44), .A2(n63), .B1(n46), .B2(n42), .ZN(N292) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[36]), .ZN(n43) );
  OAI22D1BWP30P140 U119 ( .A1(n44), .A2(n62), .B1(n46), .B2(n43), .ZN(N291) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[0]), .ZN(n58) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[32]), .ZN(n45) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  INVD2BWP30P140 U136 ( .I(n79), .ZN(n77) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n77), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n77), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n77), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n77), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n77), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n77), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n77), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n77), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n77), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n77), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n77), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n77), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  INVD2BWP30P140 U149 ( .I(n79), .ZN(n92) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n92), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_125 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD2BWP30P140 U3 ( .I(n36), .ZN(n46) );
  OAI22D1BWP30P140 U4 ( .A1(n47), .A2(n65), .B1(n46), .B2(n45), .ZN(N294) );
  OAI22D1BWP30P140 U5 ( .A1(n20), .A2(n19), .B1(n31), .B2(n78), .ZN(N306) );
  INVD1BWP30P140 U6 ( .I(n57), .ZN(n79) );
  ND2D1BWP30P140 U7 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U9 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U10 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U11 ( .A1(n20), .A2(n14), .B1(n47), .B2(n66), .ZN(N295) );
  OAI22D1BWP30P140 U12 ( .A1(n20), .A2(n7), .B1(n47), .B2(n67), .ZN(N296) );
  OAI22D1BWP30P140 U13 ( .A1(n20), .A2(n9), .B1(n47), .B2(n68), .ZN(N297) );
  OAI22D1BWP30P140 U14 ( .A1(n20), .A2(n10), .B1(n47), .B2(n69), .ZN(N298) );
  OAI22D1BWP30P140 U15 ( .A1(n20), .A2(n15), .B1(n47), .B2(n70), .ZN(N299) );
  OAI22D1BWP30P140 U16 ( .A1(n20), .A2(n13), .B1(n47), .B2(n71), .ZN(N300) );
  OAI22D1BWP30P140 U17 ( .A1(n20), .A2(n11), .B1(n47), .B2(n72), .ZN(N301) );
  OAI22D1BWP30P140 U18 ( .A1(n20), .A2(n12), .B1(n47), .B2(n73), .ZN(N302) );
  OAI22D1BWP30P140 U19 ( .A1(n20), .A2(n8), .B1(n47), .B2(n74), .ZN(N303) );
  OAI22D1BWP30P140 U20 ( .A1(n20), .A2(n16), .B1(n47), .B2(n75), .ZN(N304) );
  OAI22D1BWP30P140 U21 ( .A1(n20), .A2(n17), .B1(n47), .B2(n76), .ZN(N305) );
  OAI22D1BWP30P140 U22 ( .A1(n33), .A2(n21), .B1(n31), .B2(n80), .ZN(N307) );
  OAI22D1BWP30P140 U23 ( .A1(n33), .A2(n22), .B1(n31), .B2(n81), .ZN(N308) );
  OAI22D1BWP30P140 U24 ( .A1(n33), .A2(n23), .B1(n31), .B2(n82), .ZN(N309) );
  OAI22D1BWP30P140 U25 ( .A1(n33), .A2(n24), .B1(n31), .B2(n83), .ZN(N310) );
  OAI22D1BWP30P140 U26 ( .A1(n33), .A2(n25), .B1(n31), .B2(n84), .ZN(N311) );
  OAI22D1BWP30P140 U27 ( .A1(n33), .A2(n26), .B1(n31), .B2(n85), .ZN(N312) );
  OAI22D1BWP30P140 U28 ( .A1(n33), .A2(n27), .B1(n31), .B2(n86), .ZN(N313) );
  OAI22D1BWP30P140 U29 ( .A1(n33), .A2(n18), .B1(n31), .B2(n87), .ZN(N314) );
  OAI22D1BWP30P140 U30 ( .A1(n33), .A2(n32), .B1(n31), .B2(n88), .ZN(N315) );
  OAI22D1BWP30P140 U31 ( .A1(n33), .A2(n30), .B1(n31), .B2(n89), .ZN(N316) );
  OAI22D1BWP30P140 U32 ( .A1(n33), .A2(n29), .B1(n31), .B2(n90), .ZN(N317) );
  OAI22D1BWP30P140 U33 ( .A1(n33), .A2(n28), .B1(n31), .B2(n93), .ZN(N318) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n20) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[41]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n47) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[9]), .ZN(n67) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[48]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[16]), .ZN(n74) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n68) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[46]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[14]), .ZN(n72) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[47]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[15]), .ZN(n73) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[45]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[13]), .ZN(n71) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[40]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[44]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[12]), .ZN(n70) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n75) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n76) );
  INVD2BWP30P140 U69 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[59]), .ZN(n18) );
  INVD2BWP30P140 U71 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[27]), .ZN(n87) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[51]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[52]), .ZN(n21) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[53]), .ZN(n22) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[21]), .ZN(n81) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[54]), .ZN(n23) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[22]), .ZN(n82) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[55]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[23]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[56]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[24]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[57]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[25]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[58]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[26]), .ZN(n86) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[63]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[31]), .ZN(n93) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[62]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[30]), .ZN(n90) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[61]), .ZN(n30) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[29]), .ZN(n89) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[60]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[28]), .ZN(n88) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n43) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n43), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[33]), .ZN(n37) );
  OAI22D1BWP30P140 U101 ( .A1(n43), .A2(n59), .B1(n46), .B2(n37), .ZN(N288) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[0]), .ZN(n58) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[32]), .ZN(n38) );
  OAI22D1BWP30P140 U104 ( .A1(n43), .A2(n58), .B1(n46), .B2(n38), .ZN(N287) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U107 ( .A1(n47), .A2(n62), .B1(n46), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[6]), .ZN(n64) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[38]), .ZN(n40) );
  OAI22D1BWP30P140 U110 ( .A1(n47), .A2(n64), .B1(n46), .B2(n40), .ZN(N293) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[34]), .ZN(n41) );
  OAI22D1BWP30P140 U113 ( .A1(n43), .A2(n60), .B1(n46), .B2(n41), .ZN(N289) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[35]), .ZN(n42) );
  OAI22D1BWP30P140 U116 ( .A1(n43), .A2(n61), .B1(n46), .B2(n42), .ZN(N290) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[5]), .ZN(n63) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[37]), .ZN(n44) );
  OAI22D1BWP30P140 U119 ( .A1(n47), .A2(n63), .B1(n46), .B2(n44), .ZN(N292) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[7]), .ZN(n65) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[39]), .ZN(n45) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  INVD2BWP30P140 U136 ( .I(n79), .ZN(n77) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n77), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n77), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n77), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n77), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n77), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n77), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n77), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n77), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n77), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n77), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n77), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n77), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  INVD2BWP30P140 U149 ( .I(n79), .ZN(n92) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n92), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_126 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n33), .A2(n32), .B1(n31), .B2(n78), .ZN(N306) );
  INVD2BWP30P140 U4 ( .I(n36), .ZN(n46) );
  OAI22D1BWP30P140 U5 ( .A1(n47), .A2(n58), .B1(n46), .B2(n45), .ZN(N287) );
  INVD1BWP30P140 U6 ( .I(n57), .ZN(n79) );
  ND2D1BWP30P140 U7 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U9 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U10 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U11 ( .A1(n33), .A2(n14), .B1(n41), .B2(n66), .ZN(N295) );
  OAI22D1BWP30P140 U12 ( .A1(n33), .A2(n16), .B1(n41), .B2(n67), .ZN(N296) );
  OAI22D1BWP30P140 U13 ( .A1(n33), .A2(n17), .B1(n41), .B2(n68), .ZN(N297) );
  OAI22D1BWP30P140 U14 ( .A1(n33), .A2(n15), .B1(n41), .B2(n69), .ZN(N298) );
  OAI22D1BWP30P140 U15 ( .A1(n33), .A2(n13), .B1(n41), .B2(n70), .ZN(N299) );
  OAI22D1BWP30P140 U16 ( .A1(n33), .A2(n12), .B1(n41), .B2(n71), .ZN(N300) );
  OAI22D1BWP30P140 U17 ( .A1(n33), .A2(n11), .B1(n41), .B2(n72), .ZN(N301) );
  OAI22D1BWP30P140 U18 ( .A1(n33), .A2(n10), .B1(n41), .B2(n73), .ZN(N302) );
  OAI22D1BWP30P140 U19 ( .A1(n33), .A2(n9), .B1(n41), .B2(n74), .ZN(N303) );
  OAI22D1BWP30P140 U20 ( .A1(n33), .A2(n8), .B1(n41), .B2(n75), .ZN(N304) );
  OAI22D1BWP30P140 U21 ( .A1(n33), .A2(n7), .B1(n41), .B2(n76), .ZN(N305) );
  OAI22D1BWP30P140 U22 ( .A1(n30), .A2(n29), .B1(n31), .B2(n80), .ZN(N307) );
  OAI22D1BWP30P140 U23 ( .A1(n30), .A2(n28), .B1(n31), .B2(n81), .ZN(N308) );
  OAI22D1BWP30P140 U24 ( .A1(n30), .A2(n27), .B1(n31), .B2(n82), .ZN(N309) );
  OAI22D1BWP30P140 U25 ( .A1(n30), .A2(n26), .B1(n31), .B2(n83), .ZN(N310) );
  OAI22D1BWP30P140 U26 ( .A1(n30), .A2(n25), .B1(n31), .B2(n84), .ZN(N311) );
  OAI22D1BWP30P140 U27 ( .A1(n30), .A2(n24), .B1(n31), .B2(n85), .ZN(N312) );
  OAI22D1BWP30P140 U28 ( .A1(n30), .A2(n23), .B1(n31), .B2(n86), .ZN(N313) );
  OAI22D1BWP30P140 U29 ( .A1(n30), .A2(n22), .B1(n31), .B2(n87), .ZN(N314) );
  OAI22D1BWP30P140 U30 ( .A1(n30), .A2(n21), .B1(n31), .B2(n88), .ZN(N315) );
  OAI22D1BWP30P140 U31 ( .A1(n30), .A2(n20), .B1(n31), .B2(n89), .ZN(N316) );
  OAI22D1BWP30P140 U32 ( .A1(n30), .A2(n19), .B1(n31), .B2(n90), .ZN(N317) );
  OAI22D1BWP30P140 U33 ( .A1(n30), .A2(n18), .B1(n31), .B2(n93), .ZN(N318) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[50]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n41) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[18]), .ZN(n76) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[49]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[17]), .ZN(n75) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[48]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[16]), .ZN(n74) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[47]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[15]), .ZN(n73) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[46]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[14]), .ZN(n72) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n71) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[44]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[12]), .ZN(n70) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[40]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[43]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[41]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[9]), .ZN(n67) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[42]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[10]), .ZN(n68) );
  INVD2BWP30P140 U69 ( .I(n36), .ZN(n30) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[63]), .ZN(n18) );
  INVD2BWP30P140 U71 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[31]), .ZN(n93) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[62]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[30]), .ZN(n90) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[61]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[29]), .ZN(n89) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[60]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[28]), .ZN(n88) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[59]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[27]), .ZN(n87) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[58]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[26]), .ZN(n86) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[57]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[25]), .ZN(n85) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[56]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[24]), .ZN(n84) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[55]), .ZN(n26) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[23]), .ZN(n83) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[54]), .ZN(n27) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[22]), .ZN(n82) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[53]), .ZN(n28) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[21]), .ZN(n81) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[52]), .ZN(n29) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[51]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n47) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n47), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n65) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[39]), .ZN(n37) );
  OAI22D1BWP30P140 U101 ( .A1(n41), .A2(n65), .B1(n46), .B2(n37), .ZN(N294) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[6]), .ZN(n64) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[38]), .ZN(n38) );
  OAI22D1BWP30P140 U104 ( .A1(n41), .A2(n64), .B1(n46), .B2(n38), .ZN(N293) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[5]), .ZN(n63) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[37]), .ZN(n39) );
  OAI22D1BWP30P140 U107 ( .A1(n41), .A2(n63), .B1(n46), .B2(n39), .ZN(N292) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[4]), .ZN(n62) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[36]), .ZN(n40) );
  OAI22D1BWP30P140 U110 ( .A1(n41), .A2(n62), .B1(n46), .B2(n40), .ZN(N291) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[3]), .ZN(n61) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[35]), .ZN(n42) );
  OAI22D1BWP30P140 U113 ( .A1(n47), .A2(n61), .B1(n46), .B2(n42), .ZN(N290) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[2]), .ZN(n60) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[34]), .ZN(n43) );
  OAI22D1BWP30P140 U116 ( .A1(n47), .A2(n60), .B1(n46), .B2(n43), .ZN(N289) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[1]), .ZN(n59) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[33]), .ZN(n44) );
  OAI22D1BWP30P140 U119 ( .A1(n47), .A2(n59), .B1(n46), .B2(n44), .ZN(N288) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[0]), .ZN(n58) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[32]), .ZN(n45) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  INVD2BWP30P140 U136 ( .I(n79), .ZN(n77) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n77), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n77), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n77), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n77), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n77), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n77), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n77), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n77), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n77), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n77), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n77), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n77), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  INVD2BWP30P140 U149 ( .I(n79), .ZN(n92) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n92), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_127 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  INVD1BWP30P140 U3 ( .I(n57), .ZN(n79) );
  INVD2BWP30P140 U4 ( .I(n79), .ZN(n92) );
  NR2D1BWP30P140 U5 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  OAI22D1BWP30P140 U6 ( .A1(n26), .A2(n7), .B1(n47), .B2(n66), .ZN(N295) );
  OAI22D1BWP30P140 U7 ( .A1(n26), .A2(n8), .B1(n47), .B2(n67), .ZN(N296) );
  OAI22D1BWP30P140 U8 ( .A1(n26), .A2(n9), .B1(n47), .B2(n68), .ZN(N297) );
  OAI22D1BWP30P140 U9 ( .A1(n26), .A2(n10), .B1(n47), .B2(n69), .ZN(N298) );
  OAI22D1BWP30P140 U10 ( .A1(n26), .A2(n11), .B1(n47), .B2(n70), .ZN(N299) );
  OAI22D1BWP30P140 U11 ( .A1(n26), .A2(n12), .B1(n47), .B2(n71), .ZN(N300) );
  OAI22D1BWP30P140 U12 ( .A1(n26), .A2(n13), .B1(n47), .B2(n72), .ZN(N301) );
  OAI22D1BWP30P140 U13 ( .A1(n26), .A2(n14), .B1(n47), .B2(n73), .ZN(N302) );
  OAI22D1BWP30P140 U14 ( .A1(n26), .A2(n15), .B1(n47), .B2(n74), .ZN(N303) );
  OAI22D1BWP30P140 U15 ( .A1(n26), .A2(n16), .B1(n47), .B2(n75), .ZN(N304) );
  OAI22D1BWP30P140 U16 ( .A1(n26), .A2(n17), .B1(n47), .B2(n76), .ZN(N305) );
  OAI22D1BWP30P140 U17 ( .A1(n33), .A2(n27), .B1(n31), .B2(n80), .ZN(N307) );
  OAI22D1BWP30P140 U18 ( .A1(n33), .A2(n28), .B1(n31), .B2(n81), .ZN(N308) );
  OAI22D1BWP30P140 U19 ( .A1(n33), .A2(n29), .B1(n31), .B2(n82), .ZN(N309) );
  OAI22D1BWP30P140 U20 ( .A1(n33), .A2(n30), .B1(n31), .B2(n83), .ZN(N310) );
  OAI22D1BWP30P140 U21 ( .A1(n33), .A2(n32), .B1(n31), .B2(n84), .ZN(N311) );
  OAI22D1BWP30P140 U22 ( .A1(n33), .A2(n18), .B1(n31), .B2(n85), .ZN(N312) );
  OAI22D1BWP30P140 U23 ( .A1(n33), .A2(n24), .B1(n31), .B2(n86), .ZN(N313) );
  OAI22D1BWP30P140 U24 ( .A1(n33), .A2(n23), .B1(n31), .B2(n87), .ZN(N314) );
  OAI22D1BWP30P140 U25 ( .A1(n33), .A2(n22), .B1(n31), .B2(n88), .ZN(N315) );
  OAI22D1BWP30P140 U26 ( .A1(n33), .A2(n21), .B1(n31), .B2(n89), .ZN(N316) );
  OAI22D1BWP30P140 U27 ( .A1(n33), .A2(n20), .B1(n31), .B2(n90), .ZN(N317) );
  OAI22D1BWP30P140 U28 ( .A1(n33), .A2(n19), .B1(n31), .B2(n93), .ZN(N318) );
  ND2D1BWP30P140 U29 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U30 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U31 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U32 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U33 ( .A1(n26), .A2(n25), .B1(n31), .B2(n78), .ZN(N306) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n26) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n47) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n67) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n68) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n70) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n71) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[46]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[14]), .ZN(n72) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[47]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[15]), .ZN(n73) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[48]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[16]), .ZN(n74) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[49]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[17]), .ZN(n75) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[50]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[18]), .ZN(n76) );
  INVD2BWP30P140 U69 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[57]), .ZN(n18) );
  INVD2BWP30P140 U71 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[25]), .ZN(n85) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[63]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[31]), .ZN(n93) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[62]), .ZN(n20) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[30]), .ZN(n90) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[61]), .ZN(n21) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[29]), .ZN(n89) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[60]), .ZN(n22) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[28]), .ZN(n88) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[59]), .ZN(n23) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[27]), .ZN(n87) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[58]), .ZN(n24) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[26]), .ZN(n86) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[51]), .ZN(n25) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[52]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[53]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[21]), .ZN(n81) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[54]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[22]), .ZN(n82) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[55]), .ZN(n30) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[23]), .ZN(n83) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[56]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[24]), .ZN(n84) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n43) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n43), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[3]), .ZN(n59) );
  INVD2BWP30P140 U100 ( .I(n36), .ZN(n46) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[35]), .ZN(n37) );
  OAI22D1BWP30P140 U102 ( .A1(n43), .A2(n59), .B1(n46), .B2(n37), .ZN(N290) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[2]), .ZN(n58) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[34]), .ZN(n38) );
  OAI22D1BWP30P140 U105 ( .A1(n43), .A2(n58), .B1(n46), .B2(n38), .ZN(N289) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U108 ( .A1(n47), .A2(n60), .B1(n46), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[5]), .ZN(n61) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[37]), .ZN(n40) );
  OAI22D1BWP30P140 U111 ( .A1(n47), .A2(n61), .B1(n46), .B2(n40), .ZN(N292) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[0]), .ZN(n64) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[32]), .ZN(n41) );
  OAI22D1BWP30P140 U114 ( .A1(n43), .A2(n64), .B1(n46), .B2(n41), .ZN(N287) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[1]), .ZN(n65) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[33]), .ZN(n42) );
  OAI22D1BWP30P140 U117 ( .A1(n43), .A2(n65), .B1(n46), .B2(n42), .ZN(N288) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[6]), .ZN(n62) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[38]), .ZN(n44) );
  OAI22D1BWP30P140 U120 ( .A1(n47), .A2(n62), .B1(n46), .B2(n44), .ZN(N293) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[7]), .ZN(n63) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[39]), .ZN(n45) );
  OAI22D1BWP30P140 U123 ( .A1(n47), .A2(n63), .B1(n46), .B2(n45), .ZN(N294) );
  INVD1BWP30P140 U124 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U125 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U126 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U127 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  MUX2NUD1BWP30P140 U128 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U129 ( .A1(n58), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U130 ( .A1(n59), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U131 ( .A1(n60), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U132 ( .A1(n61), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U133 ( .A1(n62), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U134 ( .A1(n63), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U135 ( .A1(n64), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U136 ( .A1(n65), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  INVD2BWP30P140 U137 ( .I(n79), .ZN(n77) );
  MOAI22D1BWP30P140 U138 ( .A1(n66), .A2(n77), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U139 ( .A1(n67), .A2(n77), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U140 ( .A1(n68), .A2(n77), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U141 ( .A1(n69), .A2(n77), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U142 ( .A1(n70), .A2(n77), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U143 ( .A1(n71), .A2(n77), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U144 ( .A1(n72), .A2(n77), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U145 ( .A1(n73), .A2(n77), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U146 ( .A1(n74), .A2(n77), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U147 ( .A1(n75), .A2(n77), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U148 ( .A1(n76), .A2(n77), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U149 ( .A1(n78), .A2(n77), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n92), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_128 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n20), .A2(n19), .B1(n31), .B2(n78), .ZN(N306) );
  INVD2BWP30P140 U4 ( .I(n36), .ZN(n46) );
  OAI22D1BWP30P140 U5 ( .A1(n47), .A2(n65), .B1(n46), .B2(n45), .ZN(N287) );
  INVD1BWP30P140 U6 ( .I(n57), .ZN(n79) );
  ND2D1BWP30P140 U7 ( .A1(n2), .A2(i_en), .ZN(n52) );
  INVD1BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n35) );
  CKBD1BWP30P140 U9 ( .I(n57), .Z(n1) );
  INVD1BWP30P140 U10 ( .I(n91), .ZN(n50) );
  OAI22D1BWP30P140 U11 ( .A1(n20), .A2(n7), .B1(n42), .B2(n66), .ZN(N295) );
  OAI22D1BWP30P140 U12 ( .A1(n20), .A2(n8), .B1(n42), .B2(n67), .ZN(N296) );
  OAI22D1BWP30P140 U13 ( .A1(n20), .A2(n9), .B1(n42), .B2(n68), .ZN(N297) );
  OAI22D1BWP30P140 U14 ( .A1(n20), .A2(n10), .B1(n42), .B2(n69), .ZN(N298) );
  OAI22D1BWP30P140 U15 ( .A1(n20), .A2(n11), .B1(n42), .B2(n70), .ZN(N299) );
  OAI22D1BWP30P140 U16 ( .A1(n20), .A2(n12), .B1(n42), .B2(n71), .ZN(N300) );
  OAI22D1BWP30P140 U17 ( .A1(n20), .A2(n17), .B1(n42), .B2(n72), .ZN(N301) );
  OAI22D1BWP30P140 U18 ( .A1(n20), .A2(n13), .B1(n42), .B2(n73), .ZN(N302) );
  OAI22D1BWP30P140 U19 ( .A1(n20), .A2(n14), .B1(n42), .B2(n74), .ZN(N303) );
  OAI22D1BWP30P140 U20 ( .A1(n20), .A2(n15), .B1(n42), .B2(n75), .ZN(N304) );
  OAI22D1BWP30P140 U21 ( .A1(n20), .A2(n16), .B1(n42), .B2(n76), .ZN(N305) );
  OAI22D1BWP30P140 U22 ( .A1(n33), .A2(n21), .B1(n31), .B2(n80), .ZN(N307) );
  OAI22D1BWP30P140 U23 ( .A1(n33), .A2(n22), .B1(n31), .B2(n81), .ZN(N308) );
  OAI22D1BWP30P140 U24 ( .A1(n33), .A2(n23), .B1(n31), .B2(n82), .ZN(N309) );
  OAI22D1BWP30P140 U25 ( .A1(n33), .A2(n24), .B1(n31), .B2(n83), .ZN(N310) );
  OAI22D1BWP30P140 U26 ( .A1(n33), .A2(n25), .B1(n31), .B2(n84), .ZN(N311) );
  OAI22D1BWP30P140 U27 ( .A1(n33), .A2(n26), .B1(n31), .B2(n85), .ZN(N312) );
  OAI22D1BWP30P140 U28 ( .A1(n33), .A2(n27), .B1(n31), .B2(n86), .ZN(N313) );
  OAI22D1BWP30P140 U29 ( .A1(n33), .A2(n28), .B1(n31), .B2(n87), .ZN(N314) );
  OAI22D1BWP30P140 U30 ( .A1(n33), .A2(n29), .B1(n31), .B2(n88), .ZN(N315) );
  OAI22D1BWP30P140 U31 ( .A1(n33), .A2(n30), .B1(n31), .B2(n89), .ZN(N316) );
  OAI22D1BWP30P140 U32 ( .A1(n33), .A2(n32), .B1(n31), .B2(n90), .ZN(N317) );
  OAI22D1BWP30P140 U33 ( .A1(n33), .A2(n18), .B1(n31), .B2(n93), .ZN(N318) );
  CKND2D2BWP30P140 U34 ( .A1(n56), .A2(n55), .ZN(n57) );
  INVD1BWP30P140 U35 ( .I(rst), .ZN(n2) );
  NR2D1BWP30P140 U36 ( .A1(n52), .A2(n35), .ZN(n4) );
  INVD1BWP30P140 U37 ( .I(i_valid[0]), .ZN(n54) );
  INVD2BWP30P140 U38 ( .I(i_valid[1]), .ZN(n53) );
  MUX2NUD1BWP30P140 U39 ( .I0(n54), .I1(n53), .S(i_cmd[1]), .ZN(n3) );
  ND2OPTIBD1BWP30P140 U40 ( .A1(n4), .A2(n3), .ZN(n5) );
  INVD2BWP30P140 U41 ( .I(n5), .ZN(n36) );
  INVD2BWP30P140 U42 ( .I(n36), .ZN(n20) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[40]), .ZN(n7) );
  INR2D1BWP30P140 U44 ( .A1(i_valid[0]), .B1(n52), .ZN(n48) );
  CKND2D2BWP30P140 U45 ( .A1(n48), .A2(n35), .ZN(n6) );
  INVD2BWP30P140 U46 ( .I(n6), .ZN(n34) );
  INVD2BWP30P140 U47 ( .I(n34), .ZN(n42) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[8]), .ZN(n66) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[41]), .ZN(n8) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[9]), .ZN(n67) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[42]), .ZN(n9) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[10]), .ZN(n68) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[43]), .ZN(n10) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[11]), .ZN(n69) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[44]), .ZN(n11) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[12]), .ZN(n70) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[45]), .ZN(n12) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[13]), .ZN(n71) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[47]), .ZN(n13) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[15]), .ZN(n73) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[48]), .ZN(n14) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[16]), .ZN(n74) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[49]), .ZN(n15) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[17]), .ZN(n75) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[50]), .ZN(n16) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[18]), .ZN(n76) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[46]), .ZN(n17) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[14]), .ZN(n72) );
  INVD2BWP30P140 U69 ( .I(n36), .ZN(n33) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[63]), .ZN(n18) );
  INVD2BWP30P140 U71 ( .I(n34), .ZN(n31) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[31]), .ZN(n93) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[51]), .ZN(n19) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[19]), .ZN(n78) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[52]), .ZN(n21) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[20]), .ZN(n80) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[53]), .ZN(n22) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[21]), .ZN(n81) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[54]), .ZN(n23) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[22]), .ZN(n82) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[55]), .ZN(n24) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[23]), .ZN(n83) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[56]), .ZN(n25) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[24]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[57]), .ZN(n26) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[25]), .ZN(n85) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[58]), .ZN(n27) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[26]), .ZN(n86) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[59]), .ZN(n28) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[27]), .ZN(n87) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[60]), .ZN(n29) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[28]), .ZN(n88) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[61]), .ZN(n30) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[29]), .ZN(n89) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[62]), .ZN(n32) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[30]), .ZN(n90) );
  INVD1BWP30P140 U97 ( .I(n34), .ZN(n47) );
  OAI31D1BWP30P140 U98 ( .A1(n52), .A2(n53), .A3(n35), .B(n47), .ZN(N353) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[7]), .ZN(n60) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[39]), .ZN(n37) );
  OAI22D1BWP30P140 U101 ( .A1(n42), .A2(n60), .B1(n46), .B2(n37), .ZN(N294) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[6]), .ZN(n59) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[38]), .ZN(n38) );
  OAI22D1BWP30P140 U104 ( .A1(n42), .A2(n59), .B1(n46), .B2(n38), .ZN(N293) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[5]), .ZN(n58) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[37]), .ZN(n39) );
  OAI22D1BWP30P140 U107 ( .A1(n42), .A2(n58), .B1(n46), .B2(n39), .ZN(N292) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[3]), .ZN(n62) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[35]), .ZN(n40) );
  OAI22D1BWP30P140 U110 ( .A1(n47), .A2(n62), .B1(n46), .B2(n40), .ZN(N290) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[4]), .ZN(n63) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[36]), .ZN(n41) );
  OAI22D1BWP30P140 U113 ( .A1(n42), .A2(n63), .B1(n46), .B2(n41), .ZN(N291) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[1]), .ZN(n64) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[33]), .ZN(n43) );
  OAI22D1BWP30P140 U116 ( .A1(n47), .A2(n64), .B1(n46), .B2(n43), .ZN(N288) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[2]), .ZN(n61) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[34]), .ZN(n44) );
  OAI22D1BWP30P140 U119 ( .A1(n47), .A2(n61), .B1(n46), .B2(n44), .ZN(N289) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[0]), .ZN(n65) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[32]), .ZN(n45) );
  INVD1BWP30P140 U122 ( .I(n48), .ZN(n51) );
  INVD1BWP30P140 U123 ( .I(n52), .ZN(n49) );
  AN3D4BWP30P140 U124 ( .A1(i_valid[1]), .A2(i_cmd[1]), .A3(n49), .Z(n91) );
  OAI21D1BWP30P140 U125 ( .A1(n51), .A2(i_cmd[1]), .B(n50), .ZN(N354) );
  NR2D1BWP30P140 U126 ( .A1(n52), .A2(i_cmd[1]), .ZN(n56) );
  MUX2NUD1BWP30P140 U127 ( .I0(n54), .I1(n53), .S(i_cmd[0]), .ZN(n55) );
  MOAI22D1BWP30P140 U128 ( .A1(n58), .A2(n1), .B1(i_data_bus[37]), .B2(n91), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U129 ( .A1(n59), .A2(n1), .B1(i_data_bus[38]), .B2(n91), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U130 ( .A1(n60), .A2(n1), .B1(i_data_bus[39]), .B2(n91), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U131 ( .A1(n61), .A2(n1), .B1(i_data_bus[34]), .B2(n91), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U132 ( .A1(n62), .A2(n1), .B1(i_data_bus[35]), .B2(n91), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U133 ( .A1(n63), .A2(n1), .B1(i_data_bus[36]), .B2(n91), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U134 ( .A1(n64), .A2(n1), .B1(i_data_bus[33]), .B2(n91), 
        .ZN(N320) );
  MOAI22D1BWP30P140 U135 ( .A1(n65), .A2(n1), .B1(i_data_bus[32]), .B2(n91), 
        .ZN(N319) );
  INVD2BWP30P140 U136 ( .I(n79), .ZN(n77) );
  MOAI22D1BWP30P140 U137 ( .A1(n66), .A2(n77), .B1(i_data_bus[40]), .B2(n91), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U138 ( .A1(n67), .A2(n77), .B1(i_data_bus[41]), .B2(n91), 
        .ZN(N328) );
  MOAI22D1BWP30P140 U139 ( .A1(n68), .A2(n77), .B1(i_data_bus[42]), .B2(n91), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U140 ( .A1(n69), .A2(n77), .B1(i_data_bus[43]), .B2(n91), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U141 ( .A1(n70), .A2(n77), .B1(i_data_bus[44]), .B2(n91), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U142 ( .A1(n71), .A2(n77), .B1(i_data_bus[45]), .B2(n91), 
        .ZN(N332) );
  MOAI22D1BWP30P140 U143 ( .A1(n72), .A2(n77), .B1(i_data_bus[46]), .B2(n91), 
        .ZN(N333) );
  MOAI22D1BWP30P140 U144 ( .A1(n73), .A2(n77), .B1(i_data_bus[47]), .B2(n91), 
        .ZN(N334) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n77), .B1(i_data_bus[48]), .B2(n91), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U146 ( .A1(n75), .A2(n77), .B1(i_data_bus[49]), .B2(n91), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U147 ( .A1(n76), .A2(n77), .B1(i_data_bus[50]), .B2(n91), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U148 ( .A1(n78), .A2(n77), .B1(i_data_bus[51]), .B2(n91), 
        .ZN(N338) );
  INVD2BWP30P140 U149 ( .I(n79), .ZN(n92) );
  MOAI22D1BWP30P140 U150 ( .A1(n80), .A2(n92), .B1(i_data_bus[52]), .B2(n91), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U151 ( .A1(n81), .A2(n92), .B1(i_data_bus[53]), .B2(n91), 
        .ZN(N340) );
  MOAI22D1BWP30P140 U152 ( .A1(n82), .A2(n92), .B1(i_data_bus[54]), .B2(n91), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U153 ( .A1(n83), .A2(n92), .B1(i_data_bus[55]), .B2(n91), 
        .ZN(N342) );
  MOAI22D1BWP30P140 U154 ( .A1(n84), .A2(n92), .B1(i_data_bus[56]), .B2(n91), 
        .ZN(N343) );
  MOAI22D1BWP30P140 U155 ( .A1(n85), .A2(n92), .B1(i_data_bus[57]), .B2(n91), 
        .ZN(N344) );
  MOAI22D1BWP30P140 U156 ( .A1(n86), .A2(n92), .B1(i_data_bus[58]), .B2(n91), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U157 ( .A1(n87), .A2(n92), .B1(i_data_bus[59]), .B2(n91), 
        .ZN(N346) );
  MOAI22D1BWP30P140 U158 ( .A1(n88), .A2(n92), .B1(i_data_bus[60]), .B2(n91), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U159 ( .A1(n89), .A2(n92), .B1(i_data_bus[61]), .B2(n91), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U160 ( .A1(n90), .A2(n92), .B1(i_data_bus[62]), .B2(n91), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U161 ( .A1(n93), .A2(n92), .B1(i_data_bus[63]), .B2(n91), 
        .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_129 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  NR2D2BWP30P140 U3 ( .A1(i_cmd[1]), .A2(n33), .ZN(n7) );
  INVD4BWP30P140 U4 ( .I(i_cmd[1]), .ZN(n12) );
  BUFFD4BWP30P140 U5 ( .I(n70), .Z(n67) );
  ND2OPTPAD4BWP30P140 U6 ( .A1(n6), .A2(n7), .ZN(n70) );
  ND2OPTIBD12BWP30P140 U7 ( .A1(n28), .A2(n31), .ZN(n72) );
  INVD2BWP30P140 U8 ( .I(i_valid[0]), .ZN(n13) );
  INR2D6BWP30P140 U9 ( .A1(n16), .B1(n1), .ZN(n28) );
  INVD3BWP30P140 U10 ( .I(i_valid[0]), .ZN(n1) );
  INVD2BWP30P140 U11 ( .I(i_valid[1]), .ZN(n5) );
  ND2OPTIBD1BWP30P140 U12 ( .A1(n3), .A2(i_data_bus[49]), .ZN(n27) );
  CKND2D4BWP30P140 U13 ( .A1(n15), .A2(n14), .ZN(n2) );
  INVD1BWP30P140 U14 ( .I(n2), .ZN(n3) );
  INVD3BWP30P140 U15 ( .I(n70), .ZN(n36) );
  ND2D1BWP30P140 U16 ( .A1(n27), .A2(n26), .ZN(N304) );
  OR2D1BWP30P140 U17 ( .A1(n72), .A2(n51), .Z(n26) );
  ND2OPTIBD8BWP30P140 U18 ( .A1(n15), .A2(n14), .ZN(n92) );
  ND2D1BWP30P140 U19 ( .A1(n10), .A2(n9), .ZN(N349) );
  ND2D1BWP30P140 U20 ( .A1(n69), .A2(i_data_bus[62]), .ZN(n9) );
  ND2D1BWP30P140 U21 ( .A1(n36), .A2(i_data_bus[30]), .ZN(n10) );
  INVD1BWP30P140 U22 ( .I(rst), .ZN(n4) );
  ND2D1BWP30P140 U23 ( .A1(n4), .A2(i_en), .ZN(n33) );
  MUX2NOPTD4BWP30P140 U24 ( .I0(n13), .I1(n5), .S(i_cmd[0]), .ZN(n6) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[30]), .ZN(n18) );
  INVD1BWP30P140 U26 ( .I(n33), .ZN(n16) );
  ND2OPTIBD4BWP30P140 U27 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n8) );
  INR2D8BWP30P140 U28 ( .A1(n16), .B1(n8), .ZN(n69) );
  INVD1BWP30P140 U29 ( .I(i_cmd[0]), .ZN(n11) );
  NR2OPTPAD2BWP30P140 U30 ( .A1(n11), .A2(n33), .ZN(n15) );
  INVD2BWP30P140 U31 ( .I(i_valid[1]), .ZN(n32) );
  MUX2NOPTD4BWP30P140 U32 ( .I0(n32), .I1(n13), .S(n12), .ZN(n14) );
  INVD1BWP30P140 U33 ( .I(i_data_bus[63]), .ZN(n17) );
  INVD2BWP30P140 U34 ( .I(i_cmd[0]), .ZN(n31) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[31]), .ZN(n68) );
  OAI22OPTPBD1BWP30P140 U36 ( .A1(n92), .A2(n17), .B1(n72), .B2(n68), .ZN(N318) );
  INVD1BWP30P140 U37 ( .I(i_data_bus[62]), .ZN(n19) );
  OAI22OPTPBD1BWP30P140 U38 ( .A1(n92), .A2(n19), .B1(n72), .B2(n18), .ZN(N317) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[61]), .ZN(n20) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[29]), .ZN(n66) );
  OAI22OPTPBD1BWP30P140 U41 ( .A1(n92), .A2(n20), .B1(n72), .B2(n66), .ZN(N316) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[38]), .ZN(n21) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[6]), .ZN(n44) );
  OAI22OPTPBD1BWP30P140 U44 ( .A1(n92), .A2(n21), .B1(n72), .B2(n44), .ZN(N293) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[36]), .ZN(n22) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[4]), .ZN(n46) );
  OAI22OPTPBD1BWP30P140 U47 ( .A1(n92), .A2(n22), .B1(n72), .B2(n46), .ZN(N291) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[39]), .ZN(n23) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[7]), .ZN(n71) );
  OAI22OPTPBD1BWP30P140 U50 ( .A1(n92), .A2(n23), .B1(n72), .B2(n71), .ZN(N294) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[37]), .ZN(n24) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[5]), .ZN(n45) );
  OAI22OPTPBD1BWP30P140 U53 ( .A1(n92), .A2(n24), .B1(n72), .B2(n45), .ZN(N292) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[35]), .ZN(n25) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[3]), .ZN(n47) );
  OAI22OPTPBD1BWP30P140 U56 ( .A1(n92), .A2(n25), .B1(n72), .B2(n47), .ZN(N290) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[17]), .ZN(n51) );
  INVD1BWP30P140 U58 ( .I(n28), .ZN(n30) );
  INVD1BWP30P140 U59 ( .I(n69), .ZN(n29) );
  OAI21D1BWP30P140 U60 ( .A1(n30), .A2(i_cmd[1]), .B(n29), .ZN(N354) );
  OAI31D1BWP30P140 U61 ( .A1(n33), .A2(n32), .A3(n31), .B(n72), .ZN(N353) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[19]), .ZN(n53) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[51]), .ZN(n34) );
  OAI22D1BWP30P140 U64 ( .A1(n72), .A2(n53), .B1(n2), .B2(n34), .ZN(N306) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[18]), .ZN(n52) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[50]), .ZN(n35) );
  OAI22D1BWP30P140 U67 ( .A1(n72), .A2(n52), .B1(n2), .B2(n35), .ZN(N305) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[14]), .ZN(n37) );
  INVD4BWP30P140 U69 ( .I(n36), .ZN(n62) );
  MOAI22D1BWP30P140 U70 ( .A1(n37), .A2(n62), .B1(i_data_bus[46]), .B2(n69), 
        .ZN(N333) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[13]), .ZN(n38) );
  MOAI22D1BWP30P140 U72 ( .A1(n38), .A2(n67), .B1(i_data_bus[45]), .B2(n69), 
        .ZN(N332) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[12]), .ZN(n39) );
  MOAI22D1BWP30P140 U74 ( .A1(n39), .A2(n62), .B1(i_data_bus[44]), .B2(n69), 
        .ZN(N331) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[11]), .ZN(n40) );
  MOAI22D1BWP30P140 U76 ( .A1(n40), .A2(n67), .B1(i_data_bus[43]), .B2(n69), 
        .ZN(N330) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[10]), .ZN(n41) );
  MOAI22D1BWP30P140 U78 ( .A1(n41), .A2(n62), .B1(i_data_bus[42]), .B2(n69), 
        .ZN(N329) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[9]), .ZN(n42) );
  MOAI22D1BWP30P140 U80 ( .A1(n42), .A2(n67), .B1(i_data_bus[41]), .B2(n69), 
        .ZN(N328) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[8]), .ZN(n43) );
  MOAI22D1BWP30P140 U82 ( .A1(n43), .A2(n62), .B1(i_data_bus[40]), .B2(n69), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U83 ( .A1(n44), .A2(n62), .B1(i_data_bus[38]), .B2(n69), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U84 ( .A1(n45), .A2(n62), .B1(i_data_bus[37]), .B2(n69), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U85 ( .A1(n46), .A2(n62), .B1(i_data_bus[36]), .B2(n69), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U86 ( .A1(n47), .A2(n62), .B1(i_data_bus[35]), .B2(n69), 
        .ZN(N322) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[2]), .ZN(n48) );
  MOAI22D1BWP30P140 U88 ( .A1(n48), .A2(n62), .B1(i_data_bus[34]), .B2(n69), 
        .ZN(N321) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[15]), .ZN(n49) );
  MOAI22D1BWP30P140 U90 ( .A1(n49), .A2(n67), .B1(i_data_bus[47]), .B2(n69), 
        .ZN(N334) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[16]), .ZN(n50) );
  MOAI22D1BWP30P140 U92 ( .A1(n50), .A2(n62), .B1(i_data_bus[48]), .B2(n69), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U93 ( .A1(n51), .A2(n62), .B1(i_data_bus[49]), .B2(n69), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U94 ( .A1(n52), .A2(n62), .B1(i_data_bus[50]), .B2(n69), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U95 ( .A1(n53), .A2(n62), .B1(i_data_bus[51]), .B2(n69), 
        .ZN(N338) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[20]), .ZN(n54) );
  MOAI22D1BWP30P140 U97 ( .A1(n54), .A2(n62), .B1(i_data_bus[52]), .B2(n69), 
        .ZN(N339) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[21]), .ZN(n55) );
  MOAI22D1BWP30P140 U99 ( .A1(n55), .A2(n67), .B1(i_data_bus[53]), .B2(n69), 
        .ZN(N340) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[22]), .ZN(n56) );
  MOAI22D1BWP30P140 U101 ( .A1(n56), .A2(n67), .B1(i_data_bus[54]), .B2(n69), 
        .ZN(N341) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[23]), .ZN(n57) );
  MOAI22D1BWP30P140 U103 ( .A1(n57), .A2(n67), .B1(i_data_bus[55]), .B2(n69), 
        .ZN(N342) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[24]), .ZN(n58) );
  MOAI22D1BWP30P140 U105 ( .A1(n58), .A2(n67), .B1(i_data_bus[56]), .B2(n69), 
        .ZN(N343) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[25]), .ZN(n59) );
  MOAI22D1BWP30P140 U107 ( .A1(n59), .A2(n67), .B1(i_data_bus[57]), .B2(n69), 
        .ZN(N344) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[26]), .ZN(n60) );
  MOAI22D1BWP30P140 U109 ( .A1(n60), .A2(n67), .B1(i_data_bus[58]), .B2(n69), 
        .ZN(N345) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[1]), .ZN(n61) );
  MOAI22D1BWP30P140 U111 ( .A1(n61), .A2(n62), .B1(i_data_bus[33]), .B2(n69), 
        .ZN(N320) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[0]), .ZN(n63) );
  MOAI22D1BWP30P140 U113 ( .A1(n63), .A2(n62), .B1(i_data_bus[32]), .B2(n69), 
        .ZN(N319) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[27]), .ZN(n64) );
  MOAI22D1BWP30P140 U115 ( .A1(n64), .A2(n67), .B1(i_data_bus[59]), .B2(n69), 
        .ZN(N346) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[28]), .ZN(n65) );
  MOAI22D1BWP30P140 U117 ( .A1(n65), .A2(n67), .B1(i_data_bus[60]), .B2(n69), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U118 ( .A1(n66), .A2(n67), .B1(i_data_bus[61]), .B2(n69), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U119 ( .A1(n68), .A2(n67), .B1(i_data_bus[63]), .B2(n69), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U120 ( .A1(n71), .A2(n70), .B1(i_data_bus[39]), .B2(n69), 
        .ZN(N326) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[60]), .ZN(n73) );
  INVD8BWP30P140 U122 ( .I(n72), .ZN(n94) );
  MOAI22D1BWP30P140 U123 ( .A1(n92), .A2(n73), .B1(n94), .B2(i_data_bus[28]), 
        .ZN(N315) );
  INVD1BWP30P140 U124 ( .I(i_data_bus[48]), .ZN(n74) );
  MOAI22D1BWP30P140 U125 ( .A1(n92), .A2(n74), .B1(n94), .B2(i_data_bus[16]), 
        .ZN(N303) );
  INVD1BWP30P140 U126 ( .I(i_data_bus[34]), .ZN(n75) );
  MOAI22D1BWP30P140 U127 ( .A1(n92), .A2(n75), .B1(n94), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140 U128 ( .I(i_data_bus[59]), .ZN(n76) );
  MOAI22D1BWP30P140 U129 ( .A1(n92), .A2(n76), .B1(n94), .B2(i_data_bus[27]), 
        .ZN(N314) );
  INVD1BWP30P140 U130 ( .I(i_data_bus[47]), .ZN(n77) );
  MOAI22D1BWP30P140 U131 ( .A1(n92), .A2(n77), .B1(n94), .B2(i_data_bus[15]), 
        .ZN(N302) );
  INVD1BWP30P140 U132 ( .I(i_data_bus[33]), .ZN(n78) );
  MOAI22D1BWP30P140 U133 ( .A1(n92), .A2(n78), .B1(n94), .B2(i_data_bus[1]), 
        .ZN(N288) );
  INVD1BWP30P140 U134 ( .I(i_data_bus[58]), .ZN(n79) );
  MOAI22D1BWP30P140 U135 ( .A1(n92), .A2(n79), .B1(n94), .B2(i_data_bus[26]), 
        .ZN(N313) );
  INVD1BWP30P140 U136 ( .I(i_data_bus[46]), .ZN(n80) );
  MOAI22D1BWP30P140 U137 ( .A1(n92), .A2(n80), .B1(n94), .B2(i_data_bus[14]), 
        .ZN(N301) );
  INVD1BWP30P140 U138 ( .I(i_data_bus[32]), .ZN(n81) );
  MOAI22D1BWP30P140 U139 ( .A1(n92), .A2(n81), .B1(n94), .B2(i_data_bus[0]), 
        .ZN(N287) );
  INVD1BWP30P140 U140 ( .I(i_data_bus[57]), .ZN(n82) );
  MOAI22D1BWP30P140 U141 ( .A1(n92), .A2(n82), .B1(n94), .B2(i_data_bus[25]), 
        .ZN(N312) );
  INVD1BWP30P140 U142 ( .I(i_data_bus[45]), .ZN(n83) );
  MOAI22D1BWP30P140 U143 ( .A1(n92), .A2(n83), .B1(n94), .B2(i_data_bus[13]), 
        .ZN(N300) );
  INVD1BWP30P140 U144 ( .I(i_data_bus[56]), .ZN(n84) );
  MOAI22D1BWP30P140 U145 ( .A1(n92), .A2(n84), .B1(n94), .B2(i_data_bus[24]), 
        .ZN(N311) );
  INVD1BWP30P140 U146 ( .I(i_data_bus[44]), .ZN(n85) );
  MOAI22D1BWP30P140 U147 ( .A1(n92), .A2(n85), .B1(n94), .B2(i_data_bus[12]), 
        .ZN(N299) );
  INVD1BWP30P140 U148 ( .I(i_data_bus[55]), .ZN(n86) );
  MOAI22D1BWP30P140 U149 ( .A1(n92), .A2(n86), .B1(n94), .B2(i_data_bus[23]), 
        .ZN(N310) );
  INVD1BWP30P140 U150 ( .I(i_data_bus[43]), .ZN(n87) );
  MOAI22D1BWP30P140 U151 ( .A1(n92), .A2(n87), .B1(n94), .B2(i_data_bus[11]), 
        .ZN(N298) );
  INVD1BWP30P140 U152 ( .I(i_data_bus[54]), .ZN(n88) );
  MOAI22D1BWP30P140 U153 ( .A1(n92), .A2(n88), .B1(n94), .B2(i_data_bus[22]), 
        .ZN(N309) );
  INVD1BWP30P140 U154 ( .I(i_data_bus[42]), .ZN(n89) );
  MOAI22D1BWP30P140 U155 ( .A1(n92), .A2(n89), .B1(n94), .B2(i_data_bus[10]), 
        .ZN(N297) );
  INVD1BWP30P140 U156 ( .I(i_data_bus[53]), .ZN(n90) );
  MOAI22D1BWP30P140 U157 ( .A1(n92), .A2(n90), .B1(n94), .B2(i_data_bus[21]), 
        .ZN(N308) );
  INVD1BWP30P140 U158 ( .I(i_data_bus[41]), .ZN(n91) );
  MOAI22D1BWP30P140 U159 ( .A1(n92), .A2(n91), .B1(n94), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140 U160 ( .I(i_data_bus[52]), .ZN(n93) );
  MOAI22D1BWP30P140 U161 ( .A1(n92), .A2(n93), .B1(n94), .B2(i_data_bus[20]), 
        .ZN(N307) );
  INVD1BWP30P140 U162 ( .I(i_data_bus[40]), .ZN(n95) );
  MOAI22D1BWP30P140 U163 ( .A1(n2), .A2(n95), .B1(n94), .B2(i_data_bus[8]), 
        .ZN(N295) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_130 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  MOAI22D1BWP30P140 U3 ( .A1(n23), .A2(n12), .B1(i_data_bus[35]), .B2(n7), 
        .ZN(N322) );
  ND2OPTIBD1BWP30P140 U4 ( .A1(n71), .A2(i_data_bus[61]), .ZN(n6) );
  NR2OPTPAD6BWP30P140 U5 ( .A1(n13), .A2(n35), .ZN(n7) );
  CKND2D3BWP30P140 U6 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n13) );
  INVD1BWP30P140 U7 ( .I(n4), .ZN(n3) );
  BUFFD4BWP30P140 U8 ( .I(n69), .Z(n2) );
  INVD6BWP30P140 U9 ( .I(n92), .ZN(n71) );
  INVD3BWP30P140 U10 ( .I(i_cmd[1]), .ZN(n15) );
  INVD2BWP30P140 U11 ( .I(i_valid[0]), .ZN(n5) );
  ND2OPTPAD4BWP30P140 U12 ( .A1(n29), .A2(n33), .ZN(n69) );
  INVD2BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n14) );
  BUFFD4BWP30P140 U14 ( .I(n69), .Z(n1) );
  ND2OPTIBD6BWP30P140 U15 ( .A1(n17), .A2(n18), .ZN(n92) );
  ND2D1BWP30P140 U16 ( .A1(n6), .A2(n3), .ZN(N316) );
  NR2D1BWP30P140 U17 ( .A1(n1), .A2(n49), .ZN(n4) );
  INVD2BWP30P140 U18 ( .I(i_cmd[0]), .ZN(n33) );
  INR2D2BWP30P140 U19 ( .A1(n19), .B1(n5), .ZN(n29) );
  INVD1BWP30P140 U20 ( .I(n7), .ZN(n31) );
  ND2OPTPAD6BWP30P140 U21 ( .A1(n11), .A2(n10), .ZN(n12) );
  INVD1BWP30P140 U22 ( .I(i_data_bus[3]), .ZN(n23) );
  INVD2BWP30P140 U23 ( .I(n15), .ZN(n30) );
  INVD1BWP30P140 U24 ( .I(rst), .ZN(n8) );
  ND2D1BWP30P140 U25 ( .A1(n8), .A2(i_en), .ZN(n35) );
  NR2OPTPAD2BWP30P140 U26 ( .A1(n30), .A2(n35), .ZN(n11) );
  INVD3BWP30P140 U27 ( .I(i_valid[0]), .ZN(n16) );
  INVD2BWP30P140 U28 ( .I(i_valid[1]), .ZN(n9) );
  MUX2NOPTD4BWP30P140 U29 ( .I0(n16), .I1(n9), .S(i_cmd[0]), .ZN(n10) );
  INVD1BWP30P140 U30 ( .I(n35), .ZN(n19) );
  NR2OPTPAD2BWP30P140 U31 ( .A1(n14), .A2(n35), .ZN(n18) );
  INVD2BWP30P140 U32 ( .I(i_valid[1]), .ZN(n34) );
  MUX2NOPTD4BWP30P140 U33 ( .I0(n34), .I1(n16), .S(n15), .ZN(n17) );
  INVD6BWP30P140 U34 ( .I(n71), .ZN(n74) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[49]), .ZN(n20) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[17]), .ZN(n56) );
  OAI22OPTPBD1BWP30P140 U37 ( .A1(n74), .A2(n20), .B1(n2), .B2(n56), .ZN(N304)
         );
  INVD1BWP30P140 U38 ( .I(i_data_bus[51]), .ZN(n21) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[19]), .ZN(n51) );
  OAI22OPTPBD1BWP30P140 U40 ( .A1(n74), .A2(n21), .B1(n2), .B2(n51), .ZN(N306)
         );
  INVD1BWP30P140 U41 ( .I(i_data_bus[50]), .ZN(n22) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[18]), .ZN(n57) );
  OAI22OPTPBD1BWP30P140 U43 ( .A1(n74), .A2(n22), .B1(n2), .B2(n57), .ZN(N305)
         );
  INVD1BWP30P140 U44 ( .I(i_data_bus[35]), .ZN(n24) );
  OAI22OPTPBD1BWP30P140 U45 ( .A1(n74), .A2(n24), .B1(n1), .B2(n23), .ZN(N290)
         );
  INVD1BWP30P140 U46 ( .I(i_data_bus[39]), .ZN(n25) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[7]), .ZN(n45) );
  OAI22OPTPBD1BWP30P140 U48 ( .A1(n74), .A2(n25), .B1(n2), .B2(n45), .ZN(N294)
         );
  INVD1BWP30P140 U49 ( .I(i_data_bus[37]), .ZN(n26) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[5]), .ZN(n64) );
  OAI22OPTPBD1BWP30P140 U51 ( .A1(n74), .A2(n26), .B1(n2), .B2(n64), .ZN(N292)
         );
  INVD1BWP30P140 U52 ( .I(i_data_bus[38]), .ZN(n27) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[6]), .ZN(n58) );
  OAI22OPTPBD1BWP30P140 U54 ( .A1(n74), .A2(n27), .B1(n2), .B2(n58), .ZN(N293)
         );
  INVD1BWP30P140 U55 ( .I(i_data_bus[36]), .ZN(n28) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[4]), .ZN(n42) );
  OAI22OPTPBD1BWP30P140 U57 ( .A1(n74), .A2(n28), .B1(n2), .B2(n42), .ZN(N291)
         );
  INVD1BWP30P140 U58 ( .I(i_data_bus[29]), .ZN(n49) );
  INVD1BWP30P140 U59 ( .I(n29), .ZN(n32) );
  OAI21D1BWP30P140 U60 ( .A1(n32), .A2(n30), .B(n31), .ZN(N354) );
  OAI31D1BWP30P140 U61 ( .A1(n35), .A2(n34), .A3(n33), .B(n2), .ZN(N353) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[30]), .ZN(n38) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[62]), .ZN(n36) );
  OAI22D1BWP30P140 U64 ( .A1(n2), .A2(n38), .B1(n92), .B2(n36), .ZN(N317) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[31]), .ZN(n66) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[63]), .ZN(n37) );
  OAI22D1BWP30P140 U67 ( .A1(n2), .A2(n66), .B1(n92), .B2(n37), .ZN(N318) );
  MOAI22D1BWP30P140 U68 ( .A1(n38), .A2(n12), .B1(i_data_bus[62]), .B2(n7), 
        .ZN(N349) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[1]), .ZN(n39) );
  MOAI22D1BWP30P140 U70 ( .A1(n39), .A2(n12), .B1(i_data_bus[33]), .B2(n7), 
        .ZN(N320) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[13]), .ZN(n40) );
  MOAI22D1BWP30P140 U72 ( .A1(n40), .A2(n12), .B1(i_data_bus[45]), .B2(n7), 
        .ZN(N332) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[0]), .ZN(n41) );
  MOAI22D1BWP30P140 U74 ( .A1(n41), .A2(n12), .B1(i_data_bus[32]), .B2(n7), 
        .ZN(N319) );
  MOAI22D1BWP30P140 U75 ( .A1(n42), .A2(n12), .B1(i_data_bus[36]), .B2(n7), 
        .ZN(N323) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[12]), .ZN(n43) );
  MOAI22D1BWP30P140 U77 ( .A1(n43), .A2(n12), .B1(i_data_bus[44]), .B2(n7), 
        .ZN(N331) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[11]), .ZN(n44) );
  MOAI22D1BWP30P140 U79 ( .A1(n44), .A2(n12), .B1(i_data_bus[43]), .B2(n7), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U80 ( .A1(n45), .A2(n12), .B1(i_data_bus[39]), .B2(n7), 
        .ZN(N326) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[28]), .ZN(n46) );
  MOAI22D1BWP30P140 U82 ( .A1(n46), .A2(n12), .B1(i_data_bus[60]), .B2(n7), 
        .ZN(N347) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[9]), .ZN(n47) );
  MOAI22D1BWP30P140 U84 ( .A1(n47), .A2(n12), .B1(i_data_bus[41]), .B2(n7), 
        .ZN(N328) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[8]), .ZN(n48) );
  MOAI22D1BWP30P140 U86 ( .A1(n48), .A2(n12), .B1(i_data_bus[40]), .B2(n7), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U87 ( .A1(n49), .A2(n12), .B1(i_data_bus[61]), .B2(n7), 
        .ZN(N348) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[10]), .ZN(n50) );
  MOAI22D1BWP30P140 U89 ( .A1(n50), .A2(n12), .B1(i_data_bus[42]), .B2(n7), 
        .ZN(N329) );
  MOAI22D1BWP30P140 U90 ( .A1(n51), .A2(n12), .B1(i_data_bus[51]), .B2(n7), 
        .ZN(N338) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[24]), .ZN(n52) );
  MOAI22D1BWP30P140 U92 ( .A1(n52), .A2(n12), .B1(i_data_bus[56]), .B2(n7), 
        .ZN(N343) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[14]), .ZN(n53) );
  MOAI22D1BWP30P140 U94 ( .A1(n53), .A2(n12), .B1(i_data_bus[46]), .B2(n7), 
        .ZN(N333) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[15]), .ZN(n54) );
  MOAI22D1BWP30P140 U96 ( .A1(n54), .A2(n12), .B1(i_data_bus[47]), .B2(n7), 
        .ZN(N334) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[16]), .ZN(n55) );
  MOAI22D1BWP30P140 U98 ( .A1(n55), .A2(n12), .B1(i_data_bus[48]), .B2(n7), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U99 ( .A1(n56), .A2(n12), .B1(i_data_bus[49]), .B2(n7), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U100 ( .A1(n57), .A2(n12), .B1(i_data_bus[50]), .B2(n7), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U101 ( .A1(n58), .A2(n12), .B1(i_data_bus[38]), .B2(n7), 
        .ZN(N325) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[20]), .ZN(n59) );
  MOAI22D1BWP30P140 U103 ( .A1(n59), .A2(n12), .B1(i_data_bus[52]), .B2(n7), 
        .ZN(N339) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[21]), .ZN(n60) );
  MOAI22D1BWP30P140 U105 ( .A1(n60), .A2(n12), .B1(i_data_bus[53]), .B2(n7), 
        .ZN(N340) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[2]), .ZN(n61) );
  MOAI22D1BWP30P140 U107 ( .A1(n61), .A2(n12), .B1(i_data_bus[34]), .B2(n7), 
        .ZN(N321) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[23]), .ZN(n62) );
  MOAI22D1BWP30P140 U109 ( .A1(n62), .A2(n12), .B1(i_data_bus[55]), .B2(n7), 
        .ZN(N342) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[26]), .ZN(n63) );
  MOAI22D1BWP30P140 U111 ( .A1(n63), .A2(n12), .B1(i_data_bus[58]), .B2(n7), 
        .ZN(N345) );
  MOAI22D1BWP30P140 U112 ( .A1(n64), .A2(n12), .B1(i_data_bus[37]), .B2(n7), 
        .ZN(N324) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[22]), .ZN(n65) );
  MOAI22D1BWP30P140 U114 ( .A1(n65), .A2(n12), .B1(i_data_bus[54]), .B2(n7), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U115 ( .A1(n66), .A2(n12), .B1(i_data_bus[63]), .B2(n7), 
        .ZN(N350) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[27]), .ZN(n67) );
  MOAI22D1BWP30P140 U117 ( .A1(n67), .A2(n12), .B1(i_data_bus[59]), .B2(n7), 
        .ZN(N346) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[25]), .ZN(n68) );
  MOAI22D1BWP30P140 U119 ( .A1(n68), .A2(n12), .B1(i_data_bus[57]), .B2(n7), 
        .ZN(N344) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[60]), .ZN(n70) );
  INVD4BWP30P140 U121 ( .I(n69), .ZN(n93) );
  MOAI22D1BWP30P140 U122 ( .A1(n74), .A2(n70), .B1(n93), .B2(i_data_bus[28]), 
        .ZN(N315) );
  INVD4BWP30P140 U123 ( .I(n71), .ZN(n95) );
  INVD1BWP30P140 U124 ( .I(i_data_bus[48]), .ZN(n72) );
  MOAI22D1BWP30P140 U125 ( .A1(n95), .A2(n72), .B1(n93), .B2(i_data_bus[16]), 
        .ZN(N303) );
  INVD1BWP30P140 U126 ( .I(i_data_bus[34]), .ZN(n73) );
  MOAI22D1BWP30P140 U127 ( .A1(n74), .A2(n73), .B1(n93), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140 U128 ( .I(i_data_bus[59]), .ZN(n75) );
  MOAI22D1BWP30P140 U129 ( .A1(n74), .A2(n75), .B1(n93), .B2(i_data_bus[27]), 
        .ZN(N314) );
  INVD1BWP30P140 U130 ( .I(i_data_bus[47]), .ZN(n76) );
  MOAI22D1BWP30P140 U131 ( .A1(n95), .A2(n76), .B1(n93), .B2(i_data_bus[15]), 
        .ZN(N302) );
  INVD1BWP30P140 U132 ( .I(i_data_bus[33]), .ZN(n77) );
  MOAI22D1BWP30P140 U133 ( .A1(n95), .A2(n77), .B1(n93), .B2(i_data_bus[1]), 
        .ZN(N288) );
  INVD1BWP30P140 U134 ( .I(i_data_bus[58]), .ZN(n78) );
  MOAI22D1BWP30P140 U135 ( .A1(n74), .A2(n78), .B1(n93), .B2(i_data_bus[26]), 
        .ZN(N313) );
  INVD1BWP30P140 U136 ( .I(i_data_bus[46]), .ZN(n79) );
  MOAI22D1BWP30P140 U137 ( .A1(n95), .A2(n79), .B1(n93), .B2(i_data_bus[14]), 
        .ZN(N301) );
  INVD1BWP30P140 U138 ( .I(i_data_bus[32]), .ZN(n80) );
  MOAI22D1BWP30P140 U139 ( .A1(n74), .A2(n80), .B1(n93), .B2(i_data_bus[0]), 
        .ZN(N287) );
  INVD1BWP30P140 U140 ( .I(i_data_bus[57]), .ZN(n81) );
  MOAI22D1BWP30P140 U141 ( .A1(n74), .A2(n81), .B1(n93), .B2(i_data_bus[25]), 
        .ZN(N312) );
  INVD1BWP30P140 U142 ( .I(i_data_bus[45]), .ZN(n82) );
  MOAI22D1BWP30P140 U143 ( .A1(n95), .A2(n82), .B1(n93), .B2(i_data_bus[13]), 
        .ZN(N300) );
  INVD1BWP30P140 U144 ( .I(i_data_bus[56]), .ZN(n83) );
  MOAI22D1BWP30P140 U145 ( .A1(n74), .A2(n83), .B1(n93), .B2(i_data_bus[24]), 
        .ZN(N311) );
  INVD1BWP30P140 U146 ( .I(i_data_bus[44]), .ZN(n84) );
  MOAI22D1BWP30P140 U147 ( .A1(n95), .A2(n84), .B1(n93), .B2(i_data_bus[12]), 
        .ZN(N299) );
  INVD1BWP30P140 U148 ( .I(i_data_bus[55]), .ZN(n85) );
  MOAI22D1BWP30P140 U149 ( .A1(n74), .A2(n85), .B1(n93), .B2(i_data_bus[23]), 
        .ZN(N310) );
  INVD1BWP30P140 U150 ( .I(i_data_bus[43]), .ZN(n86) );
  MOAI22D1BWP30P140 U151 ( .A1(n95), .A2(n86), .B1(n93), .B2(i_data_bus[11]), 
        .ZN(N298) );
  INVD1BWP30P140 U152 ( .I(i_data_bus[54]), .ZN(n87) );
  MOAI22D1BWP30P140 U153 ( .A1(n74), .A2(n87), .B1(n93), .B2(i_data_bus[22]), 
        .ZN(N309) );
  INVD1BWP30P140 U154 ( .I(i_data_bus[42]), .ZN(n88) );
  MOAI22D1BWP30P140 U155 ( .A1(n95), .A2(n88), .B1(n93), .B2(i_data_bus[10]), 
        .ZN(N297) );
  INVD1BWP30P140 U156 ( .I(i_data_bus[53]), .ZN(n89) );
  MOAI22D1BWP30P140 U157 ( .A1(n92), .A2(n89), .B1(n93), .B2(i_data_bus[21]), 
        .ZN(N308) );
  INVD1BWP30P140 U158 ( .I(i_data_bus[41]), .ZN(n90) );
  MOAI22D1BWP30P140 U159 ( .A1(n95), .A2(n90), .B1(n93), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140 U160 ( .I(i_data_bus[52]), .ZN(n91) );
  MOAI22D1BWP30P140 U161 ( .A1(n92), .A2(n91), .B1(n93), .B2(i_data_bus[20]), 
        .ZN(N307) );
  INVD1BWP30P140 U162 ( .I(i_data_bus[40]), .ZN(n94) );
  MOAI22D1BWP30P140 U163 ( .A1(n95), .A2(n94), .B1(n93), .B2(i_data_bus[8]), 
        .ZN(N295) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_131 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n105), .A2(n10), .B1(n98), .B2(n73), .ZN(N291) );
  OAI22D1BWP30P140 U4 ( .A1(n105), .A2(n11), .B1(n98), .B2(n30), .ZN(N292) );
  OAI22D1BWP30P140 U5 ( .A1(n105), .A2(n12), .B1(n98), .B2(n28), .ZN(N293) );
  OAI22D1BWP30P140 U6 ( .A1(n105), .A2(n13), .B1(n98), .B2(n44), .ZN(N290) );
  OAI22D1BWP30P140 U7 ( .A1(n105), .A2(n14), .B1(n98), .B2(n40), .ZN(N294) );
  OAI21D1BWP30P140 U8 ( .A1(n91), .A2(n71), .B(n70), .ZN(N343) );
  INVD9BWP30P140 U9 ( .I(n98), .ZN(n121) );
  INVD4BWP30P140 U10 ( .I(n123), .ZN(n97) );
  ND2OPTIBD6BWP30P140 U11 ( .A1(n5), .A2(n6), .ZN(n123) );
  INVD3BWP30P140 U12 ( .I(i_cmd[1]), .ZN(n15) );
  BUFFD4BWP30P140 U13 ( .I(n123), .Z(n1) );
  INVD4BWP30P140 U14 ( .I(n20), .ZN(n26) );
  INVD8BWP30P140 U15 ( .I(n26), .ZN(n91) );
  INVD4BWP30P140 U16 ( .I(n2), .ZN(n78) );
  INVD4BWP30P140 U17 ( .I(i_valid[0]), .ZN(n17) );
  INVD6BWP30P140 U18 ( .I(n26), .ZN(n95) );
  OAI21D2BWP30P140 U19 ( .A1(n95), .A2(n75), .B(n74), .ZN(N331) );
  CKND2D4BWP30P140 U20 ( .A1(i_valid[0]), .A2(n22), .ZN(n2) );
  ND2D1BWP30P140 U21 ( .A1(n77), .A2(n76), .ZN(N304) );
  ND2OPTPAD6BWP30P140 U22 ( .A1(n78), .A2(n82), .ZN(n98) );
  INVD8BWP30P140 U23 ( .I(n80), .ZN(n94) );
  CKND2D3BWP30P140 U24 ( .A1(n19), .A2(n18), .ZN(n20) );
  INVD1BWP30P140 U25 ( .I(i_cmd[0]), .ZN(n3) );
  NR2OPTPAD2BWP30P140 U26 ( .A1(n3), .A2(n84), .ZN(n6) );
  OR2D1BWP30P140 U27 ( .A1(n98), .A2(n93), .Z(n76) );
  ND2OPTIBD1BWP30P140 U28 ( .A1(n97), .A2(i_data_bus[49]), .ZN(n77) );
  ND2D1BWP30P140 U29 ( .A1(n94), .A2(i_data_bus[40]), .ZN(n31) );
  ND2D1BWP30P140 U30 ( .A1(n94), .A2(i_data_bus[42]), .ZN(n35) );
  ND2D1BWP30P140 U31 ( .A1(n94), .A2(i_data_bus[44]), .ZN(n74) );
  ND2D1BWP30P140 U32 ( .A1(n94), .A2(i_data_bus[45]), .ZN(n41) );
  ND2D1BWP30P140 U33 ( .A1(n94), .A2(i_data_bus[46]), .ZN(n64) );
  ND2D1BWP30P140 U34 ( .A1(n94), .A2(i_data_bus[47]), .ZN(n60) );
  ND2D1BWP30P140 U35 ( .A1(n94), .A2(i_data_bus[48]), .ZN(n47) );
  ND2D1BWP30P140 U36 ( .A1(n94), .A2(i_data_bus[50]), .ZN(n51) );
  ND2D1BWP30P140 U37 ( .A1(n94), .A2(i_data_bus[54]), .ZN(n58) );
  ND2D1BWP30P140 U38 ( .A1(n94), .A2(i_data_bus[55]), .ZN(n62) );
  ND2D1BWP30P140 U39 ( .A1(n94), .A2(i_data_bus[56]), .ZN(n70) );
  ND2D1BWP30P140 U40 ( .A1(n94), .A2(i_data_bus[57]), .ZN(n24) );
  ND2D1BWP30P140 U41 ( .A1(n94), .A2(i_data_bus[58]), .ZN(n33) );
  ND2D1BWP30P140 U42 ( .A1(n94), .A2(i_data_bus[59]), .ZN(n37) );
  ND2D1BWP30P140 U43 ( .A1(n94), .A2(i_data_bus[60]), .ZN(n45) );
  ND2D1BWP30P140 U44 ( .A1(n94), .A2(i_data_bus[61]), .ZN(n49) );
  ND2D1BWP30P140 U45 ( .A1(n94), .A2(i_data_bus[62]), .ZN(n52) );
  ND2D1BWP30P140 U46 ( .A1(n94), .A2(i_data_bus[63]), .ZN(n54) );
  CKND2D2BWP30P140 U47 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n21) );
  ND2D1BWP30P140 U48 ( .A1(n94), .A2(i_data_bus[33]), .ZN(n66) );
  ND2D1BWP30P140 U49 ( .A1(n94), .A2(i_data_bus[34]), .ZN(n68) );
  ND2D1BWP30P140 U50 ( .A1(n94), .A2(i_data_bus[35]), .ZN(n43) );
  ND2D1BWP30P140 U51 ( .A1(n94), .A2(i_data_bus[36]), .ZN(n72) );
  ND2D1BWP30P140 U52 ( .A1(n94), .A2(i_data_bus[37]), .ZN(n29) );
  ND2D1BWP30P140 U53 ( .A1(n94), .A2(i_data_bus[38]), .ZN(n27) );
  ND2D1BWP30P140 U54 ( .A1(n94), .A2(i_data_bus[39]), .ZN(n39) );
  INVD1BWP30P140 U55 ( .I(rst), .ZN(n4) );
  ND2D1BWP30P140 U56 ( .A1(n4), .A2(i_en), .ZN(n84) );
  INVD2BWP30P140 U57 ( .I(i_valid[1]), .ZN(n83) );
  MUX2NOPTD4BWP30P140 U58 ( .I0(n83), .I1(n17), .S(n15), .ZN(n5) );
  INVD4BWP30P140 U59 ( .I(n97), .ZN(n105) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[61]), .ZN(n7) );
  INVD1BWP30P140 U61 ( .I(n84), .ZN(n22) );
  INVD2BWP30P140 U62 ( .I(i_cmd[0]), .ZN(n82) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[29]), .ZN(n50) );
  OAI22OPTPBD1BWP30P140 U64 ( .A1(n105), .A2(n7), .B1(n98), .B2(n50), .ZN(N316) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[62]), .ZN(n8) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[30]), .ZN(n53) );
  OAI22OPTPBD1BWP30P140 U67 ( .A1(n105), .A2(n8), .B1(n98), .B2(n53), .ZN(N317) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[63]), .ZN(n9) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[31]), .ZN(n55) );
  OAI22OPTPBD1BWP30P140 U70 ( .A1(n105), .A2(n9), .B1(n98), .B2(n55), .ZN(N318) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[36]), .ZN(n10) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[4]), .ZN(n73) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[37]), .ZN(n11) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[5]), .ZN(n30) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[38]), .ZN(n12) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[6]), .ZN(n28) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[35]), .ZN(n13) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[3]), .ZN(n44) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[39]), .ZN(n14) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[7]), .ZN(n40) );
  INVD2BWP30P140 U81 ( .I(n15), .ZN(n79) );
  NR2OPTPAD2BWP30P140 U82 ( .A1(n79), .A2(n84), .ZN(n19) );
  INVD2BWP30P140 U83 ( .I(i_valid[1]), .ZN(n16) );
  MUX2NOPTD2BWP30P140 U84 ( .I0(n17), .I1(n16), .S(i_cmd[0]), .ZN(n18) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[25]), .ZN(n25) );
  INVD2BWP30P140 U86 ( .I(n21), .ZN(n23) );
  ND2OPTPAD4BWP30P140 U87 ( .A1(n23), .A2(n22), .ZN(n80) );
  OAI21D1BWP30P140 U88 ( .A1(n91), .A2(n25), .B(n24), .ZN(N344) );
  OAI21D1BWP30P140 U89 ( .A1(n95), .A2(n28), .B(n27), .ZN(N325) );
  OAI21D1BWP30P140 U90 ( .A1(n95), .A2(n30), .B(n29), .ZN(N324) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[8]), .ZN(n32) );
  OAI21D1BWP30P140 U92 ( .A1(n95), .A2(n32), .B(n31), .ZN(N327) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[26]), .ZN(n34) );
  OAI21D1BWP30P140 U94 ( .A1(n91), .A2(n34), .B(n33), .ZN(N345) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[10]), .ZN(n36) );
  OAI21D1BWP30P140 U96 ( .A1(n95), .A2(n36), .B(n35), .ZN(N329) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[27]), .ZN(n38) );
  OAI21D1BWP30P140 U98 ( .A1(n91), .A2(n38), .B(n37), .ZN(N346) );
  OAI21D1BWP30P140 U99 ( .A1(n95), .A2(n40), .B(n39), .ZN(N326) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[13]), .ZN(n42) );
  OAI21D1BWP30P140 U101 ( .A1(n91), .A2(n42), .B(n41), .ZN(N332) );
  OAI21D1BWP30P140 U102 ( .A1(n95), .A2(n44), .B(n43), .ZN(N322) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[28]), .ZN(n46) );
  OAI21D1BWP30P140 U104 ( .A1(n91), .A2(n46), .B(n45), .ZN(N347) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[16]), .ZN(n48) );
  OAI21D1BWP30P140 U106 ( .A1(n95), .A2(n48), .B(n47), .ZN(N335) );
  OAI21D1BWP30P140 U107 ( .A1(n91), .A2(n50), .B(n49), .ZN(N348) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[18]), .ZN(n87) );
  OAI21D1BWP30P140 U109 ( .A1(n95), .A2(n87), .B(n51), .ZN(N337) );
  OAI21D1BWP30P140 U110 ( .A1(n91), .A2(n53), .B(n52), .ZN(N349) );
  OAI21D1BWP30P140 U111 ( .A1(n91), .A2(n55), .B(n54), .ZN(N350) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[21]), .ZN(n57) );
  ND2D1BWP30P140 U113 ( .A1(n94), .A2(i_data_bus[53]), .ZN(n56) );
  OAI21D1BWP30P140 U114 ( .A1(n91), .A2(n57), .B(n56), .ZN(N340) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[22]), .ZN(n59) );
  OAI21D1BWP30P140 U116 ( .A1(n91), .A2(n59), .B(n58), .ZN(N341) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[15]), .ZN(n61) );
  OAI21D1BWP30P140 U118 ( .A1(n91), .A2(n61), .B(n60), .ZN(N334) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[23]), .ZN(n63) );
  OAI21D1BWP30P140 U120 ( .A1(n91), .A2(n63), .B(n62), .ZN(N342) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[14]), .ZN(n65) );
  OAI21D1BWP30P140 U122 ( .A1(n95), .A2(n65), .B(n64), .ZN(N333) );
  INVD1BWP30P140 U123 ( .I(i_data_bus[1]), .ZN(n67) );
  OAI21D1BWP30P140 U124 ( .A1(n95), .A2(n67), .B(n66), .ZN(N320) );
  INVD1BWP30P140 U125 ( .I(i_data_bus[2]), .ZN(n69) );
  OAI21D1BWP30P140 U126 ( .A1(n95), .A2(n69), .B(n68), .ZN(N321) );
  INVD1BWP30P140 U127 ( .I(i_data_bus[24]), .ZN(n71) );
  OAI21D1BWP30P140 U128 ( .A1(n95), .A2(n73), .B(n72), .ZN(N323) );
  INVD1BWP30P140 U129 ( .I(i_data_bus[12]), .ZN(n75) );
  INVD1BWP30P140 U130 ( .I(i_data_bus[17]), .ZN(n93) );
  INVD1BWP30P140 U131 ( .I(n78), .ZN(n81) );
  OAI21D1BWP30P140 U132 ( .A1(n81), .A2(n79), .B(n80), .ZN(N354) );
  OAI31D1BWP30P140 U133 ( .A1(n84), .A2(n83), .A3(n82), .B(n98), .ZN(N353) );
  INVD1BWP30P140 U134 ( .I(i_data_bus[19]), .ZN(n90) );
  INVD1BWP30P140 U135 ( .I(i_data_bus[51]), .ZN(n85) );
  OAI22D1BWP30P140 U136 ( .A1(n98), .A2(n90), .B1(n123), .B2(n85), .ZN(N306)
         );
  INVD1BWP30P140 U137 ( .I(i_data_bus[50]), .ZN(n86) );
  OAI22D1BWP30P140 U138 ( .A1(n98), .A2(n87), .B1(n123), .B2(n86), .ZN(N305)
         );
  INVD1BWP30P140 U139 ( .I(i_data_bus[9]), .ZN(n88) );
  MOAI22D1BWP30P140 U140 ( .A1(n88), .A2(n91), .B1(i_data_bus[41]), .B2(n94), 
        .ZN(N328) );
  INVD1BWP30P140 U141 ( .I(i_data_bus[20]), .ZN(n89) );
  MOAI22D1BWP30P140 U142 ( .A1(n89), .A2(n95), .B1(i_data_bus[52]), .B2(n94), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U143 ( .A1(n90), .A2(n91), .B1(i_data_bus[51]), .B2(n94), 
        .ZN(N338) );
  INVD1BWP30P140 U144 ( .I(i_data_bus[11]), .ZN(n92) );
  MOAI22D1BWP30P140 U145 ( .A1(n92), .A2(n91), .B1(i_data_bus[43]), .B2(n94), 
        .ZN(N330) );
  MOAI22D1BWP30P140 U146 ( .A1(n93), .A2(n95), .B1(i_data_bus[49]), .B2(n94), 
        .ZN(N336) );
  INVD1BWP30P140 U147 ( .I(i_data_bus[0]), .ZN(n96) );
  MOAI22D1BWP30P140 U148 ( .A1(n96), .A2(n91), .B1(i_data_bus[32]), .B2(n94), 
        .ZN(N319) );
  INVD4BWP30P140 U149 ( .I(n97), .ZN(n120) );
  INVD1BWP30P140 U150 ( .I(i_data_bus[60]), .ZN(n99) );
  MOAI22D1BWP30P140 U151 ( .A1(n120), .A2(n99), .B1(n121), .B2(i_data_bus[28]), 
        .ZN(N315) );
  INVD1BWP30P140 U152 ( .I(i_data_bus[48]), .ZN(n100) );
  MOAI22D1BWP30P140 U153 ( .A1(n1), .A2(n100), .B1(n121), .B2(i_data_bus[16]), 
        .ZN(N303) );
  INVD1BWP30P140 U154 ( .I(i_data_bus[34]), .ZN(n101) );
  MOAI22D1BWP30P140 U155 ( .A1(n120), .A2(n101), .B1(n121), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140 U156 ( .I(i_data_bus[59]), .ZN(n102) );
  MOAI22D1BWP30P140 U157 ( .A1(n120), .A2(n102), .B1(n121), .B2(i_data_bus[27]), .ZN(N314) );
  INVD1BWP30P140 U158 ( .I(i_data_bus[47]), .ZN(n103) );
  MOAI22D1BWP30P140 U159 ( .A1(n1), .A2(n103), .B1(n121), .B2(i_data_bus[15]), 
        .ZN(N302) );
  INVD1BWP30P140 U160 ( .I(i_data_bus[33]), .ZN(n104) );
  MOAI22D1BWP30P140 U161 ( .A1(n105), .A2(n104), .B1(n121), .B2(i_data_bus[1]), 
        .ZN(N288) );
  INVD1BWP30P140 U162 ( .I(i_data_bus[58]), .ZN(n106) );
  MOAI22D1BWP30P140 U163 ( .A1(n120), .A2(n106), .B1(n121), .B2(i_data_bus[26]), .ZN(N313) );
  INVD1BWP30P140 U164 ( .I(i_data_bus[46]), .ZN(n107) );
  MOAI22D1BWP30P140 U165 ( .A1(n1), .A2(n107), .B1(n121), .B2(i_data_bus[14]), 
        .ZN(N301) );
  INVD1BWP30P140 U166 ( .I(i_data_bus[32]), .ZN(n108) );
  MOAI22D1BWP30P140 U167 ( .A1(n120), .A2(n108), .B1(n121), .B2(i_data_bus[0]), 
        .ZN(N287) );
  INVD1BWP30P140 U168 ( .I(i_data_bus[57]), .ZN(n109) );
  MOAI22D1BWP30P140 U169 ( .A1(n120), .A2(n109), .B1(n121), .B2(i_data_bus[25]), .ZN(N312) );
  INVD1BWP30P140 U170 ( .I(i_data_bus[45]), .ZN(n110) );
  MOAI22D1BWP30P140 U171 ( .A1(n1), .A2(n110), .B1(n121), .B2(i_data_bus[13]), 
        .ZN(N300) );
  INVD1BWP30P140 U172 ( .I(i_data_bus[56]), .ZN(n111) );
  MOAI22D1BWP30P140 U173 ( .A1(n120), .A2(n111), .B1(n121), .B2(i_data_bus[24]), .ZN(N311) );
  INVD1BWP30P140 U174 ( .I(i_data_bus[44]), .ZN(n112) );
  MOAI22D1BWP30P140 U175 ( .A1(n1), .A2(n112), .B1(n121), .B2(i_data_bus[12]), 
        .ZN(N299) );
  INVD1BWP30P140 U176 ( .I(i_data_bus[55]), .ZN(n113) );
  MOAI22D1BWP30P140 U177 ( .A1(n120), .A2(n113), .B1(n121), .B2(i_data_bus[23]), .ZN(N310) );
  INVD1BWP30P140 U178 ( .I(i_data_bus[43]), .ZN(n114) );
  MOAI22D1BWP30P140 U179 ( .A1(n1), .A2(n114), .B1(n121), .B2(i_data_bus[11]), 
        .ZN(N298) );
  INVD1BWP30P140 U180 ( .I(i_data_bus[54]), .ZN(n115) );
  MOAI22D1BWP30P140 U181 ( .A1(n120), .A2(n115), .B1(n121), .B2(i_data_bus[22]), .ZN(N309) );
  INVD1BWP30P140 U182 ( .I(i_data_bus[42]), .ZN(n116) );
  MOAI22D1BWP30P140 U183 ( .A1(n1), .A2(n116), .B1(n121), .B2(i_data_bus[10]), 
        .ZN(N297) );
  INVD1BWP30P140 U184 ( .I(i_data_bus[53]), .ZN(n117) );
  MOAI22D1BWP30P140 U185 ( .A1(n120), .A2(n117), .B1(n121), .B2(i_data_bus[21]), .ZN(N308) );
  INVD1BWP30P140 U186 ( .I(i_data_bus[41]), .ZN(n118) );
  MOAI22D1BWP30P140 U187 ( .A1(n1), .A2(n118), .B1(n121), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140 U188 ( .I(i_data_bus[52]), .ZN(n119) );
  MOAI22D1BWP30P140 U189 ( .A1(n120), .A2(n119), .B1(n121), .B2(i_data_bus[20]), .ZN(N307) );
  INVD1BWP30P140 U190 ( .I(i_data_bus[40]), .ZN(n122) );
  MOAI22D1BWP30P140 U191 ( .A1(n1), .A2(n122), .B1(n121), .B2(i_data_bus[8]), 
        .ZN(N295) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_132 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n110), .A2(n33), .B1(n101), .B2(n32), .ZN(N317) );
  OAI22D1BWP30P140 U4 ( .A1(n110), .A2(n36), .B1(n101), .B2(n51), .ZN(N291) );
  OAI22D1BWP30P140 U5 ( .A1(n110), .A2(n39), .B1(n101), .B2(n38), .ZN(N294) );
  OAI21D2BWP30P140 U6 ( .A1(n86), .A2(n38), .B(n23), .ZN(N326) );
  OAI22D1BWP30P140 U7 ( .A1(n110), .A2(n40), .B1(n101), .B2(n55), .ZN(N293) );
  OAI21D2BWP30P140 U8 ( .A1(n86), .A2(n30), .B(n24), .ZN(N350) );
  OAI22D1BWP30P140 U9 ( .A1(n110), .A2(n41), .B1(n101), .B2(n53), .ZN(N292) );
  CKND2D3BWP30P140 U10 ( .A1(n83), .A2(i_data_bus[47]), .ZN(n70) );
  CKND2D3BWP30P140 U11 ( .A1(n83), .A2(i_data_bus[49]), .ZN(n74) );
  CKND2D3BWP30P140 U12 ( .A1(n83), .A2(i_data_bus[50]), .ZN(n75) );
  CKND2D3BWP30P140 U13 ( .A1(n83), .A2(i_data_bus[48]), .ZN(n72) );
  CKND2D3BWP30P140 U14 ( .A1(n83), .A2(i_data_bus[51]), .ZN(n76) );
  CKND2D3BWP30P140 U15 ( .A1(n83), .A2(i_data_bus[52]), .ZN(n77) );
  CKND2D3BWP30P140 U16 ( .A1(n83), .A2(i_data_bus[53]), .ZN(n79) );
  CKND2D3BWP30P140 U17 ( .A1(n83), .A2(i_data_bus[54]), .ZN(n81) );
  INVD9BWP30P140 U18 ( .I(n101), .ZN(n125) );
  INVD3BWP30P140 U19 ( .I(n3), .ZN(n90) );
  INVD2BWP30P140 U20 ( .I(i_valid[1]), .ZN(n5) );
  ND2OPTPAD6BWP30P140 U21 ( .A1(n28), .A2(n27), .ZN(n103) );
  INVD6BWP30P140 U22 ( .I(n103), .ZN(n100) );
  INVD3BWP30P140 U23 ( .I(n9), .ZN(n10) );
  OAI21D2BWP30P140 U24 ( .A1(n86), .A2(n87), .B(n76), .ZN(N338) );
  OAI21D2BWP30P140 U25 ( .A1(n86), .A2(n78), .B(n77), .ZN(N339) );
  OAI21D2BWP30P140 U26 ( .A1(n86), .A2(n80), .B(n79), .ZN(N340) );
  OAI21D2BWP30P140 U27 ( .A1(n86), .A2(n82), .B(n81), .ZN(N341) );
  OAI21D2BWP30P140 U28 ( .A1(n86), .A2(n12), .B(n11), .ZN(N343) );
  OAI21D2BWP30P140 U29 ( .A1(n86), .A2(n14), .B(n13), .ZN(N344) );
  OAI21D2BWP30P140 U30 ( .A1(n86), .A2(n16), .B(n15), .ZN(N345) );
  OAI21D2BWP30P140 U31 ( .A1(n86), .A2(n18), .B(n17), .ZN(N346) );
  OAI21D2BWP30P140 U32 ( .A1(n1), .A2(n43), .B(n42), .ZN(N319) );
  INVD6BWP30P140 U33 ( .I(n2), .ZN(n8) );
  INVD15BWP30P140 U34 ( .I(n8), .ZN(n86) );
  OAI22D1BWP30P140 U35 ( .A1(n110), .A2(n37), .B1(n101), .B2(n49), .ZN(N290)
         );
  OAI22D1BWP30P140 U36 ( .A1(n110), .A2(n35), .B1(n101), .B2(n34), .ZN(N316)
         );
  ND2OPTPAD6BWP30P140 U37 ( .A1(n90), .A2(n93), .ZN(n101) );
  OAI21OPTREPBD2BWP30P140 U38 ( .A1(n86), .A2(n34), .B(n21), .ZN(N348) );
  OAI21OPTREPBD2BWP30P140 U39 ( .A1(n86), .A2(n32), .B(n22), .ZN(N349) );
  NR2OPTPAD1BWP30P140 U40 ( .A1(i_cmd[1]), .A2(n95), .ZN(n7) );
  INVD4BWP30P140 U41 ( .I(i_cmd[1]), .ZN(n25) );
  CKBD1BWP30P140 U42 ( .I(n2), .Z(n1) );
  CKND2D3BWP30P140 U43 ( .A1(i_valid[1]), .A2(i_cmd[1]), .ZN(n9) );
  OAI21OPTREPBD2BWP30P140 U44 ( .A1(n86), .A2(n85), .B(n84), .ZN(N342) );
  OAI21OPTREPBD2BWP30P140 U45 ( .A1(n86), .A2(n20), .B(n19), .ZN(N347) );
  OAI21D2BWP30P140 U46 ( .A1(n86), .A2(n45), .B(n44), .ZN(N320) );
  OAI21D2BWP30P140 U47 ( .A1(n86), .A2(n47), .B(n46), .ZN(N321) );
  OAI21D2BWP30P140 U48 ( .A1(n86), .A2(n49), .B(n48), .ZN(N322) );
  OAI21D2BWP30P140 U49 ( .A1(n86), .A2(n51), .B(n50), .ZN(N323) );
  OAI21D2BWP30P140 U50 ( .A1(n86), .A2(n53), .B(n52), .ZN(N324) );
  OAI21D2BWP30P140 U51 ( .A1(n86), .A2(n55), .B(n54), .ZN(N325) );
  OAI21D2BWP30P140 U52 ( .A1(n86), .A2(n57), .B(n56), .ZN(N327) );
  OAI21D2BWP30P140 U53 ( .A1(n86), .A2(n59), .B(n58), .ZN(N328) );
  OAI21D2BWP30P140 U54 ( .A1(n86), .A2(n61), .B(n60), .ZN(N329) );
  OAI21D2BWP30P140 U55 ( .A1(n86), .A2(n63), .B(n62), .ZN(N330) );
  OAI21D2BWP30P140 U56 ( .A1(n1), .A2(n65), .B(n64), .ZN(N331) );
  OAI21D2BWP30P140 U57 ( .A1(n86), .A2(n67), .B(n66), .ZN(N332) );
  OAI21D2BWP30P140 U58 ( .A1(n86), .A2(n69), .B(n68), .ZN(N333) );
  OAI21D2BWP30P140 U59 ( .A1(n86), .A2(n71), .B(n70), .ZN(N334) );
  OAI21D2BWP30P140 U60 ( .A1(n86), .A2(n73), .B(n72), .ZN(N335) );
  OAI21D2BWP30P140 U61 ( .A1(n86), .A2(n97), .B(n74), .ZN(N336) );
  OAI21D2BWP30P140 U62 ( .A1(n86), .A2(n99), .B(n75), .ZN(N337) );
  CKND2D4BWP30P140 U63 ( .A1(n6), .A2(n7), .ZN(n2) );
  CKND2D3BWP30P140 U64 ( .A1(i_valid[0]), .A2(n29), .ZN(n3) );
  MUX2NOPTD4BWP30P140 U65 ( .I0(n26), .I1(n5), .S(i_cmd[0]), .ZN(n6) );
  ND2D1BWP30P140 U66 ( .A1(n89), .A2(n88), .ZN(N306) );
  OR2D1BWP30P140 U67 ( .A1(n101), .A2(n87), .Z(n88) );
  ND2OPTIBD1BWP30P140 U68 ( .A1(n100), .A2(i_data_bus[51]), .ZN(n89) );
  CKND2D2BWP30P140 U69 ( .A1(n83), .A2(i_data_bus[55]), .ZN(n84) );
  CKND2D2BWP30P140 U70 ( .A1(n83), .A2(i_data_bus[60]), .ZN(n19) );
  CKND2D2BWP30P140 U71 ( .A1(n83), .A2(i_data_bus[61]), .ZN(n21) );
  CKND2D2BWP30P140 U72 ( .A1(n83), .A2(i_data_bus[62]), .ZN(n22) );
  INVD1BWP30P140 U73 ( .I(rst), .ZN(n4) );
  ND2D1BWP30P140 U74 ( .A1(n4), .A2(i_en), .ZN(n95) );
  INVD3BWP30P140 U75 ( .I(i_valid[0]), .ZN(n26) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[24]), .ZN(n12) );
  INVD1BWP30P140 U77 ( .I(n95), .ZN(n29) );
  ND2OPTPAD6BWP30P140 U78 ( .A1(n10), .A2(n29), .ZN(n91) );
  INVD15BWP30P140 U79 ( .I(n91), .ZN(n83) );
  ND2OPTIBD4BWP30P140 U80 ( .A1(n83), .A2(i_data_bus[56]), .ZN(n11) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[25]), .ZN(n14) );
  ND2OPTIBD4BWP30P140 U82 ( .A1(n83), .A2(i_data_bus[57]), .ZN(n13) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[26]), .ZN(n16) );
  ND2OPTIBD4BWP30P140 U84 ( .A1(n83), .A2(i_data_bus[58]), .ZN(n15) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[27]), .ZN(n18) );
  ND2OPTIBD4BWP30P140 U86 ( .A1(n83), .A2(i_data_bus[59]), .ZN(n17) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[28]), .ZN(n20) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[29]), .ZN(n34) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[30]), .ZN(n32) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[7]), .ZN(n38) );
  CKND2D3BWP30P140 U91 ( .A1(n83), .A2(i_data_bus[39]), .ZN(n23) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[31]), .ZN(n30) );
  CKND2D3BWP30P140 U93 ( .A1(n83), .A2(i_data_bus[63]), .ZN(n24) );
  INR2D4BWP30P140 U94 ( .A1(i_cmd[0]), .B1(n95), .ZN(n28) );
  INVD2BWP30P140 U95 ( .I(i_valid[1]), .ZN(n94) );
  MUX2NOPTD4BWP30P140 U96 ( .I0(n94), .I1(n26), .S(n25), .ZN(n27) );
  INVD4BWP30P140 U97 ( .I(n100), .ZN(n110) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[63]), .ZN(n31) );
  INVD3BWP30P140 U99 ( .I(i_cmd[0]), .ZN(n93) );
  OAI22OPTPBD1BWP30P140 U100 ( .A1(n110), .A2(n31), .B1(n101), .B2(n30), .ZN(
        N318) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[62]), .ZN(n33) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[61]), .ZN(n35) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[36]), .ZN(n36) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[4]), .ZN(n51) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[35]), .ZN(n37) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[3]), .ZN(n49) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[39]), .ZN(n39) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[38]), .ZN(n40) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[6]), .ZN(n55) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[37]), .ZN(n41) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[5]), .ZN(n53) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[0]), .ZN(n43) );
  ND2OPTIBD4BWP30P140 U113 ( .A1(n83), .A2(i_data_bus[32]), .ZN(n42) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[1]), .ZN(n45) );
  ND2OPTIBD4BWP30P140 U115 ( .A1(n83), .A2(i_data_bus[33]), .ZN(n44) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[2]), .ZN(n47) );
  ND2OPTIBD4BWP30P140 U117 ( .A1(n83), .A2(i_data_bus[34]), .ZN(n46) );
  ND2OPTIBD4BWP30P140 U118 ( .A1(n83), .A2(i_data_bus[35]), .ZN(n48) );
  ND2OPTIBD4BWP30P140 U119 ( .A1(n83), .A2(i_data_bus[36]), .ZN(n50) );
  ND2OPTIBD4BWP30P140 U120 ( .A1(n83), .A2(i_data_bus[37]), .ZN(n52) );
  ND2OPTIBD4BWP30P140 U121 ( .A1(n83), .A2(i_data_bus[38]), .ZN(n54) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[8]), .ZN(n57) );
  ND2OPTIBD4BWP30P140 U123 ( .A1(n83), .A2(i_data_bus[40]), .ZN(n56) );
  INVD1BWP30P140 U124 ( .I(i_data_bus[9]), .ZN(n59) );
  ND2OPTIBD4BWP30P140 U125 ( .A1(n83), .A2(i_data_bus[41]), .ZN(n58) );
  INVD1BWP30P140 U126 ( .I(i_data_bus[10]), .ZN(n61) );
  ND2OPTIBD4BWP30P140 U127 ( .A1(n83), .A2(i_data_bus[42]), .ZN(n60) );
  INVD1BWP30P140 U128 ( .I(i_data_bus[11]), .ZN(n63) );
  ND2OPTIBD4BWP30P140 U129 ( .A1(n83), .A2(i_data_bus[43]), .ZN(n62) );
  INVD1BWP30P140 U130 ( .I(i_data_bus[12]), .ZN(n65) );
  ND2OPTIBD4BWP30P140 U131 ( .A1(n83), .A2(i_data_bus[44]), .ZN(n64) );
  INVD1BWP30P140 U132 ( .I(i_data_bus[13]), .ZN(n67) );
  ND2OPTIBD4BWP30P140 U133 ( .A1(n83), .A2(i_data_bus[45]), .ZN(n66) );
  INVD1BWP30P140 U134 ( .I(i_data_bus[14]), .ZN(n69) );
  ND2OPTIBD4BWP30P140 U135 ( .A1(n83), .A2(i_data_bus[46]), .ZN(n68) );
  INVD1BWP30P140 U136 ( .I(i_data_bus[15]), .ZN(n71) );
  INVD1BWP30P140 U137 ( .I(i_data_bus[16]), .ZN(n73) );
  INVD1BWP30P140 U138 ( .I(i_data_bus[17]), .ZN(n97) );
  INVD1BWP30P140 U139 ( .I(i_data_bus[18]), .ZN(n99) );
  INVD1BWP30P140 U140 ( .I(i_data_bus[19]), .ZN(n87) );
  INVD1BWP30P140 U141 ( .I(i_data_bus[20]), .ZN(n78) );
  INVD1BWP30P140 U142 ( .I(i_data_bus[21]), .ZN(n80) );
  INVD1BWP30P140 U143 ( .I(i_data_bus[22]), .ZN(n82) );
  INVD1BWP30P140 U144 ( .I(i_data_bus[23]), .ZN(n85) );
  INVD1BWP30P140 U145 ( .I(n90), .ZN(n92) );
  OAI21D1BWP30P140 U146 ( .A1(n92), .A2(i_cmd[1]), .B(n91), .ZN(N354) );
  OAI31D1BWP30P140 U147 ( .A1(n95), .A2(n94), .A3(n93), .B(n101), .ZN(N353) );
  INVD1BWP30P140 U148 ( .I(i_data_bus[49]), .ZN(n96) );
  OAI22D1BWP30P140 U149 ( .A1(n101), .A2(n97), .B1(n103), .B2(n96), .ZN(N304)
         );
  INVD1BWP30P140 U150 ( .I(i_data_bus[50]), .ZN(n98) );
  OAI22D1BWP30P140 U151 ( .A1(n101), .A2(n99), .B1(n103), .B2(n98), .ZN(N305)
         );
  INVD4BWP30P140 U152 ( .I(n100), .ZN(n124) );
  INVD1BWP30P140 U153 ( .I(i_data_bus[60]), .ZN(n102) );
  MOAI22D1BWP30P140 U154 ( .A1(n124), .A2(n102), .B1(n125), .B2(i_data_bus[28]), .ZN(N315) );
  BUFFD4BWP30P140 U155 ( .I(n103), .Z(n127) );
  INVD1BWP30P140 U156 ( .I(i_data_bus[48]), .ZN(n104) );
  MOAI22D1BWP30P140 U157 ( .A1(n127), .A2(n104), .B1(n125), .B2(i_data_bus[16]), .ZN(N303) );
  INVD1BWP30P140 U158 ( .I(i_data_bus[34]), .ZN(n105) );
  MOAI22D1BWP30P140 U159 ( .A1(n124), .A2(n105), .B1(n125), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140 U160 ( .I(i_data_bus[59]), .ZN(n106) );
  MOAI22D1BWP30P140 U161 ( .A1(n124), .A2(n106), .B1(n125), .B2(i_data_bus[27]), .ZN(N314) );
  INVD1BWP30P140 U162 ( .I(i_data_bus[47]), .ZN(n107) );
  MOAI22D1BWP30P140 U163 ( .A1(n127), .A2(n107), .B1(n125), .B2(i_data_bus[15]), .ZN(N302) );
  INVD1BWP30P140 U164 ( .I(i_data_bus[33]), .ZN(n108) );
  MOAI22D1BWP30P140 U165 ( .A1(n124), .A2(n108), .B1(n125), .B2(i_data_bus[1]), 
        .ZN(N288) );
  INVD1BWP30P140 U166 ( .I(i_data_bus[58]), .ZN(n109) );
  MOAI22D1BWP30P140 U167 ( .A1(n110), .A2(n109), .B1(n125), .B2(i_data_bus[26]), .ZN(N313) );
  INVD1BWP30P140 U168 ( .I(i_data_bus[46]), .ZN(n111) );
  MOAI22D1BWP30P140 U169 ( .A1(n127), .A2(n111), .B1(n125), .B2(i_data_bus[14]), .ZN(N301) );
  INVD1BWP30P140 U170 ( .I(i_data_bus[32]), .ZN(n112) );
  MOAI22D1BWP30P140 U171 ( .A1(n124), .A2(n112), .B1(n125), .B2(i_data_bus[0]), 
        .ZN(N287) );
  INVD1BWP30P140 U172 ( .I(i_data_bus[57]), .ZN(n113) );
  MOAI22D1BWP30P140 U173 ( .A1(n124), .A2(n113), .B1(n125), .B2(i_data_bus[25]), .ZN(N312) );
  INVD1BWP30P140 U174 ( .I(i_data_bus[45]), .ZN(n114) );
  MOAI22D1BWP30P140 U175 ( .A1(n127), .A2(n114), .B1(n125), .B2(i_data_bus[13]), .ZN(N300) );
  INVD1BWP30P140 U176 ( .I(i_data_bus[56]), .ZN(n115) );
  MOAI22D1BWP30P140 U177 ( .A1(n124), .A2(n115), .B1(n125), .B2(i_data_bus[24]), .ZN(N311) );
  INVD1BWP30P140 U178 ( .I(i_data_bus[44]), .ZN(n116) );
  MOAI22D1BWP30P140 U179 ( .A1(n127), .A2(n116), .B1(n125), .B2(i_data_bus[12]), .ZN(N299) );
  INVD1BWP30P140 U180 ( .I(i_data_bus[55]), .ZN(n117) );
  MOAI22D1BWP30P140 U181 ( .A1(n124), .A2(n117), .B1(n125), .B2(i_data_bus[23]), .ZN(N310) );
  INVD1BWP30P140 U182 ( .I(i_data_bus[43]), .ZN(n118) );
  MOAI22D1BWP30P140 U183 ( .A1(n127), .A2(n118), .B1(n125), .B2(i_data_bus[11]), .ZN(N298) );
  INVD1BWP30P140 U184 ( .I(i_data_bus[54]), .ZN(n119) );
  MOAI22D1BWP30P140 U185 ( .A1(n124), .A2(n119), .B1(n125), .B2(i_data_bus[22]), .ZN(N309) );
  INVD1BWP30P140 U186 ( .I(i_data_bus[42]), .ZN(n120) );
  MOAI22D1BWP30P140 U187 ( .A1(n127), .A2(n120), .B1(n125), .B2(i_data_bus[10]), .ZN(N297) );
  INVD1BWP30P140 U188 ( .I(i_data_bus[53]), .ZN(n121) );
  MOAI22D1BWP30P140 U189 ( .A1(n124), .A2(n121), .B1(n125), .B2(i_data_bus[21]), .ZN(N308) );
  INVD1BWP30P140 U190 ( .I(i_data_bus[41]), .ZN(n122) );
  MOAI22D1BWP30P140 U191 ( .A1(n127), .A2(n122), .B1(n125), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140 U192 ( .I(i_data_bus[52]), .ZN(n123) );
  MOAI22D1BWP30P140 U193 ( .A1(n124), .A2(n123), .B1(n125), .B2(i_data_bus[20]), .ZN(N307) );
  INVD1BWP30P140 U194 ( .I(i_data_bus[40]), .ZN(n126) );
  MOAI22D1BWP30P140 U195 ( .A1(n127), .A2(n126), .B1(n125), .B2(i_data_bus[8]), 
        .ZN(N295) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_133 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI21D1P5BWP30P140 U3 ( .A1(n5), .A2(n101), .B(n30), .ZN(N336) );
  OAI21D1P5BWP30P140 U4 ( .A1(n5), .A2(n34), .B(n33), .ZN(N331) );
  OAI21D1P5BWP30P140 U5 ( .A1(n57), .A2(n36), .B(n35), .ZN(N329) );
  OAI21D1P5BWP30P140 U6 ( .A1(n5), .A2(n38), .B(n37), .ZN(N328) );
  OAI21D1P5BWP30P140 U7 ( .A1(n57), .A2(n40), .B(n39), .ZN(N327) );
  OAI21D1P5BWP30P140 U8 ( .A1(n5), .A2(n52), .B(n51), .ZN(N321) );
  OAI21D1P5BWP30P140 U9 ( .A1(n89), .A2(n26), .B(n25), .ZN(N346) );
  OAI21D1P5BWP30P140 U10 ( .A1(n57), .A2(n56), .B(n55), .ZN(N319) );
  CKND2D2BWP30P140 U11 ( .A1(n86), .A2(i_data_bus[58]), .ZN(n68) );
  CKND2D2BWP30P140 U12 ( .A1(n86), .A2(i_data_bus[54]), .ZN(n70) );
  CKND2D3BWP30P140 U13 ( .A1(n86), .A2(i_data_bus[63]), .ZN(n72) );
  CKND2D3BWP30P140 U14 ( .A1(n86), .A2(i_data_bus[53]), .ZN(n76) );
  CKND2D3BWP30P140 U15 ( .A1(n86), .A2(i_data_bus[56]), .ZN(n78) );
  CKND2D3BWP30P140 U16 ( .A1(n86), .A2(i_data_bus[55]), .ZN(n80) );
  CKND2D3BWP30P140 U17 ( .A1(n86), .A2(i_data_bus[61]), .ZN(n87) );
  CKND2D3BWP30P140 U18 ( .A1(n86), .A2(i_data_bus[57]), .ZN(n82) );
  ND2OPTPAD6BWP30P140 U19 ( .A1(n93), .A2(n97), .ZN(n105) );
  INVD12BWP30P140 U20 ( .I(n95), .ZN(n86) );
  CKND2D4BWP30P140 U21 ( .A1(n8), .A2(n7), .ZN(n126) );
  INVD8BWP30P140 U22 ( .I(n22), .ZN(n27) );
  CKND2D3BWP30P140 U23 ( .A1(i_valid[0]), .A2(n23), .ZN(n3) );
  INVD8BWP30P140 U24 ( .I(n105), .ZN(n128) );
  OAI21D2BWP30P140 U25 ( .A1(n57), .A2(n77), .B(n76), .ZN(N340) );
  OAI21D2BWP30P140 U26 ( .A1(n5), .A2(n54), .B(n53), .ZN(N320) );
  OAI21D2BWP30P140 U27 ( .A1(n89), .A2(n69), .B(n68), .ZN(N345) );
  BUFFD4BWP30P140 U28 ( .I(n126), .Z(n1) );
  OAI21D2BWP30P140 U29 ( .A1(n89), .A2(n71), .B(n70), .ZN(N341) );
  OAI21D2BWP30P140 U30 ( .A1(n5), .A2(n79), .B(n78), .ZN(N343) );
  OAI21D2BWP30P140 U31 ( .A1(n57), .A2(n83), .B(n82), .ZN(N344) );
  OAI21D2BWP30P140 U32 ( .A1(n89), .A2(n73), .B(n72), .ZN(N350) );
  OAI21D2BWP30P140 U33 ( .A1(n5), .A2(n81), .B(n80), .ZN(N342) );
  INVD2BWP30P140 U34 ( .I(i_valid[1]), .ZN(n18) );
  INVD2BWP30P140 U35 ( .I(n2), .ZN(n24) );
  ND2OPTIBD1BWP30P140 U36 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n2) );
  OAI21OPTREPBD2BWP30P140 U37 ( .A1(n89), .A2(n75), .B(n74), .ZN(N347) );
  OAI21OPTREPBD2BWP30P140 U38 ( .A1(n5), .A2(n85), .B(n84), .ZN(N349) );
  INVD3BWP30P140 U39 ( .I(i_valid[0]), .ZN(n19) );
  INVD3BWP30P140 U40 ( .I(n3), .ZN(n93) );
  INVD4BWP30P140 U41 ( .I(n104), .ZN(n109) );
  INVD1BWP30P140 U42 ( .I(i_cmd[0]), .ZN(n4) );
  NR2OPTPAD1BWP30P140 U43 ( .A1(n4), .A2(n99), .ZN(n8) );
  NR2OPTPAD2BWP30P140 U44 ( .A1(n94), .A2(n99), .ZN(n21) );
  OAI21D2BWP30P140 U45 ( .A1(n57), .A2(n88), .B(n87), .ZN(N348) );
  ND2D1BWP30P140 U46 ( .A1(n92), .A2(n91), .ZN(N305) );
  OR2D1BWP30P140 U47 ( .A1(n105), .A2(n90), .Z(n91) );
  ND2D1BWP30P140 U48 ( .A1(n104), .A2(i_data_bus[50]), .ZN(n92) );
  INVD9BWP30P140 U49 ( .I(n27), .ZN(n5) );
  INVD1BWP30P140 U50 ( .I(rst), .ZN(n6) );
  ND2D1BWP30P140 U51 ( .A1(n6), .A2(i_en), .ZN(n99) );
  INVD2BWP30P140 U52 ( .I(i_valid[1]), .ZN(n98) );
  INVD3BWP30P140 U53 ( .I(i_cmd[1]), .ZN(n17) );
  MUX2NOPTD4BWP30P140 U54 ( .I0(n98), .I1(n19), .S(n17), .ZN(n7) );
  INVD4BWP30P140 U55 ( .I(n126), .ZN(n104) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[61]), .ZN(n9) );
  INVD1BWP30P140 U57 ( .I(n99), .ZN(n23) );
  INVD2BWP30P140 U58 ( .I(i_cmd[0]), .ZN(n97) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[29]), .ZN(n88) );
  OAI22OPTPBD1BWP30P140 U60 ( .A1(n109), .A2(n9), .B1(n105), .B2(n88), .ZN(
        N316) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[63]), .ZN(n10) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[31]), .ZN(n73) );
  OAI22OPTPBD1BWP30P140 U63 ( .A1(n109), .A2(n10), .B1(n105), .B2(n73), .ZN(
        N318) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[62]), .ZN(n11) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[30]), .ZN(n85) );
  OAI22OPTPBD1BWP30P140 U66 ( .A1(n109), .A2(n11), .B1(n105), .B2(n85), .ZN(
        N317) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[39]), .ZN(n12) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[7]), .ZN(n42) );
  OAI22OPTPBD1BWP30P140 U69 ( .A1(n109), .A2(n12), .B1(n105), .B2(n42), .ZN(
        N294) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[38]), .ZN(n13) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[6]), .ZN(n44) );
  OAI22OPTPBD1BWP30P140 U72 ( .A1(n109), .A2(n13), .B1(n105), .B2(n44), .ZN(
        N293) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[37]), .ZN(n14) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[5]), .ZN(n46) );
  OAI22OPTPBD1BWP30P140 U75 ( .A1(n109), .A2(n14), .B1(n105), .B2(n46), .ZN(
        N292) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[36]), .ZN(n15) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[4]), .ZN(n48) );
  OAI22OPTPBD1BWP30P140 U78 ( .A1(n109), .A2(n15), .B1(n105), .B2(n48), .ZN(
        N291) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[35]), .ZN(n16) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[3]), .ZN(n50) );
  OAI22OPTPBD1BWP30P140 U81 ( .A1(n109), .A2(n16), .B1(n105), .B2(n50), .ZN(
        N290) );
  INVD2BWP30P140 U82 ( .I(n17), .ZN(n94) );
  MUX2NOPTD4BWP30P140 U83 ( .I0(n19), .I1(n18), .S(i_cmd[0]), .ZN(n20) );
  ND2OPTPAD4BWP30P140 U84 ( .A1(n21), .A2(n20), .ZN(n22) );
  INVD9BWP30P140 U85 ( .I(n27), .ZN(n89) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[27]), .ZN(n26) );
  ND2OPTPAD6BWP30P140 U87 ( .A1(n24), .A2(n23), .ZN(n95) );
  CKND2D2BWP30P140 U88 ( .A1(n86), .A2(i_data_bus[59]), .ZN(n25) );
  INVD8BWP30P140 U89 ( .I(n27), .ZN(n57) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[19]), .ZN(n103) );
  ND2OPTIBD2BWP30P140 U91 ( .A1(n86), .A2(i_data_bus[51]), .ZN(n28) );
  OAI21OPTREPBD2BWP30P140 U92 ( .A1(n5), .A2(n103), .B(n28), .ZN(N338) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[18]), .ZN(n90) );
  ND2OPTIBD2BWP30P140 U94 ( .A1(n86), .A2(i_data_bus[50]), .ZN(n29) );
  OAI21OPTREPBD2BWP30P140 U95 ( .A1(n57), .A2(n90), .B(n29), .ZN(N337) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[17]), .ZN(n101) );
  ND2OPTIBD2BWP30P140 U97 ( .A1(n86), .A2(i_data_bus[49]), .ZN(n30) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[16]), .ZN(n32) );
  ND2OPTIBD2BWP30P140 U99 ( .A1(n86), .A2(i_data_bus[48]), .ZN(n31) );
  OAI21OPTREPBD2BWP30P140 U100 ( .A1(n57), .A2(n32), .B(n31), .ZN(N335) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[12]), .ZN(n34) );
  ND2OPTIBD2BWP30P140 U102 ( .A1(n86), .A2(i_data_bus[44]), .ZN(n33) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[10]), .ZN(n36) );
  ND2OPTIBD2BWP30P140 U104 ( .A1(n86), .A2(i_data_bus[42]), .ZN(n35) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[9]), .ZN(n38) );
  ND2OPTIBD2BWP30P140 U106 ( .A1(n86), .A2(i_data_bus[41]), .ZN(n37) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[8]), .ZN(n40) );
  ND2OPTIBD2BWP30P140 U108 ( .A1(n86), .A2(i_data_bus[40]), .ZN(n39) );
  ND2OPTIBD2BWP30P140 U109 ( .A1(n86), .A2(i_data_bus[39]), .ZN(n41) );
  OAI21OPTREPBD2BWP30P140 U110 ( .A1(n89), .A2(n42), .B(n41), .ZN(N326) );
  ND2OPTIBD2BWP30P140 U111 ( .A1(n86), .A2(i_data_bus[38]), .ZN(n43) );
  OAI21OPTREPBD2BWP30P140 U112 ( .A1(n5), .A2(n44), .B(n43), .ZN(N325) );
  ND2OPTIBD2BWP30P140 U113 ( .A1(n86), .A2(i_data_bus[37]), .ZN(n45) );
  OAI21OPTREPBD2BWP30P140 U114 ( .A1(n57), .A2(n46), .B(n45), .ZN(N324) );
  ND2OPTIBD2BWP30P140 U115 ( .A1(n86), .A2(i_data_bus[36]), .ZN(n47) );
  OAI21OPTREPBD2BWP30P140 U116 ( .A1(n5), .A2(n48), .B(n47), .ZN(N323) );
  ND2OPTIBD2BWP30P140 U117 ( .A1(n86), .A2(i_data_bus[35]), .ZN(n49) );
  OAI21OPTREPBD2BWP30P140 U118 ( .A1(n57), .A2(n50), .B(n49), .ZN(N322) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[2]), .ZN(n52) );
  ND2OPTIBD2BWP30P140 U120 ( .A1(n86), .A2(i_data_bus[34]), .ZN(n51) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[1]), .ZN(n54) );
  ND2OPTIBD4BWP30P140 U122 ( .A1(n86), .A2(i_data_bus[33]), .ZN(n53) );
  INVD1BWP30P140 U123 ( .I(i_data_bus[0]), .ZN(n56) );
  ND2OPTIBD2BWP30P140 U124 ( .A1(n86), .A2(i_data_bus[32]), .ZN(n55) );
  INVD1BWP30P140 U125 ( .I(i_data_bus[15]), .ZN(n59) );
  ND2OPTIBD2BWP30P140 U126 ( .A1(n86), .A2(i_data_bus[47]), .ZN(n58) );
  OAI21OPTREPBD2BWP30P140 U127 ( .A1(n89), .A2(n59), .B(n58), .ZN(N334) );
  INVD1BWP30P140 U128 ( .I(i_data_bus[14]), .ZN(n61) );
  ND2OPTIBD2BWP30P140 U129 ( .A1(n86), .A2(i_data_bus[46]), .ZN(n60) );
  OAI21OPTREPBD2BWP30P140 U130 ( .A1(n89), .A2(n61), .B(n60), .ZN(N333) );
  INVD1BWP30P140 U131 ( .I(i_data_bus[13]), .ZN(n63) );
  ND2OPTIBD2BWP30P140 U132 ( .A1(n86), .A2(i_data_bus[45]), .ZN(n62) );
  OAI21OPTREPBD2BWP30P140 U133 ( .A1(n89), .A2(n63), .B(n62), .ZN(N332) );
  INVD1BWP30P140 U134 ( .I(i_data_bus[11]), .ZN(n65) );
  ND2OPTIBD2BWP30P140 U135 ( .A1(n86), .A2(i_data_bus[43]), .ZN(n64) );
  OAI21OPTREPBD2BWP30P140 U136 ( .A1(n89), .A2(n65), .B(n64), .ZN(N330) );
  INVD1BWP30P140 U137 ( .I(i_data_bus[20]), .ZN(n67) );
  ND2OPTIBD2BWP30P140 U138 ( .A1(n86), .A2(i_data_bus[52]), .ZN(n66) );
  OAI21OPTREPBD2BWP30P140 U139 ( .A1(n89), .A2(n67), .B(n66), .ZN(N339) );
  INVD1BWP30P140 U140 ( .I(i_data_bus[26]), .ZN(n69) );
  INVD1BWP30P140 U141 ( .I(i_data_bus[22]), .ZN(n71) );
  INVD1BWP30P140 U142 ( .I(i_data_bus[28]), .ZN(n75) );
  ND2OPTIBD2BWP30P140 U143 ( .A1(n86), .A2(i_data_bus[60]), .ZN(n74) );
  INVD1BWP30P140 U144 ( .I(i_data_bus[21]), .ZN(n77) );
  INVD1BWP30P140 U145 ( .I(i_data_bus[24]), .ZN(n79) );
  INVD1BWP30P140 U146 ( .I(i_data_bus[23]), .ZN(n81) );
  INVD1BWP30P140 U147 ( .I(i_data_bus[25]), .ZN(n83) );
  ND2OPTIBD2BWP30P140 U148 ( .A1(n86), .A2(i_data_bus[62]), .ZN(n84) );
  INVD1BWP30P140 U149 ( .I(n93), .ZN(n96) );
  OAI21D1BWP30P140 U150 ( .A1(n94), .A2(n96), .B(n95), .ZN(N354) );
  OAI31D1BWP30P140 U151 ( .A1(n99), .A2(n98), .A3(n97), .B(n105), .ZN(N353) );
  INVD1BWP30P140 U152 ( .I(i_data_bus[49]), .ZN(n100) );
  OAI22D1BWP30P140 U153 ( .A1(n105), .A2(n101), .B1(n126), .B2(n100), .ZN(N304) );
  INVD1BWP30P140 U154 ( .I(i_data_bus[51]), .ZN(n102) );
  OAI22D1BWP30P140 U155 ( .A1(n105), .A2(n103), .B1(n126), .B2(n102), .ZN(N306) );
  INVD4BWP30P140 U156 ( .I(n104), .ZN(n130) );
  INVD1BWP30P140 U157 ( .I(i_data_bus[60]), .ZN(n106) );
  MOAI22D1BWP30P140 U158 ( .A1(n130), .A2(n106), .B1(n128), .B2(i_data_bus[28]), .ZN(N315) );
  INVD1BWP30P140 U159 ( .I(i_data_bus[48]), .ZN(n107) );
  MOAI22D1BWP30P140 U160 ( .A1(n1), .A2(n107), .B1(n128), .B2(i_data_bus[16]), 
        .ZN(N303) );
  INVD1BWP30P140 U161 ( .I(i_data_bus[34]), .ZN(n108) );
  MOAI22D1BWP30P140 U162 ( .A1(n130), .A2(n108), .B1(n128), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140 U163 ( .I(i_data_bus[59]), .ZN(n110) );
  MOAI22D1BWP30P140 U164 ( .A1(n130), .A2(n110), .B1(n128), .B2(i_data_bus[27]), .ZN(N314) );
  INVD1BWP30P140 U165 ( .I(i_data_bus[47]), .ZN(n111) );
  MOAI22D1BWP30P140 U166 ( .A1(n1), .A2(n111), .B1(n128), .B2(i_data_bus[15]), 
        .ZN(N302) );
  INVD1BWP30P140 U167 ( .I(i_data_bus[33]), .ZN(n112) );
  MOAI22D1BWP30P140 U168 ( .A1(n130), .A2(n112), .B1(n128), .B2(i_data_bus[1]), 
        .ZN(N288) );
  INVD1BWP30P140 U169 ( .I(i_data_bus[58]), .ZN(n113) );
  MOAI22D1BWP30P140 U170 ( .A1(n130), .A2(n113), .B1(n128), .B2(i_data_bus[26]), .ZN(N313) );
  INVD1BWP30P140 U171 ( .I(i_data_bus[46]), .ZN(n114) );
  MOAI22D1BWP30P140 U172 ( .A1(n1), .A2(n114), .B1(n128), .B2(i_data_bus[14]), 
        .ZN(N301) );
  INVD1BWP30P140 U173 ( .I(i_data_bus[32]), .ZN(n115) );
  MOAI22D1BWP30P140 U174 ( .A1(n130), .A2(n115), .B1(n128), .B2(i_data_bus[0]), 
        .ZN(N287) );
  INVD1BWP30P140 U175 ( .I(i_data_bus[57]), .ZN(n116) );
  MOAI22D1BWP30P140 U176 ( .A1(n1), .A2(n116), .B1(n128), .B2(i_data_bus[25]), 
        .ZN(N312) );
  INVD1BWP30P140 U177 ( .I(i_data_bus[45]), .ZN(n117) );
  MOAI22D1BWP30P140 U178 ( .A1(n1), .A2(n117), .B1(n128), .B2(i_data_bus[13]), 
        .ZN(N300) );
  INVD1BWP30P140 U179 ( .I(i_data_bus[56]), .ZN(n118) );
  MOAI22D1BWP30P140 U180 ( .A1(n109), .A2(n118), .B1(n128), .B2(i_data_bus[24]), .ZN(N311) );
  INVD1BWP30P140 U181 ( .I(i_data_bus[44]), .ZN(n119) );
  MOAI22D1BWP30P140 U182 ( .A1(n1), .A2(n119), .B1(n128), .B2(i_data_bus[12]), 
        .ZN(N299) );
  INVD1BWP30P140 U183 ( .I(i_data_bus[55]), .ZN(n120) );
  MOAI22D1BWP30P140 U184 ( .A1(n130), .A2(n120), .B1(n128), .B2(i_data_bus[23]), .ZN(N310) );
  INVD1BWP30P140 U185 ( .I(i_data_bus[43]), .ZN(n121) );
  MOAI22D1BWP30P140 U186 ( .A1(n1), .A2(n121), .B1(n128), .B2(i_data_bus[11]), 
        .ZN(N298) );
  INVD1BWP30P140 U187 ( .I(i_data_bus[54]), .ZN(n122) );
  MOAI22D1BWP30P140 U188 ( .A1(n130), .A2(n122), .B1(n128), .B2(i_data_bus[22]), .ZN(N309) );
  INVD1BWP30P140 U189 ( .I(i_data_bus[42]), .ZN(n123) );
  MOAI22D1BWP30P140 U190 ( .A1(n1), .A2(n123), .B1(n128), .B2(i_data_bus[10]), 
        .ZN(N297) );
  INVD1BWP30P140 U191 ( .I(i_data_bus[53]), .ZN(n124) );
  MOAI22D1BWP30P140 U192 ( .A1(n130), .A2(n124), .B1(n128), .B2(i_data_bus[21]), .ZN(N308) );
  INVD1BWP30P140 U193 ( .I(i_data_bus[41]), .ZN(n125) );
  MOAI22D1BWP30P140 U194 ( .A1(n1), .A2(n125), .B1(n128), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140 U195 ( .I(i_data_bus[52]), .ZN(n127) );
  MOAI22D1BWP30P140 U196 ( .A1(n130), .A2(n127), .B1(n128), .B2(i_data_bus[20]), .ZN(N307) );
  INVD1BWP30P140 U197 ( .I(i_data_bus[40]), .ZN(n129) );
  MOAI22D1BWP30P140 U198 ( .A1(n130), .A2(n129), .B1(n128), .B2(i_data_bus[8]), 
        .ZN(N295) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_134 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  CKND2D2BWP30P140 U3 ( .A1(n63), .A2(i_data_bus[55]), .ZN(n31) );
  CKND2D2BWP30P140 U4 ( .A1(n63), .A2(i_data_bus[37]), .ZN(n45) );
  CKND2D2BWP30P140 U5 ( .A1(n63), .A2(i_data_bus[54]), .ZN(n33) );
  CKND2D2BWP30P140 U6 ( .A1(n63), .A2(i_data_bus[36]), .ZN(n46) );
  CKND2D2BWP30P140 U7 ( .A1(n63), .A2(i_data_bus[35]), .ZN(n47) );
  CKND2D2BWP30P140 U8 ( .A1(n63), .A2(i_data_bus[42]), .ZN(n35) );
  CKND2D2BWP30P140 U9 ( .A1(n63), .A2(i_data_bus[40]), .ZN(n39) );
  CKND2D2BWP30P140 U10 ( .A1(n63), .A2(i_data_bus[53]), .ZN(n37) );
  CKND2D3BWP30P140 U11 ( .A1(i_valid[0]), .A2(n70), .ZN(n2) );
  CKND2D2BWP30P140 U12 ( .A1(n63), .A2(i_data_bus[63]), .ZN(n10) );
  INVD1BWP30P140 U13 ( .I(i_cmd[0]), .ZN(n1) );
  NR2OPTPAD2BWP30P140 U14 ( .A1(n1), .A2(n94), .ZN(n69) );
  INVD3BWP30P140 U15 ( .I(i_valid[0]), .ZN(n67) );
  INVD4BWP30P140 U16 ( .I(i_valid[1]), .ZN(n3) );
  CKND2D3BWP30P140 U17 ( .A1(n63), .A2(i_data_bus[45]), .ZN(n58) );
  INVD4BWP30P140 U18 ( .I(n2), .ZN(n90) );
  MUX2NOPTD4BWP30P140 U19 ( .I0(n67), .I1(n3), .S(i_cmd[1]), .ZN(n68) );
  INVD6BWP30P140 U20 ( .I(n7), .ZN(n13) );
  IOA21D2BWP30P140 U21 ( .A1(n13), .A2(i_data_bus[31]), .B(n10), .ZN(N350) );
  ND2OPTPAD6BWP30P140 U22 ( .A1(n90), .A2(n93), .ZN(n99) );
  ND2OPTPAD4BWP30P140 U23 ( .A1(n69), .A2(n68), .ZN(n123) );
  NR2OPTPAD1BWP30P140 U24 ( .A1(i_cmd[1]), .A2(n94), .ZN(n5) );
  OAI21D2BWP30P140 U25 ( .A1(n62), .A2(n59), .B(n58), .ZN(N332) );
  CKND2D4BWP30P140 U26 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n8) );
  INVD3BWP30P140 U27 ( .I(n8), .ZN(n9) );
  CKND2D2BWP30P140 U28 ( .A1(n63), .A2(i_data_bus[33]), .ZN(n50) );
  CKND2D2BWP30P140 U29 ( .A1(n63), .A2(i_data_bus[43]), .ZN(n60) );
  INVD3BWP30P140 U30 ( .I(i_cmd[0]), .ZN(n93) );
  OAI21D2BWP30P140 U31 ( .A1(n62), .A2(n61), .B(n60), .ZN(N330) );
  OAI21D2BWP30P140 U32 ( .A1(n66), .A2(n51), .B(n50), .ZN(N320) );
  CKND2D3BWP30P140 U33 ( .A1(n63), .A2(i_data_bus[34]), .ZN(n64) );
  OAI21D2BWP30P140 U34 ( .A1(n66), .A2(n65), .B(n64), .ZN(N321) );
  CKND2D4BWP30P140 U35 ( .A1(n6), .A2(n5), .ZN(n7) );
  ND2OPTIBD1BWP30P140 U36 ( .A1(n89), .A2(n88), .ZN(N318) );
  OR2D1BWP30P140 U37 ( .A1(n99), .A2(n87), .Z(n88) );
  ND2OPTIBD1BWP30P140 U38 ( .A1(n101), .A2(i_data_bus[63]), .ZN(n89) );
  MUX2NOPTD4BWP30P140 U39 ( .I0(n67), .I1(n3), .S(i_cmd[0]), .ZN(n6) );
  INVD1BWP30P140 U40 ( .I(rst), .ZN(n4) );
  ND2D1BWP30P140 U41 ( .A1(n4), .A2(i_en), .ZN(n94) );
  INVD1BWP30P140 U42 ( .I(n94), .ZN(n70) );
  ND2OPTPAD6BWP30P140 U43 ( .A1(n9), .A2(n70), .ZN(n91) );
  INVD15BWP30P140 U44 ( .I(n91), .ZN(n63) );
  INVD6BWP30P140 U45 ( .I(n13), .ZN(n66) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[27]), .ZN(n12) );
  ND2OPTIBD4BWP30P140 U47 ( .A1(n63), .A2(i_data_bus[59]), .ZN(n11) );
  OAI21D2BWP30P140 U48 ( .A1(n66), .A2(n12), .B(n11), .ZN(N346) );
  INVD8BWP30P140 U49 ( .I(n13), .ZN(n62) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[30]), .ZN(n96) );
  ND2OPTIBD4BWP30P140 U51 ( .A1(n63), .A2(i_data_bus[62]), .ZN(n14) );
  OAI21D2BWP30P140 U52 ( .A1(n62), .A2(n96), .B(n14), .ZN(N349) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[19]), .ZN(n71) );
  ND2OPTIBD4BWP30P140 U54 ( .A1(n63), .A2(i_data_bus[51]), .ZN(n15) );
  OAI21D2BWP30P140 U55 ( .A1(n66), .A2(n71), .B(n15), .ZN(N338) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[29]), .ZN(n98) );
  ND2OPTIBD4BWP30P140 U57 ( .A1(n63), .A2(i_data_bus[61]), .ZN(n16) );
  OAI21D2BWP30P140 U58 ( .A1(n62), .A2(n98), .B(n16), .ZN(N348) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[18]), .ZN(n73) );
  ND2OPTIBD4BWP30P140 U60 ( .A1(n63), .A2(i_data_bus[50]), .ZN(n17) );
  OAI21D2BWP30P140 U61 ( .A1(n66), .A2(n73), .B(n17), .ZN(N337) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[28]), .ZN(n19) );
  ND2OPTIBD4BWP30P140 U63 ( .A1(n63), .A2(i_data_bus[60]), .ZN(n18) );
  OAI21D2BWP30P140 U64 ( .A1(n62), .A2(n19), .B(n18), .ZN(N347) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[26]), .ZN(n21) );
  ND2OPTIBD4BWP30P140 U66 ( .A1(n63), .A2(i_data_bus[58]), .ZN(n20) );
  OAI21D2BWP30P140 U67 ( .A1(n62), .A2(n21), .B(n20), .ZN(N345) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[17]), .ZN(n75) );
  ND2OPTIBD4BWP30P140 U69 ( .A1(n63), .A2(i_data_bus[49]), .ZN(n22) );
  OAI21D2BWP30P140 U70 ( .A1(n66), .A2(n75), .B(n22), .ZN(N336) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[25]), .ZN(n24) );
  ND2OPTIBD4BWP30P140 U72 ( .A1(n63), .A2(i_data_bus[57]), .ZN(n23) );
  OAI21D2BWP30P140 U73 ( .A1(n62), .A2(n24), .B(n23), .ZN(N344) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[14]), .ZN(n26) );
  ND2OPTIBD4BWP30P140 U75 ( .A1(n63), .A2(i_data_bus[46]), .ZN(n25) );
  OAI21D2BWP30P140 U76 ( .A1(n66), .A2(n26), .B(n25), .ZN(N333) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[24]), .ZN(n28) );
  ND2OPTIBD4BWP30P140 U78 ( .A1(n63), .A2(i_data_bus[56]), .ZN(n27) );
  OAI21D2BWP30P140 U79 ( .A1(n62), .A2(n28), .B(n27), .ZN(N343) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[12]), .ZN(n30) );
  ND2OPTIBD4BWP30P140 U81 ( .A1(n63), .A2(i_data_bus[44]), .ZN(n29) );
  OAI21D2BWP30P140 U82 ( .A1(n66), .A2(n30), .B(n29), .ZN(N331) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[23]), .ZN(n32) );
  OAI21D2BWP30P140 U84 ( .A1(n62), .A2(n32), .B(n31), .ZN(N342) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[22]), .ZN(n34) );
  OAI21D2BWP30P140 U86 ( .A1(n62), .A2(n34), .B(n33), .ZN(N341) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[10]), .ZN(n36) );
  OAI21D2BWP30P140 U88 ( .A1(n66), .A2(n36), .B(n35), .ZN(N329) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[21]), .ZN(n38) );
  OAI21D2BWP30P140 U90 ( .A1(n62), .A2(n38), .B(n37), .ZN(N340) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[8]), .ZN(n40) );
  OAI21D2BWP30P140 U92 ( .A1(n66), .A2(n40), .B(n39), .ZN(N327) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[0]), .ZN(n42) );
  CKND2D3BWP30P140 U94 ( .A1(n63), .A2(i_data_bus[32]), .ZN(n41) );
  OAI21D2BWP30P140 U95 ( .A1(n62), .A2(n42), .B(n41), .ZN(N319) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[7]), .ZN(n79) );
  ND2OPTIBD4BWP30P140 U97 ( .A1(n63), .A2(i_data_bus[39]), .ZN(n43) );
  OAI21D2BWP30P140 U98 ( .A1(n66), .A2(n79), .B(n43), .ZN(N326) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[6]), .ZN(n83) );
  ND2OPTIBD4BWP30P140 U100 ( .A1(n63), .A2(i_data_bus[38]), .ZN(n44) );
  OAI21D2BWP30P140 U101 ( .A1(n66), .A2(n83), .B(n44), .ZN(N325) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[5]), .ZN(n85) );
  OAI21D2BWP30P140 U103 ( .A1(n66), .A2(n85), .B(n45), .ZN(N324) );
  INVD1BWP30P140 U104 ( .I(i_data_bus[4]), .ZN(n81) );
  OAI21D2BWP30P140 U105 ( .A1(n66), .A2(n81), .B(n46), .ZN(N323) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[3]), .ZN(n77) );
  OAI21D2BWP30P140 U107 ( .A1(n66), .A2(n77), .B(n47), .ZN(N322) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[9]), .ZN(n49) );
  ND2D2BWP30P140 U109 ( .A1(n63), .A2(i_data_bus[41]), .ZN(n48) );
  OAI21OPTREPBD2BWP30P140 U110 ( .A1(n62), .A2(n49), .B(n48), .ZN(N328) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[1]), .ZN(n51) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[20]), .ZN(n53) );
  ND2D2BWP30P140 U113 ( .A1(n63), .A2(i_data_bus[52]), .ZN(n52) );
  OAI21OPTREPBD2BWP30P140 U114 ( .A1(n62), .A2(n53), .B(n52), .ZN(N339) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[16]), .ZN(n55) );
  ND2D2BWP30P140 U116 ( .A1(n63), .A2(i_data_bus[48]), .ZN(n54) );
  OAI21OPTREPBD2BWP30P140 U117 ( .A1(n62), .A2(n55), .B(n54), .ZN(N335) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[15]), .ZN(n57) );
  ND2D2BWP30P140 U119 ( .A1(n63), .A2(i_data_bus[47]), .ZN(n56) );
  OAI21OPTREPBD2BWP30P140 U120 ( .A1(n62), .A2(n57), .B(n56), .ZN(N334) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[13]), .ZN(n59) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[11]), .ZN(n61) );
  INVD1BWP30P140 U123 ( .I(i_data_bus[2]), .ZN(n65) );
  INVD4BWP30P140 U124 ( .I(n123), .ZN(n101) );
  INVD4BWP30P140 U125 ( .I(n101), .ZN(n112) );
  INVD1BWP30P140 U126 ( .I(i_data_bus[51]), .ZN(n72) );
  OAI22OPTPBD1BWP30P140 U127 ( .A1(n112), .A2(n72), .B1(n99), .B2(n71), .ZN(
        N306) );
  INVD1BWP30P140 U128 ( .I(i_data_bus[50]), .ZN(n74) );
  OAI22OPTPBD1BWP30P140 U129 ( .A1(n112), .A2(n74), .B1(n99), .B2(n73), .ZN(
        N305) );
  INVD1BWP30P140 U130 ( .I(i_data_bus[49]), .ZN(n76) );
  OAI22OPTPBD1BWP30P140 U131 ( .A1(n112), .A2(n76), .B1(n99), .B2(n75), .ZN(
        N304) );
  INVD1BWP30P140 U132 ( .I(i_data_bus[35]), .ZN(n78) );
  OAI22OPTPBD1BWP30P140 U133 ( .A1(n112), .A2(n78), .B1(n99), .B2(n77), .ZN(
        N290) );
  INVD1BWP30P140 U134 ( .I(i_data_bus[39]), .ZN(n80) );
  OAI22OPTPBD1BWP30P140 U135 ( .A1(n112), .A2(n80), .B1(n99), .B2(n79), .ZN(
        N294) );
  INVD1BWP30P140 U136 ( .I(i_data_bus[36]), .ZN(n82) );
  OAI22OPTPBD1BWP30P140 U137 ( .A1(n112), .A2(n82), .B1(n99), .B2(n81), .ZN(
        N291) );
  INVD1BWP30P140 U138 ( .I(i_data_bus[38]), .ZN(n84) );
  OAI22OPTPBD1BWP30P140 U139 ( .A1(n112), .A2(n84), .B1(n99), .B2(n83), .ZN(
        N293) );
  INVD1BWP30P140 U140 ( .I(i_data_bus[37]), .ZN(n86) );
  OAI22OPTPBD1BWP30P140 U141 ( .A1(n112), .A2(n86), .B1(n99), .B2(n85), .ZN(
        N292) );
  INVD1BWP30P140 U142 ( .I(i_data_bus[31]), .ZN(n87) );
  INVD1BWP30P140 U143 ( .I(n90), .ZN(n92) );
  OAI21D1BWP30P140 U144 ( .A1(n92), .A2(i_cmd[1]), .B(n91), .ZN(N354) );
  OAI31D1BWP30P140 U145 ( .A1(n94), .A2(n3), .A3(n93), .B(n99), .ZN(N353) );
  INVD1BWP30P140 U146 ( .I(i_data_bus[62]), .ZN(n95) );
  OAI22D1BWP30P140 U147 ( .A1(n99), .A2(n96), .B1(n123), .B2(n95), .ZN(N317)
         );
  INVD1BWP30P140 U148 ( .I(i_data_bus[61]), .ZN(n97) );
  OAI22D1BWP30P140 U149 ( .A1(n99), .A2(n98), .B1(n123), .B2(n97), .ZN(N316)
         );
  BUFFD4BWP30P140 U150 ( .I(n123), .Z(n120) );
  INVD1BWP30P140 U151 ( .I(i_data_bus[60]), .ZN(n100) );
  INVD8BWP30P140 U152 ( .I(n99), .ZN(n124) );
  MOAI22D1BWP30P140 U153 ( .A1(n120), .A2(n100), .B1(n124), .B2(i_data_bus[28]), .ZN(N315) );
  INVD4BWP30P140 U154 ( .I(n101), .ZN(n126) );
  INVD1BWP30P140 U155 ( .I(i_data_bus[48]), .ZN(n102) );
  MOAI22D1BWP30P140 U156 ( .A1(n126), .A2(n102), .B1(n124), .B2(i_data_bus[16]), .ZN(N303) );
  INVD1BWP30P140 U157 ( .I(i_data_bus[34]), .ZN(n103) );
  MOAI22D1BWP30P140 U158 ( .A1(n126), .A2(n103), .B1(n124), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140 U159 ( .I(i_data_bus[59]), .ZN(n104) );
  MOAI22D1BWP30P140 U160 ( .A1(n120), .A2(n104), .B1(n124), .B2(i_data_bus[27]), .ZN(N314) );
  INVD1BWP30P140 U161 ( .I(i_data_bus[47]), .ZN(n105) );
  MOAI22D1BWP30P140 U162 ( .A1(n126), .A2(n105), .B1(n124), .B2(i_data_bus[15]), .ZN(N302) );
  INVD1BWP30P140 U163 ( .I(i_data_bus[33]), .ZN(n106) );
  MOAI22D1BWP30P140 U164 ( .A1(n126), .A2(n106), .B1(n124), .B2(i_data_bus[1]), 
        .ZN(N288) );
  INVD1BWP30P140 U165 ( .I(i_data_bus[58]), .ZN(n107) );
  MOAI22D1BWP30P140 U166 ( .A1(n120), .A2(n107), .B1(n124), .B2(i_data_bus[26]), .ZN(N313) );
  INVD1BWP30P140 U167 ( .I(i_data_bus[46]), .ZN(n108) );
  MOAI22D1BWP30P140 U168 ( .A1(n126), .A2(n108), .B1(n124), .B2(i_data_bus[14]), .ZN(N301) );
  INVD1BWP30P140 U169 ( .I(i_data_bus[32]), .ZN(n109) );
  MOAI22D1BWP30P140 U170 ( .A1(n126), .A2(n109), .B1(n124), .B2(i_data_bus[0]), 
        .ZN(N287) );
  INVD1BWP30P140 U171 ( .I(i_data_bus[57]), .ZN(n110) );
  MOAI22D1BWP30P140 U172 ( .A1(n120), .A2(n110), .B1(n124), .B2(i_data_bus[25]), .ZN(N312) );
  INVD1BWP30P140 U173 ( .I(i_data_bus[45]), .ZN(n111) );
  MOAI22D1BWP30P140 U174 ( .A1(n112), .A2(n111), .B1(n124), .B2(i_data_bus[13]), .ZN(N300) );
  INVD1BWP30P140 U175 ( .I(i_data_bus[56]), .ZN(n113) );
  MOAI22D1BWP30P140 U176 ( .A1(n120), .A2(n113), .B1(n124), .B2(i_data_bus[24]), .ZN(N311) );
  INVD1BWP30P140 U177 ( .I(i_data_bus[44]), .ZN(n114) );
  MOAI22D1BWP30P140 U178 ( .A1(n126), .A2(n114), .B1(n124), .B2(i_data_bus[12]), .ZN(N299) );
  INVD1BWP30P140 U179 ( .I(i_data_bus[55]), .ZN(n115) );
  MOAI22D1BWP30P140 U180 ( .A1(n120), .A2(n115), .B1(n124), .B2(i_data_bus[23]), .ZN(N310) );
  INVD1BWP30P140 U181 ( .I(i_data_bus[43]), .ZN(n116) );
  MOAI22D1BWP30P140 U182 ( .A1(n126), .A2(n116), .B1(n124), .B2(i_data_bus[11]), .ZN(N298) );
  INVD1BWP30P140 U183 ( .I(i_data_bus[54]), .ZN(n117) );
  MOAI22D1BWP30P140 U184 ( .A1(n120), .A2(n117), .B1(n124), .B2(i_data_bus[22]), .ZN(N309) );
  INVD1BWP30P140 U185 ( .I(i_data_bus[42]), .ZN(n118) );
  MOAI22D1BWP30P140 U186 ( .A1(n126), .A2(n118), .B1(n124), .B2(i_data_bus[10]), .ZN(N297) );
  INVD1BWP30P140 U187 ( .I(i_data_bus[53]), .ZN(n119) );
  MOAI22D1BWP30P140 U188 ( .A1(n120), .A2(n119), .B1(n124), .B2(i_data_bus[21]), .ZN(N308) );
  INVD1BWP30P140 U189 ( .I(i_data_bus[41]), .ZN(n121) );
  MOAI22D1BWP30P140 U190 ( .A1(n126), .A2(n121), .B1(n124), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140 U191 ( .I(i_data_bus[52]), .ZN(n122) );
  MOAI22D1BWP30P140 U192 ( .A1(n123), .A2(n122), .B1(n124), .B2(i_data_bus[20]), .ZN(N307) );
  INVD1BWP30P140 U193 ( .I(i_data_bus[40]), .ZN(n125) );
  MOAI22D1BWP30P140 U194 ( .A1(n126), .A2(n125), .B1(n124), .B2(i_data_bus[8]), 
        .ZN(N295) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_135 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI21D1BWP30P140 U3 ( .A1(n90), .A2(n72), .B(n71), .ZN(N339) );
  ND2OPTPAD6BWP30P140 U4 ( .A1(n76), .A2(n79), .ZN(n96) );
  CKND2D3BWP30P140 U5 ( .A1(i_valid[0]), .A2(n1), .ZN(n5) );
  INVD12BWP30P140 U6 ( .I(n96), .ZN(n119) );
  INVD4BWP30P140 U7 ( .I(i_valid[0]), .ZN(n18) );
  ND2OPTPAD6BWP30P140 U8 ( .A1(n7), .A2(n3), .ZN(n121) );
  BUFFD2BWP30P140 U9 ( .I(n121), .Z(n2) );
  INVD4BWP30P140 U10 ( .I(n42), .ZN(n90) );
  INVD3BWP30P140 U11 ( .I(i_cmd[1]), .ZN(n16) );
  OAI21D1BWP30P140 U12 ( .A1(n93), .A2(n83), .B(n73), .ZN(N338) );
  ND2D1BWP30P140 U13 ( .A1(n75), .A2(n74), .ZN(N305) );
  INVD1BWP30P140 U14 ( .I(n81), .ZN(n1) );
  INVD3BWP30P140 U15 ( .I(n4), .ZN(n3) );
  INVD8BWP30P140 U16 ( .I(n77), .ZN(n92) );
  INVD3BWP30P140 U17 ( .I(n21), .ZN(n42) );
  CKND2D2BWP30P140 U18 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n22) );
  INVD3BWP30P140 U19 ( .I(i_cmd[0]), .ZN(n79) );
  CKND2D3BWP30P140 U20 ( .A1(i_cmd[0]), .A2(n1), .ZN(n4) );
  INVD6BWP30P140 U21 ( .I(n121), .ZN(n95) );
  MUX2NOPTD4BWP30P140 U22 ( .I0(n18), .I1(n17), .S(i_cmd[0]), .ZN(n19) );
  INVD4BWP30P140 U23 ( .I(n42), .ZN(n93) );
  INVD4BWP30P140 U24 ( .I(n5), .ZN(n76) );
  OR2D1BWP30P140 U25 ( .A1(n96), .A2(n85), .Z(n74) );
  ND2OPTIBD1BWP30P140 U26 ( .A1(n95), .A2(i_data_bus[50]), .ZN(n75) );
  ND2D1BWP30P140 U27 ( .A1(n92), .A2(i_data_bus[40]), .ZN(n40) );
  ND2D1BWP30P140 U28 ( .A1(n92), .A2(i_data_bus[41]), .ZN(n43) );
  ND2D1BWP30P140 U29 ( .A1(n92), .A2(i_data_bus[42]), .ZN(n45) );
  ND2D1BWP30P140 U30 ( .A1(n92), .A2(i_data_bus[44]), .ZN(n47) );
  ND2D1BWP30P140 U31 ( .A1(n92), .A2(i_data_bus[52]), .ZN(n71) );
  ND2D1BWP30P140 U32 ( .A1(n92), .A2(i_data_bus[53]), .ZN(n69) );
  ND2D1BWP30P140 U33 ( .A1(n92), .A2(i_data_bus[54]), .ZN(n67) );
  ND2D1BWP30P140 U34 ( .A1(n92), .A2(i_data_bus[55]), .ZN(n65) );
  ND2D1BWP30P140 U35 ( .A1(n92), .A2(i_data_bus[56]), .ZN(n63) );
  ND2D1BWP30P140 U36 ( .A1(n92), .A2(i_data_bus[57]), .ZN(n61) );
  ND2D1BWP30P140 U37 ( .A1(n92), .A2(i_data_bus[58]), .ZN(n59) );
  ND2D1BWP30P140 U38 ( .A1(n92), .A2(i_data_bus[59]), .ZN(n57) );
  ND2D1BWP30P140 U39 ( .A1(n92), .A2(i_data_bus[60]), .ZN(n55) );
  ND2D1BWP30P140 U40 ( .A1(n92), .A2(i_data_bus[61]), .ZN(n53) );
  ND2D1BWP30P140 U41 ( .A1(n92), .A2(i_data_bus[62]), .ZN(n51) );
  ND2D1BWP30P140 U42 ( .A1(n92), .A2(i_data_bus[63]), .ZN(n49) );
  ND2D1BWP30P140 U43 ( .A1(n92), .A2(i_data_bus[32]), .ZN(n36) );
  ND2D1BWP30P140 U44 ( .A1(n92), .A2(i_data_bus[33]), .ZN(n34) );
  ND2D1BWP30P140 U45 ( .A1(n92), .A2(i_data_bus[34]), .ZN(n32) );
  ND2D1BWP30P140 U46 ( .A1(n92), .A2(i_data_bus[35]), .ZN(n24) );
  ND2D1BWP30P140 U47 ( .A1(n92), .A2(i_data_bus[36]), .ZN(n26) );
  ND2D1BWP30P140 U48 ( .A1(n92), .A2(i_data_bus[37]), .ZN(n28) );
  ND2D1BWP30P140 U49 ( .A1(n92), .A2(i_data_bus[38]), .ZN(n30) );
  ND2D1BWP30P140 U50 ( .A1(n92), .A2(i_data_bus[39]), .ZN(n38) );
  ND2D1BWP30P140 U51 ( .A1(n92), .A2(i_data_bus[51]), .ZN(n73) );
  INVD1BWP30P140 U52 ( .I(rst), .ZN(n6) );
  ND2D1BWP30P140 U53 ( .A1(n6), .A2(i_en), .ZN(n81) );
  INVD2BWP30P140 U54 ( .I(i_valid[1]), .ZN(n80) );
  MUX2NOPTD4BWP30P140 U55 ( .I0(n80), .I1(n18), .S(n16), .ZN(n7) );
  INVD4BWP30P140 U56 ( .I(n95), .ZN(n104) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[63]), .ZN(n8) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[31]), .ZN(n50) );
  OAI22OPTPBD1BWP30P140 U59 ( .A1(n104), .A2(n8), .B1(n96), .B2(n50), .ZN(N318) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[62]), .ZN(n9) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[30]), .ZN(n52) );
  OAI22OPTPBD1BWP30P140 U62 ( .A1(n104), .A2(n9), .B1(n96), .B2(n52), .ZN(N317) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[61]), .ZN(n10) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[29]), .ZN(n54) );
  OAI22OPTPBD1BWP30P140 U65 ( .A1(n104), .A2(n10), .B1(n96), .B2(n54), .ZN(
        N316) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[39]), .ZN(n11) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[7]), .ZN(n39) );
  OAI22OPTPBD1BWP30P140 U68 ( .A1(n104), .A2(n11), .B1(n96), .B2(n39), .ZN(
        N294) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[37]), .ZN(n12) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[5]), .ZN(n29) );
  OAI22OPTPBD1BWP30P140 U71 ( .A1(n104), .A2(n12), .B1(n96), .B2(n29), .ZN(
        N292) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[36]), .ZN(n13) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[4]), .ZN(n27) );
  OAI22OPTPBD1BWP30P140 U74 ( .A1(n104), .A2(n13), .B1(n96), .B2(n27), .ZN(
        N291) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[35]), .ZN(n14) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[3]), .ZN(n25) );
  OAI22OPTPBD1BWP30P140 U77 ( .A1(n104), .A2(n14), .B1(n96), .B2(n25), .ZN(
        N290) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[38]), .ZN(n15) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[6]), .ZN(n31) );
  OAI22OPTPBD1BWP30P140 U80 ( .A1(n104), .A2(n15), .B1(n96), .B2(n31), .ZN(
        N293) );
  NR2OPTPAD1BWP30P140 U81 ( .A1(i_cmd[1]), .A2(n81), .ZN(n20) );
  INVD2BWP30P140 U82 ( .I(i_valid[1]), .ZN(n17) );
  CKND2D3BWP30P140 U83 ( .A1(n19), .A2(n20), .ZN(n21) );
  INVD2BWP30P140 U84 ( .I(n22), .ZN(n23) );
  ND2OPTPAD4BWP30P140 U85 ( .A1(n23), .A2(n1), .ZN(n77) );
  OAI21D1BWP30P140 U86 ( .A1(n93), .A2(n25), .B(n24), .ZN(N322) );
  OAI21D1BWP30P140 U87 ( .A1(n93), .A2(n27), .B(n26), .ZN(N323) );
  OAI21D1BWP30P140 U88 ( .A1(n93), .A2(n29), .B(n28), .ZN(N324) );
  OAI21D1BWP30P140 U89 ( .A1(n93), .A2(n31), .B(n30), .ZN(N325) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[2]), .ZN(n33) );
  OAI21D1BWP30P140 U91 ( .A1(n93), .A2(n33), .B(n32), .ZN(N321) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[1]), .ZN(n35) );
  OAI21D1BWP30P140 U93 ( .A1(n93), .A2(n35), .B(n34), .ZN(N320) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[0]), .ZN(n37) );
  OAI21D1BWP30P140 U95 ( .A1(n93), .A2(n37), .B(n36), .ZN(N319) );
  OAI21D1BWP30P140 U96 ( .A1(n93), .A2(n39), .B(n38), .ZN(N326) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[8]), .ZN(n41) );
  OAI21D1BWP30P140 U98 ( .A1(n93), .A2(n41), .B(n40), .ZN(N327) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[9]), .ZN(n44) );
  OAI21D1BWP30P140 U100 ( .A1(n90), .A2(n44), .B(n43), .ZN(N328) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[10]), .ZN(n46) );
  OAI21D1BWP30P140 U102 ( .A1(n93), .A2(n46), .B(n45), .ZN(N329) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[12]), .ZN(n48) );
  OAI21D1BWP30P140 U104 ( .A1(n93), .A2(n48), .B(n47), .ZN(N331) );
  OAI21D1BWP30P140 U105 ( .A1(n90), .A2(n50), .B(n49), .ZN(N350) );
  OAI21D1BWP30P140 U106 ( .A1(n90), .A2(n52), .B(n51), .ZN(N349) );
  OAI21D1BWP30P140 U107 ( .A1(n90), .A2(n54), .B(n53), .ZN(N348) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[28]), .ZN(n56) );
  OAI21D1BWP30P140 U109 ( .A1(n90), .A2(n56), .B(n55), .ZN(N347) );
  INVD1BWP30P140 U110 ( .I(i_data_bus[27]), .ZN(n58) );
  OAI21D1BWP30P140 U111 ( .A1(n90), .A2(n58), .B(n57), .ZN(N346) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[26]), .ZN(n60) );
  OAI21D1BWP30P140 U113 ( .A1(n90), .A2(n60), .B(n59), .ZN(N345) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[25]), .ZN(n62) );
  OAI21D1BWP30P140 U115 ( .A1(n90), .A2(n62), .B(n61), .ZN(N344) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[24]), .ZN(n64) );
  OAI21D1BWP30P140 U117 ( .A1(n90), .A2(n64), .B(n63), .ZN(N343) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[23]), .ZN(n66) );
  OAI21D1BWP30P140 U119 ( .A1(n90), .A2(n66), .B(n65), .ZN(N342) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[22]), .ZN(n68) );
  OAI21D1BWP30P140 U121 ( .A1(n90), .A2(n68), .B(n67), .ZN(N341) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[21]), .ZN(n70) );
  OAI21D1BWP30P140 U123 ( .A1(n90), .A2(n70), .B(n69), .ZN(N340) );
  INVD1BWP30P140 U124 ( .I(i_data_bus[20]), .ZN(n72) );
  INVD1BWP30P140 U125 ( .I(i_data_bus[19]), .ZN(n83) );
  INVD1BWP30P140 U126 ( .I(i_data_bus[18]), .ZN(n85) );
  INVD1BWP30P140 U127 ( .I(n76), .ZN(n78) );
  OAI21D1BWP30P140 U128 ( .A1(i_cmd[1]), .A2(n78), .B(n77), .ZN(N354) );
  OAI31D1BWP30P140 U129 ( .A1(n81), .A2(n80), .A3(n79), .B(n96), .ZN(N353) );
  INVD1BWP30P140 U130 ( .I(i_data_bus[51]), .ZN(n82) );
  OAI22D1BWP30P140 U131 ( .A1(n96), .A2(n83), .B1(n121), .B2(n82), .ZN(N306)
         );
  INVD1BWP30P140 U132 ( .I(i_data_bus[17]), .ZN(n86) );
  INVD1BWP30P140 U133 ( .I(i_data_bus[49]), .ZN(n84) );
  OAI22D1BWP30P140 U134 ( .A1(n96), .A2(n86), .B1(n121), .B2(n84), .ZN(N304)
         );
  MOAI22D1BWP30P140 U135 ( .A1(n85), .A2(n93), .B1(i_data_bus[50]), .B2(n92), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U136 ( .A1(n86), .A2(n93), .B1(i_data_bus[49]), .B2(n92), 
        .ZN(N336) );
  INVD1BWP30P140 U137 ( .I(i_data_bus[16]), .ZN(n87) );
  MOAI22D1BWP30P140 U138 ( .A1(n87), .A2(n93), .B1(i_data_bus[48]), .B2(n92), 
        .ZN(N335) );
  INVD1BWP30P140 U139 ( .I(i_data_bus[15]), .ZN(n88) );
  MOAI22D1BWP30P140 U140 ( .A1(n88), .A2(n90), .B1(i_data_bus[47]), .B2(n92), 
        .ZN(N334) );
  INVD1BWP30P140 U141 ( .I(i_data_bus[14]), .ZN(n89) );
  MOAI22D1BWP30P140 U142 ( .A1(n89), .A2(n93), .B1(i_data_bus[46]), .B2(n92), 
        .ZN(N333) );
  INVD1BWP30P140 U143 ( .I(i_data_bus[13]), .ZN(n91) );
  MOAI22D1BWP30P140 U144 ( .A1(n91), .A2(n90), .B1(i_data_bus[45]), .B2(n92), 
        .ZN(N332) );
  INVD1BWP30P140 U145 ( .I(i_data_bus[11]), .ZN(n94) );
  MOAI22D1BWP30P140 U146 ( .A1(n94), .A2(n93), .B1(i_data_bus[43]), .B2(n92), 
        .ZN(N330) );
  INVD4BWP30P140 U147 ( .I(n95), .ZN(n118) );
  INVD1BWP30P140 U148 ( .I(i_data_bus[60]), .ZN(n97) );
  MOAI22D1BWP30P140 U149 ( .A1(n118), .A2(n97), .B1(n119), .B2(i_data_bus[28]), 
        .ZN(N315) );
  INVD1BWP30P140 U150 ( .I(i_data_bus[48]), .ZN(n98) );
  MOAI22D1BWP30P140 U151 ( .A1(n2), .A2(n98), .B1(n119), .B2(i_data_bus[16]), 
        .ZN(N303) );
  INVD1BWP30P140 U152 ( .I(i_data_bus[34]), .ZN(n99) );
  MOAI22D1BWP30P140 U153 ( .A1(n118), .A2(n99), .B1(n119), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140 U154 ( .I(i_data_bus[59]), .ZN(n100) );
  MOAI22D1BWP30P140 U155 ( .A1(n118), .A2(n100), .B1(n119), .B2(i_data_bus[27]), .ZN(N314) );
  INVD1BWP30P140 U156 ( .I(i_data_bus[47]), .ZN(n101) );
  MOAI22D1BWP30P140 U157 ( .A1(n2), .A2(n101), .B1(n119), .B2(i_data_bus[15]), 
        .ZN(N302) );
  INVD1BWP30P140 U158 ( .I(i_data_bus[33]), .ZN(n102) );
  MOAI22D1BWP30P140 U159 ( .A1(n118), .A2(n102), .B1(n119), .B2(i_data_bus[1]), 
        .ZN(N288) );
  INVD1BWP30P140 U160 ( .I(i_data_bus[58]), .ZN(n103) );
  MOAI22D1BWP30P140 U161 ( .A1(n104), .A2(n103), .B1(n119), .B2(i_data_bus[26]), .ZN(N313) );
  INVD1BWP30P140 U162 ( .I(i_data_bus[46]), .ZN(n105) );
  MOAI22D1BWP30P140 U163 ( .A1(n121), .A2(n105), .B1(n119), .B2(i_data_bus[14]), .ZN(N301) );
  INVD1BWP30P140 U164 ( .I(i_data_bus[32]), .ZN(n106) );
  MOAI22D1BWP30P140 U165 ( .A1(n118), .A2(n106), .B1(n119), .B2(i_data_bus[0]), 
        .ZN(N287) );
  INVD1BWP30P140 U166 ( .I(i_data_bus[57]), .ZN(n107) );
  MOAI22D1BWP30P140 U167 ( .A1(n118), .A2(n107), .B1(n119), .B2(i_data_bus[25]), .ZN(N312) );
  INVD1BWP30P140 U168 ( .I(i_data_bus[45]), .ZN(n108) );
  MOAI22D1BWP30P140 U169 ( .A1(n121), .A2(n108), .B1(n119), .B2(i_data_bus[13]), .ZN(N300) );
  INVD1BWP30P140 U170 ( .I(i_data_bus[56]), .ZN(n109) );
  MOAI22D1BWP30P140 U171 ( .A1(n118), .A2(n109), .B1(n119), .B2(i_data_bus[24]), .ZN(N311) );
  INVD1BWP30P140 U172 ( .I(i_data_bus[44]), .ZN(n110) );
  MOAI22D1BWP30P140 U173 ( .A1(n121), .A2(n110), .B1(n119), .B2(i_data_bus[12]), .ZN(N299) );
  INVD1BWP30P140 U174 ( .I(i_data_bus[55]), .ZN(n111) );
  MOAI22D1BWP30P140 U175 ( .A1(n118), .A2(n111), .B1(n119), .B2(i_data_bus[23]), .ZN(N310) );
  INVD1BWP30P140 U176 ( .I(i_data_bus[43]), .ZN(n112) );
  MOAI22D1BWP30P140 U177 ( .A1(n121), .A2(n112), .B1(n119), .B2(i_data_bus[11]), .ZN(N298) );
  INVD1BWP30P140 U178 ( .I(i_data_bus[54]), .ZN(n113) );
  MOAI22D1BWP30P140 U179 ( .A1(n118), .A2(n113), .B1(n119), .B2(i_data_bus[22]), .ZN(N309) );
  INVD1BWP30P140 U180 ( .I(i_data_bus[42]), .ZN(n114) );
  MOAI22D1BWP30P140 U181 ( .A1(n121), .A2(n114), .B1(n119), .B2(i_data_bus[10]), .ZN(N297) );
  INVD1BWP30P140 U182 ( .I(i_data_bus[53]), .ZN(n115) );
  MOAI22D1BWP30P140 U183 ( .A1(n118), .A2(n115), .B1(n119), .B2(i_data_bus[21]), .ZN(N308) );
  INVD1BWP30P140 U184 ( .I(i_data_bus[41]), .ZN(n116) );
  MOAI22D1BWP30P140 U185 ( .A1(n121), .A2(n116), .B1(n119), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140 U186 ( .I(i_data_bus[52]), .ZN(n117) );
  MOAI22D1BWP30P140 U187 ( .A1(n118), .A2(n117), .B1(n119), .B2(i_data_bus[20]), .ZN(N307) );
  INVD1BWP30P140 U188 ( .I(i_data_bus[40]), .ZN(n120) );
  MOAI22D1BWP30P140 U189 ( .A1(n121), .A2(n120), .B1(n119), .B2(i_data_bus[8]), 
        .ZN(N295) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_136 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  CKND2D4BWP30P140 U3 ( .A1(n9), .A2(n11), .ZN(n90) );
  INVD4BWP30P140 U4 ( .I(i_cmd[1]), .ZN(n12) );
  INVD8BWP30P140 U5 ( .I(n102), .ZN(n105) );
  OAI22OPTPBD2BWP30P140 U6 ( .A1(n100), .A2(n17), .B1(n105), .B2(n16), .ZN(
        N304) );
  OAI21D1BWP30P140 U7 ( .A1(n26), .A2(n7), .B(n25), .ZN(N346) );
  INVD8BWP30P140 U8 ( .I(n90), .ZN(n82) );
  INVD2BWP30P140 U9 ( .I(n8), .ZN(n9) );
  NR2D3BWP30P140 U10 ( .A1(n89), .A2(n94), .ZN(n6) );
  MUX2NOPTD2BWP30P140 U11 ( .I0(n13), .I1(n4), .S(i_cmd[0]), .ZN(n5) );
  INVD1BWP30P140 U12 ( .I(i_valid[1]), .ZN(n4) );
  INVD1BWP30P140 U13 ( .I(n12), .ZN(n89) );
  OAI22D1BWP30P140 U14 ( .A1(n105), .A2(n22), .B1(n100), .B2(n49), .ZN(N290)
         );
  OAI22D1BWP30P140 U15 ( .A1(n105), .A2(n21), .B1(n100), .B2(n51), .ZN(N291)
         );
  OAI22D1BWP30P140 U16 ( .A1(n105), .A2(n20), .B1(n100), .B2(n53), .ZN(N292)
         );
  OAI22D1BWP30P140 U17 ( .A1(n105), .A2(n24), .B1(n100), .B2(n55), .ZN(N293)
         );
  OAI22D1BWP30P140 U18 ( .A1(n105), .A2(n23), .B1(n100), .B2(n57), .ZN(N294)
         );
  OAI22D1BWP30P140 U19 ( .A1(n105), .A2(n18), .B1(n100), .B2(n34), .ZN(N305)
         );
  OAI22D1BWP30P140 U20 ( .A1(n105), .A2(n19), .B1(n100), .B2(n67), .ZN(N306)
         );
  ND2D1BWP30P140 U21 ( .A1(n87), .A2(n86), .ZN(N318) );
  ND2OPTIBD1BWP30P140 U22 ( .A1(n102), .A2(i_data_bus[63]), .ZN(n87) );
  OR2D1BWP30P140 U23 ( .A1(n100), .A2(n85), .Z(n86) );
  ND2D1BWP30P140 U24 ( .A1(n82), .A2(i_data_bus[32]), .ZN(n42) );
  ND2D1BWP30P140 U25 ( .A1(n82), .A2(i_data_bus[33]), .ZN(n44) );
  ND2D1BWP30P140 U26 ( .A1(n82), .A2(i_data_bus[34]), .ZN(n46) );
  ND2D1BWP30P140 U27 ( .A1(n82), .A2(i_data_bus[35]), .ZN(n48) );
  ND2D1BWP30P140 U28 ( .A1(n82), .A2(i_data_bus[36]), .ZN(n50) );
  ND2D1BWP30P140 U29 ( .A1(n82), .A2(i_data_bus[37]), .ZN(n52) );
  ND2D1BWP30P140 U30 ( .A1(n82), .A2(i_data_bus[38]), .ZN(n54) );
  ND2D1BWP30P140 U31 ( .A1(n82), .A2(i_data_bus[39]), .ZN(n56) );
  ND2D1BWP30P140 U32 ( .A1(n82), .A2(i_data_bus[40]), .ZN(n58) );
  ND2D1BWP30P140 U33 ( .A1(n82), .A2(i_data_bus[41]), .ZN(n60) );
  ND2D1BWP30P140 U34 ( .A1(n82), .A2(i_data_bus[42]), .ZN(n62) );
  ND2D1BWP30P140 U35 ( .A1(n82), .A2(i_data_bus[43]), .ZN(n64) );
  ND2D1BWP30P140 U36 ( .A1(n82), .A2(i_data_bus[44]), .ZN(n68) );
  ND2D1BWP30P140 U37 ( .A1(n82), .A2(i_data_bus[45]), .ZN(n70) );
  ND2D1BWP30P140 U38 ( .A1(n82), .A2(i_data_bus[46]), .ZN(n72) );
  ND2D1BWP30P140 U39 ( .A1(n82), .A2(i_data_bus[47]), .ZN(n74) );
  ND2D1BWP30P140 U40 ( .A1(n82), .A2(i_data_bus[48]), .ZN(n76) );
  OAI21D1BWP30P140 U41 ( .A1(n7), .A2(n17), .B(n10), .ZN(N336) );
  ND2D1BWP30P140 U42 ( .A1(n82), .A2(i_data_bus[49]), .ZN(n10) );
  ND2D1BWP30P140 U43 ( .A1(n82), .A2(i_data_bus[58]), .ZN(n31) );
  ND2OPTIBD6BWP30P140 U44 ( .A1(n15), .A2(n14), .ZN(n99) );
  CKND2D4BWP30P140 U45 ( .A1(n6), .A2(n5), .ZN(n1) );
  CKND2D4BWP30P140 U46 ( .A1(n6), .A2(n5), .ZN(n2) );
  INVD1BWP30P140 U47 ( .I(rst), .ZN(n3) );
  ND2D1BWP30P140 U48 ( .A1(n3), .A2(i_en), .ZN(n94) );
  INVD3BWP30P140 U49 ( .I(i_valid[0]), .ZN(n13) );
  CKND2D3BWP30P140 U50 ( .A1(n6), .A2(n5), .ZN(n7) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[17]), .ZN(n17) );
  CKND2D2BWP30P140 U52 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n8) );
  INVD1BWP30P140 U53 ( .I(n94), .ZN(n11) );
  AN2D4BWP30P140 U54 ( .A1(i_valid[0]), .A2(n11), .Z(n88) );
  INVD2BWP30P140 U55 ( .I(i_cmd[0]), .ZN(n92) );
  ND2OPTPAD8BWP30P140 U56 ( .A1(n88), .A2(n92), .ZN(n100) );
  INR2D4BWP30P140 U57 ( .A1(i_cmd[0]), .B1(n94), .ZN(n15) );
  INVD2BWP30P140 U58 ( .I(i_valid[1]), .ZN(n93) );
  MUX2NOPTD4BWP30P140 U59 ( .I0(n93), .I1(n13), .S(n12), .ZN(n14) );
  INVD6BWP30P140 U60 ( .I(n99), .ZN(n102) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[49]), .ZN(n16) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[50]), .ZN(n18) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[18]), .ZN(n34) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[51]), .ZN(n19) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[19]), .ZN(n67) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[37]), .ZN(n20) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[5]), .ZN(n53) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[36]), .ZN(n21) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[4]), .ZN(n51) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[35]), .ZN(n22) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[3]), .ZN(n49) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[39]), .ZN(n23) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[7]), .ZN(n57) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[38]), .ZN(n24) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[6]), .ZN(n55) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[27]), .ZN(n26) );
  ND2D1BWP30P140 U77 ( .A1(n82), .A2(i_data_bus[59]), .ZN(n25) );
  INVD1BWP30P140 U78 ( .I(i_data_bus[31]), .ZN(n85) );
  ND2D1BWP30P140 U79 ( .A1(n82), .A2(i_data_bus[63]), .ZN(n27) );
  OAI21D1BWP30P140 U80 ( .A1(n85), .A2(n7), .B(n27), .ZN(N350) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[29]), .ZN(n96) );
  ND2D1BWP30P140 U82 ( .A1(n82), .A2(i_data_bus[61]), .ZN(n28) );
  OAI21D1BWP30P140 U83 ( .A1(n96), .A2(n7), .B(n28), .ZN(N348) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[28]), .ZN(n30) );
  ND2D1BWP30P140 U85 ( .A1(n82), .A2(i_data_bus[60]), .ZN(n29) );
  OAI21D1BWP30P140 U86 ( .A1(n30), .A2(n7), .B(n29), .ZN(N347) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[26]), .ZN(n32) );
  OAI21D1BWP30P140 U88 ( .A1(n7), .A2(n32), .B(n31), .ZN(N345) );
  ND2D1BWP30P140 U89 ( .A1(n82), .A2(i_data_bus[50]), .ZN(n33) );
  OAI21D1BWP30P140 U90 ( .A1(n1), .A2(n34), .B(n33), .ZN(N337) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[30]), .ZN(n98) );
  ND2D1BWP30P140 U92 ( .A1(n82), .A2(i_data_bus[62]), .ZN(n35) );
  OAI21D1BWP30P140 U93 ( .A1(n2), .A2(n98), .B(n35), .ZN(N349) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[25]), .ZN(n37) );
  ND2D1BWP30P140 U95 ( .A1(n82), .A2(i_data_bus[57]), .ZN(n36) );
  OAI21D1BWP30P140 U96 ( .A1(n1), .A2(n37), .B(n36), .ZN(N344) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[24]), .ZN(n39) );
  ND2D1BWP30P140 U98 ( .A1(n82), .A2(i_data_bus[56]), .ZN(n38) );
  OAI21D1BWP30P140 U99 ( .A1(n2), .A2(n39), .B(n38), .ZN(N343) );
  INVD1BWP30P140 U100 ( .I(i_data_bus[23]), .ZN(n41) );
  ND2D1BWP30P140 U101 ( .A1(n82), .A2(i_data_bus[55]), .ZN(n40) );
  OAI21D1BWP30P140 U102 ( .A1(n1), .A2(n41), .B(n40), .ZN(N342) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[0]), .ZN(n43) );
  OAI21D1BWP30P140 U104 ( .A1(n2), .A2(n43), .B(n42), .ZN(N319) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[1]), .ZN(n45) );
  OAI21D1BWP30P140 U106 ( .A1(n1), .A2(n45), .B(n44), .ZN(N320) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[2]), .ZN(n47) );
  OAI21D1BWP30P140 U108 ( .A1(n2), .A2(n47), .B(n46), .ZN(N321) );
  OAI21D1BWP30P140 U109 ( .A1(n1), .A2(n49), .B(n48), .ZN(N322) );
  OAI21D1BWP30P140 U110 ( .A1(n2), .A2(n51), .B(n50), .ZN(N323) );
  OAI21D1BWP30P140 U111 ( .A1(n1), .A2(n53), .B(n52), .ZN(N324) );
  OAI21D1BWP30P140 U112 ( .A1(n2), .A2(n55), .B(n54), .ZN(N325) );
  OAI21D1BWP30P140 U113 ( .A1(n1), .A2(n57), .B(n56), .ZN(N326) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[8]), .ZN(n59) );
  OAI21D1BWP30P140 U115 ( .A1(n2), .A2(n59), .B(n58), .ZN(N327) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[9]), .ZN(n61) );
  OAI21D1BWP30P140 U117 ( .A1(n1), .A2(n61), .B(n60), .ZN(N328) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[10]), .ZN(n63) );
  OAI21D1BWP30P140 U119 ( .A1(n2), .A2(n63), .B(n62), .ZN(N329) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[11]), .ZN(n65) );
  OAI21D1BWP30P140 U121 ( .A1(n1), .A2(n65), .B(n64), .ZN(N330) );
  ND2D1BWP30P140 U122 ( .A1(n82), .A2(i_data_bus[51]), .ZN(n66) );
  OAI21D1BWP30P140 U123 ( .A1(n2), .A2(n67), .B(n66), .ZN(N338) );
  INVD1BWP30P140 U124 ( .I(i_data_bus[12]), .ZN(n69) );
  OAI21D1BWP30P140 U125 ( .A1(n1), .A2(n69), .B(n68), .ZN(N331) );
  INVD1BWP30P140 U126 ( .I(i_data_bus[13]), .ZN(n71) );
  OAI21D1BWP30P140 U127 ( .A1(n2), .A2(n71), .B(n70), .ZN(N332) );
  INVD1BWP30P140 U128 ( .I(i_data_bus[14]), .ZN(n73) );
  OAI21D1BWP30P140 U129 ( .A1(n1), .A2(n73), .B(n72), .ZN(N333) );
  INVD1BWP30P140 U130 ( .I(i_data_bus[15]), .ZN(n75) );
  OAI21D1BWP30P140 U131 ( .A1(n2), .A2(n75), .B(n74), .ZN(N334) );
  INVD1BWP30P140 U132 ( .I(i_data_bus[16]), .ZN(n77) );
  OAI21D1BWP30P140 U133 ( .A1(n1), .A2(n77), .B(n76), .ZN(N335) );
  INVD1BWP30P140 U134 ( .I(i_data_bus[22]), .ZN(n79) );
  ND2D1BWP30P140 U135 ( .A1(n82), .A2(i_data_bus[54]), .ZN(n78) );
  OAI21D1BWP30P140 U136 ( .A1(n2), .A2(n79), .B(n78), .ZN(N341) );
  INVD1BWP30P140 U137 ( .I(i_data_bus[21]), .ZN(n81) );
  ND2D1BWP30P140 U138 ( .A1(n82), .A2(i_data_bus[53]), .ZN(n80) );
  OAI21D1BWP30P140 U139 ( .A1(n1), .A2(n81), .B(n80), .ZN(N340) );
  INVD1BWP30P140 U140 ( .I(i_data_bus[20]), .ZN(n84) );
  ND2D1BWP30P140 U141 ( .A1(n82), .A2(i_data_bus[52]), .ZN(n83) );
  OAI21D1BWP30P140 U142 ( .A1(n2), .A2(n84), .B(n83), .ZN(N339) );
  INVD1BWP30P140 U143 ( .I(n88), .ZN(n91) );
  OAI21D1BWP30P140 U144 ( .A1(n91), .A2(n89), .B(n90), .ZN(N354) );
  OAI31D1BWP30P140 U145 ( .A1(n94), .A2(n93), .A3(n92), .B(n100), .ZN(N353) );
  INVD1BWP30P140 U146 ( .I(i_data_bus[61]), .ZN(n95) );
  OAI22D1BWP30P140 U147 ( .A1(n100), .A2(n96), .B1(n99), .B2(n95), .ZN(N316)
         );
  INVD1BWP30P140 U148 ( .I(i_data_bus[62]), .ZN(n97) );
  OAI22D1BWP30P140 U149 ( .A1(n100), .A2(n98), .B1(n99), .B2(n97), .ZN(N317)
         );
  INVD1BWP30P140 U150 ( .I(i_data_bus[60]), .ZN(n101) );
  INVD8BWP30P140 U151 ( .I(n100), .ZN(n123) );
  MOAI22D1BWP30P140 U152 ( .A1(n105), .A2(n101), .B1(n123), .B2(i_data_bus[28]), .ZN(N315) );
  INVD3BWP30P140 U153 ( .I(n102), .ZN(n125) );
  INVD1BWP30P140 U154 ( .I(i_data_bus[48]), .ZN(n103) );
  MOAI22D1BWP30P140 U155 ( .A1(n125), .A2(n103), .B1(n123), .B2(i_data_bus[16]), .ZN(N303) );
  INVD1BWP30P140 U156 ( .I(i_data_bus[34]), .ZN(n104) );
  MOAI22D1BWP30P140 U157 ( .A1(n105), .A2(n104), .B1(n123), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140 U158 ( .I(i_data_bus[59]), .ZN(n106) );
  MOAI22D1BWP30P140 U159 ( .A1(n105), .A2(n106), .B1(n123), .B2(i_data_bus[27]), .ZN(N314) );
  INVD1BWP30P140 U160 ( .I(i_data_bus[47]), .ZN(n107) );
  MOAI22D1BWP30P140 U161 ( .A1(n125), .A2(n107), .B1(n123), .B2(i_data_bus[15]), .ZN(N302) );
  INVD1BWP30P140 U162 ( .I(i_data_bus[33]), .ZN(n108) );
  MOAI22D1BWP30P140 U163 ( .A1(n125), .A2(n108), .B1(n123), .B2(i_data_bus[1]), 
        .ZN(N288) );
  INVD1BWP30P140 U164 ( .I(i_data_bus[58]), .ZN(n109) );
  MOAI22D1BWP30P140 U165 ( .A1(n105), .A2(n109), .B1(n123), .B2(i_data_bus[26]), .ZN(N313) );
  INVD1BWP30P140 U166 ( .I(i_data_bus[46]), .ZN(n110) );
  MOAI22D1BWP30P140 U167 ( .A1(n125), .A2(n110), .B1(n123), .B2(i_data_bus[14]), .ZN(N301) );
  INVD1BWP30P140 U168 ( .I(i_data_bus[32]), .ZN(n111) );
  MOAI22D1BWP30P140 U169 ( .A1(n125), .A2(n111), .B1(n123), .B2(i_data_bus[0]), 
        .ZN(N287) );
  INVD1BWP30P140 U170 ( .I(i_data_bus[57]), .ZN(n112) );
  MOAI22D1BWP30P140 U171 ( .A1(n105), .A2(n112), .B1(n123), .B2(i_data_bus[25]), .ZN(N312) );
  INVD1BWP30P140 U172 ( .I(i_data_bus[45]), .ZN(n113) );
  MOAI22D1BWP30P140 U173 ( .A1(n125), .A2(n113), .B1(n123), .B2(i_data_bus[13]), .ZN(N300) );
  INVD1BWP30P140 U174 ( .I(i_data_bus[56]), .ZN(n114) );
  MOAI22D1BWP30P140 U175 ( .A1(n105), .A2(n114), .B1(n123), .B2(i_data_bus[24]), .ZN(N311) );
  INVD1BWP30P140 U176 ( .I(i_data_bus[44]), .ZN(n115) );
  MOAI22D1BWP30P140 U177 ( .A1(n125), .A2(n115), .B1(n123), .B2(i_data_bus[12]), .ZN(N299) );
  INVD1BWP30P140 U178 ( .I(i_data_bus[55]), .ZN(n116) );
  MOAI22D1BWP30P140 U179 ( .A1(n105), .A2(n116), .B1(n123), .B2(i_data_bus[23]), .ZN(N310) );
  INVD1BWP30P140 U180 ( .I(i_data_bus[43]), .ZN(n117) );
  MOAI22D1BWP30P140 U181 ( .A1(n125), .A2(n117), .B1(n123), .B2(i_data_bus[11]), .ZN(N298) );
  INVD1BWP30P140 U182 ( .I(i_data_bus[54]), .ZN(n118) );
  MOAI22D1BWP30P140 U183 ( .A1(n105), .A2(n118), .B1(n123), .B2(i_data_bus[22]), .ZN(N309) );
  INVD1BWP30P140 U184 ( .I(i_data_bus[42]), .ZN(n119) );
  MOAI22D1BWP30P140 U185 ( .A1(n125), .A2(n119), .B1(n123), .B2(i_data_bus[10]), .ZN(N297) );
  INVD1BWP30P140 U186 ( .I(i_data_bus[53]), .ZN(n120) );
  MOAI22D1BWP30P140 U187 ( .A1(n105), .A2(n120), .B1(n123), .B2(i_data_bus[21]), .ZN(N308) );
  INVD1BWP30P140 U188 ( .I(i_data_bus[41]), .ZN(n121) );
  MOAI22D1BWP30P140 U189 ( .A1(n125), .A2(n121), .B1(n123), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140 U190 ( .I(i_data_bus[52]), .ZN(n122) );
  MOAI22D1BWP30P140 U191 ( .A1(n105), .A2(n122), .B1(n123), .B2(i_data_bus[20]), .ZN(N307) );
  INVD1BWP30P140 U192 ( .I(i_data_bus[40]), .ZN(n124) );
  MOAI22D1BWP30P140 U193 ( .A1(n125), .A2(n124), .B1(n123), .B2(i_data_bus[8]), 
        .ZN(N295) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_137 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI21D1BWP30P140 U3 ( .A1(n1), .A2(n59), .B(n58), .ZN(N334) );
  OAI21D1BWP30P140 U4 ( .A1(n1), .A2(n61), .B(n60), .ZN(N335) );
  OAI21D1BWP30P140 U5 ( .A1(n1), .A2(n68), .B(n67), .ZN(N340) );
  OAI21D1BWP30P140 U6 ( .A1(n1), .A2(n70), .B(n69), .ZN(N341) );
  OAI21D1BWP30P140 U7 ( .A1(n1), .A2(n17), .B(n16), .ZN(N320) );
  OAI21D1BWP30P140 U8 ( .A1(n1), .A2(n23), .B(n14), .ZN(N350) );
  OAI21D1BWP30P140 U9 ( .A1(n1), .A2(n84), .B(n83), .ZN(N348) );
  ND2OPTIBD1BWP30P140 U10 ( .A1(n87), .A2(i_data_bus[44]), .ZN(n52) );
  ND2OPTIBD1BWP30P140 U11 ( .A1(n87), .A2(i_data_bus[45]), .ZN(n54) );
  CKND2D2BWP30P140 U12 ( .A1(n87), .A2(i_data_bus[34]), .ZN(n88) );
  CKND2D2BWP30P140 U13 ( .A1(n87), .A2(i_data_bus[46]), .ZN(n56) );
  CKND2D2BWP30P140 U14 ( .A1(n87), .A2(i_data_bus[47]), .ZN(n58) );
  CKND2D2BWP30P140 U15 ( .A1(n87), .A2(i_data_bus[48]), .ZN(n60) );
  CKND2D2BWP30P140 U16 ( .A1(n87), .A2(i_data_bus[53]), .ZN(n67) );
  CKND2D2BWP30P140 U17 ( .A1(n87), .A2(i_data_bus[54]), .ZN(n69) );
  INVD4BWP30P140 U18 ( .I(n104), .ZN(n128) );
  NR2D1BWP30P140 U19 ( .A1(i_cmd[0]), .A2(i_valid[0]), .ZN(n6) );
  NR2D3BWP30P140 U20 ( .A1(n2), .A2(n98), .ZN(n21) );
  OAI21D1BWP30P140 U21 ( .A1(n1), .A2(n72), .B(n71), .ZN(N342) );
  CKND2D4BWP30P140 U22 ( .A1(n8), .A2(n9), .ZN(n7) );
  CKND2D4BWP30P140 U23 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n12) );
  INVD4BWP30P140 U24 ( .I(n12), .ZN(n13) );
  OAI21OPTREPBD1BWP30P140 U25 ( .A1(n1), .A2(n33), .B(n32), .ZN(N319) );
  INVD6BWP30P140 U26 ( .I(n103), .ZN(n108) );
  INVD4BWP30P140 U27 ( .I(i_cmd[1]), .ZN(n18) );
  INVD9BWP30P140 U28 ( .I(n15), .ZN(n1) );
  ND2OPTIBD8BWP30P140 U29 ( .A1(n20), .A2(n21), .ZN(n126) );
  OAI21D1BWP30P140 U30 ( .A1(n1), .A2(n74), .B(n73), .ZN(N343) );
  OAI21D1BWP30P140 U31 ( .A1(n1), .A2(n90), .B(n62), .ZN(N336) );
  OAI21D1BWP30P140 U32 ( .A1(n1), .A2(n76), .B(n75), .ZN(N344) );
  OAI21D1BWP30P140 U33 ( .A1(n1), .A2(n78), .B(n77), .ZN(N345) );
  OAI21D1BWP30P140 U34 ( .A1(n1), .A2(n80), .B(n79), .ZN(N346) );
  OAI21D1BWP30P140 U35 ( .A1(n1), .A2(n102), .B(n63), .ZN(N337) );
  OAI21D1BWP30P140 U36 ( .A1(n1), .A2(n100), .B(n64), .ZN(N338) );
  OAI21D1BWP30P140 U37 ( .A1(n1), .A2(n82), .B(n81), .ZN(N347) );
  ND2OPTPAD4BWP30P140 U38 ( .A1(n93), .A2(n96), .ZN(n104) );
  OAI21OPTREPBD1BWP30P140 U39 ( .A1(n1), .A2(n86), .B(n85), .ZN(N349) );
  INR2D4BWP30P140 U40 ( .A1(n22), .B1(n5), .ZN(n93) );
  OAI21D1BWP30P140 U41 ( .A1(n1), .A2(n66), .B(n65), .ZN(N339) );
  OAI21D1BWP30P140 U42 ( .A1(n1), .A2(n89), .B(n88), .ZN(N321) );
  INVD2BWP30P140 U43 ( .I(i_valid[1]), .ZN(n10) );
  INVD2BWP30P140 U44 ( .I(i_cmd[0]), .ZN(n2) );
  BUFFD4BWP30P140 U45 ( .I(n104), .Z(n3) );
  INVD1P5BWP30P140 U46 ( .I(i_cmd[0]), .ZN(n96) );
  OAI21D1BWP30P140 U47 ( .A1(n126), .A2(n125), .B(n4), .ZN(N296) );
  ND2D1BWP30P140 U48 ( .A1(n128), .A2(i_data_bus[9]), .ZN(n4) );
  INVD2BWP30P140 U49 ( .I(i_valid[0]), .ZN(n5) );
  NR2OPTPAD2BWP30P140 U50 ( .A1(i_cmd[1]), .A2(n98), .ZN(n8) );
  INVD2BWP30P140 U51 ( .I(i_valid[0]), .ZN(n19) );
  NR2OPTPAD4BWP30P140 U52 ( .A1(n7), .A2(n6), .ZN(n15) );
  ND2D2BWP30P140 U53 ( .A1(n10), .A2(i_cmd[0]), .ZN(n9) );
  ND2OPTIBD1BWP30P140 U54 ( .A1(n92), .A2(n91), .ZN(N304) );
  OR2D1BWP30P140 U55 ( .A1(n104), .A2(n90), .Z(n91) );
  ND2OPTIBD1BWP30P140 U56 ( .A1(n103), .A2(i_data_bus[49]), .ZN(n92) );
  OAI22D1BWP30P140 U57 ( .A1(n108), .A2(n26), .B1(n3), .B2(n84), .ZN(N316) );
  OAI22D1BWP30P140 U58 ( .A1(n108), .A2(n25), .B1(n3), .B2(n86), .ZN(N317) );
  OAI22D1BWP30P140 U59 ( .A1(n108), .A2(n24), .B1(n104), .B2(n23), .ZN(N318)
         );
  OAI22D1BWP30P140 U60 ( .A1(n108), .A2(n29), .B1(n3), .B2(n37), .ZN(N290) );
  OAI22D1BWP30P140 U61 ( .A1(n108), .A2(n28), .B1(n3), .B2(n39), .ZN(N291) );
  OAI22D1BWP30P140 U62 ( .A1(n108), .A2(n31), .B1(n3), .B2(n35), .ZN(N292) );
  OAI22D1BWP30P140 U63 ( .A1(n108), .A2(n30), .B1(n3), .B2(n41), .ZN(N293) );
  OAI22D1BWP30P140 U64 ( .A1(n108), .A2(n27), .B1(n3), .B2(n43), .ZN(N294) );
  CKND2D2BWP30P140 U65 ( .A1(n87), .A2(i_data_bus[32]), .ZN(n32) );
  CKND2D2BWP30P140 U66 ( .A1(n87), .A2(i_data_bus[61]), .ZN(n83) );
  CKND2D2BWP30P140 U67 ( .A1(n87), .A2(i_data_bus[62]), .ZN(n85) );
  INVD1BWP30P140 U68 ( .I(rst), .ZN(n11) );
  ND2D1BWP30P140 U69 ( .A1(n11), .A2(i_en), .ZN(n98) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[31]), .ZN(n23) );
  INVD1BWP30P140 U71 ( .I(n98), .ZN(n22) );
  ND2OPTPAD6BWP30P140 U72 ( .A1(n13), .A2(n22), .ZN(n94) );
  INVD15BWP30P140 U73 ( .I(n94), .ZN(n87) );
  ND2OPTIBD4BWP30P140 U74 ( .A1(n87), .A2(i_data_bus[63]), .ZN(n14) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[1]), .ZN(n17) );
  ND2OPTIBD4BWP30P140 U76 ( .A1(n87), .A2(i_data_bus[33]), .ZN(n16) );
  INVD2BWP30P140 U77 ( .I(i_valid[1]), .ZN(n97) );
  MUX2NOPTD4BWP30P140 U78 ( .I0(n97), .I1(n19), .S(n18), .ZN(n20) );
  INVD6BWP30P140 U79 ( .I(n126), .ZN(n103) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[63]), .ZN(n24) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[62]), .ZN(n25) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[30]), .ZN(n86) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[61]), .ZN(n26) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[29]), .ZN(n84) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[39]), .ZN(n27) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[7]), .ZN(n43) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[36]), .ZN(n28) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[4]), .ZN(n39) );
  INVD1BWP30P140 U89 ( .I(i_data_bus[35]), .ZN(n29) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[3]), .ZN(n37) );
  INVD1BWP30P140 U91 ( .I(i_data_bus[38]), .ZN(n30) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[6]), .ZN(n41) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[37]), .ZN(n31) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[5]), .ZN(n35) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[0]), .ZN(n33) );
  ND2OPTIBD4BWP30P140 U96 ( .A1(n87), .A2(i_data_bus[37]), .ZN(n34) );
  OAI21OPTREPBD1BWP30P140 U97 ( .A1(n1), .A2(n35), .B(n34), .ZN(N324) );
  ND2OPTIBD4BWP30P140 U98 ( .A1(n87), .A2(i_data_bus[35]), .ZN(n36) );
  OAI21OPTREPBD1BWP30P140 U99 ( .A1(n1), .A2(n37), .B(n36), .ZN(N322) );
  ND2OPTIBD4BWP30P140 U100 ( .A1(n87), .A2(i_data_bus[36]), .ZN(n38) );
  OAI21OPTREPBD1BWP30P140 U101 ( .A1(n1), .A2(n39), .B(n38), .ZN(N323) );
  ND2OPTIBD4BWP30P140 U102 ( .A1(n87), .A2(i_data_bus[38]), .ZN(n40) );
  OAI21OPTREPBD1BWP30P140 U103 ( .A1(n1), .A2(n41), .B(n40), .ZN(N325) );
  ND2OPTIBD4BWP30P140 U104 ( .A1(n87), .A2(i_data_bus[39]), .ZN(n42) );
  OAI21OPTREPBD1BWP30P140 U105 ( .A1(n1), .A2(n43), .B(n42), .ZN(N326) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[8]), .ZN(n45) );
  ND2OPTIBD4BWP30P140 U107 ( .A1(n87), .A2(i_data_bus[40]), .ZN(n44) );
  OAI21OPTREPBD1BWP30P140 U108 ( .A1(n1), .A2(n45), .B(n44), .ZN(N327) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[9]), .ZN(n47) );
  ND2OPTIBD4BWP30P140 U110 ( .A1(n87), .A2(i_data_bus[41]), .ZN(n46) );
  OAI21OPTREPBD1BWP30P140 U111 ( .A1(n1), .A2(n47), .B(n46), .ZN(N328) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[10]), .ZN(n49) );
  ND2OPTIBD4BWP30P140 U113 ( .A1(n87), .A2(i_data_bus[42]), .ZN(n48) );
  OAI21OPTREPBD1BWP30P140 U114 ( .A1(n1), .A2(n49), .B(n48), .ZN(N329) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[11]), .ZN(n51) );
  ND2OPTIBD4BWP30P140 U116 ( .A1(n87), .A2(i_data_bus[43]), .ZN(n50) );
  OAI21OPTREPBD1BWP30P140 U117 ( .A1(n1), .A2(n51), .B(n50), .ZN(N330) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[12]), .ZN(n53) );
  OAI21OPTREPBD1BWP30P140 U119 ( .A1(n1), .A2(n53), .B(n52), .ZN(N331) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[13]), .ZN(n55) );
  OAI21OPTREPBD1BWP30P140 U121 ( .A1(n1), .A2(n55), .B(n54), .ZN(N332) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[14]), .ZN(n57) );
  OAI21OPTREPBD1BWP30P140 U123 ( .A1(n1), .A2(n57), .B(n56), .ZN(N333) );
  INVD1BWP30P140 U124 ( .I(i_data_bus[15]), .ZN(n59) );
  INVD1BWP30P140 U125 ( .I(i_data_bus[16]), .ZN(n61) );
  INVD1BWP30P140 U126 ( .I(i_data_bus[17]), .ZN(n90) );
  ND2OPTIBD4BWP30P140 U127 ( .A1(n87), .A2(i_data_bus[49]), .ZN(n62) );
  INVD1BWP30P140 U128 ( .I(i_data_bus[18]), .ZN(n102) );
  ND2OPTIBD4BWP30P140 U129 ( .A1(n87), .A2(i_data_bus[50]), .ZN(n63) );
  INVD1BWP30P140 U130 ( .I(i_data_bus[19]), .ZN(n100) );
  ND2OPTIBD4BWP30P140 U131 ( .A1(n87), .A2(i_data_bus[51]), .ZN(n64) );
  INVD1BWP30P140 U132 ( .I(i_data_bus[20]), .ZN(n66) );
  ND2OPTIBD4BWP30P140 U133 ( .A1(n87), .A2(i_data_bus[52]), .ZN(n65) );
  INVD1BWP30P140 U134 ( .I(i_data_bus[21]), .ZN(n68) );
  INVD1BWP30P140 U135 ( .I(i_data_bus[22]), .ZN(n70) );
  INVD1BWP30P140 U136 ( .I(i_data_bus[23]), .ZN(n72) );
  ND2OPTIBD4BWP30P140 U137 ( .A1(n87), .A2(i_data_bus[55]), .ZN(n71) );
  INVD1BWP30P140 U138 ( .I(i_data_bus[24]), .ZN(n74) );
  ND2OPTIBD4BWP30P140 U139 ( .A1(n87), .A2(i_data_bus[56]), .ZN(n73) );
  INVD1BWP30P140 U140 ( .I(i_data_bus[25]), .ZN(n76) );
  ND2OPTIBD4BWP30P140 U141 ( .A1(n87), .A2(i_data_bus[57]), .ZN(n75) );
  INVD1BWP30P140 U142 ( .I(i_data_bus[26]), .ZN(n78) );
  ND2OPTIBD4BWP30P140 U143 ( .A1(n87), .A2(i_data_bus[58]), .ZN(n77) );
  INVD1BWP30P140 U144 ( .I(i_data_bus[27]), .ZN(n80) );
  ND2OPTIBD4BWP30P140 U145 ( .A1(n87), .A2(i_data_bus[59]), .ZN(n79) );
  INVD1BWP30P140 U146 ( .I(i_data_bus[28]), .ZN(n82) );
  ND2OPTIBD4BWP30P140 U147 ( .A1(n87), .A2(i_data_bus[60]), .ZN(n81) );
  INVD1BWP30P140 U148 ( .I(i_data_bus[2]), .ZN(n89) );
  INVD1BWP30P140 U149 ( .I(n93), .ZN(n95) );
  OAI21D1BWP30P140 U150 ( .A1(n95), .A2(i_cmd[1]), .B(n94), .ZN(N354) );
  OAI31D1BWP30P140 U151 ( .A1(n98), .A2(n97), .A3(n96), .B(n3), .ZN(N353) );
  INVD1BWP30P140 U152 ( .I(i_data_bus[51]), .ZN(n99) );
  OAI22D1BWP30P140 U153 ( .A1(n3), .A2(n100), .B1(n126), .B2(n99), .ZN(N306)
         );
  INVD1BWP30P140 U154 ( .I(i_data_bus[50]), .ZN(n101) );
  OAI22D1BWP30P140 U155 ( .A1(n3), .A2(n102), .B1(n126), .B2(n101), .ZN(N305)
         );
  INVD6BWP30P140 U156 ( .I(n103), .ZN(n130) );
  INVD1BWP30P140 U157 ( .I(i_data_bus[60]), .ZN(n105) );
  MOAI22D1BWP30P140 U158 ( .A1(n130), .A2(n105), .B1(n128), .B2(i_data_bus[28]), .ZN(N315) );
  BUFFD4BWP30P140 U159 ( .I(n126), .Z(n123) );
  INVD1BWP30P140 U160 ( .I(i_data_bus[48]), .ZN(n106) );
  MOAI22D1BWP30P140 U161 ( .A1(n123), .A2(n106), .B1(n128), .B2(i_data_bus[16]), .ZN(N303) );
  INVD1BWP30P140 U162 ( .I(i_data_bus[34]), .ZN(n107) );
  MOAI22D1BWP30P140 U163 ( .A1(n108), .A2(n107), .B1(n128), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140 U164 ( .I(i_data_bus[59]), .ZN(n109) );
  MOAI22D1BWP30P140 U165 ( .A1(n130), .A2(n109), .B1(n128), .B2(i_data_bus[27]), .ZN(N314) );
  INVD1BWP30P140 U166 ( .I(i_data_bus[47]), .ZN(n110) );
  MOAI22D1BWP30P140 U167 ( .A1(n123), .A2(n110), .B1(n128), .B2(i_data_bus[15]), .ZN(N302) );
  INVD1BWP30P140 U168 ( .I(i_data_bus[33]), .ZN(n111) );
  MOAI22D1BWP30P140 U169 ( .A1(n130), .A2(n111), .B1(n128), .B2(i_data_bus[1]), 
        .ZN(N288) );
  INVD1BWP30P140 U170 ( .I(i_data_bus[58]), .ZN(n112) );
  MOAI22D1BWP30P140 U171 ( .A1(n130), .A2(n112), .B1(n128), .B2(i_data_bus[26]), .ZN(N313) );
  INVD1BWP30P140 U172 ( .I(i_data_bus[46]), .ZN(n113) );
  MOAI22D1BWP30P140 U173 ( .A1(n123), .A2(n113), .B1(n128), .B2(i_data_bus[14]), .ZN(N301) );
  INVD1BWP30P140 U174 ( .I(i_data_bus[32]), .ZN(n114) );
  MOAI22D1BWP30P140 U175 ( .A1(n130), .A2(n114), .B1(n128), .B2(i_data_bus[0]), 
        .ZN(N287) );
  INVD1BWP30P140 U176 ( .I(i_data_bus[57]), .ZN(n115) );
  MOAI22D1BWP30P140 U177 ( .A1(n123), .A2(n115), .B1(n128), .B2(i_data_bus[25]), .ZN(N312) );
  INVD1BWP30P140 U178 ( .I(i_data_bus[45]), .ZN(n116) );
  MOAI22D1BWP30P140 U179 ( .A1(n123), .A2(n116), .B1(n128), .B2(i_data_bus[13]), .ZN(N300) );
  INVD1BWP30P140 U180 ( .I(i_data_bus[56]), .ZN(n117) );
  MOAI22D1BWP30P140 U181 ( .A1(n130), .A2(n117), .B1(n128), .B2(i_data_bus[24]), .ZN(N311) );
  INVD1BWP30P140 U182 ( .I(i_data_bus[44]), .ZN(n118) );
  MOAI22D1BWP30P140 U183 ( .A1(n123), .A2(n118), .B1(n128), .B2(i_data_bus[12]), .ZN(N299) );
  INVD1BWP30P140 U184 ( .I(i_data_bus[55]), .ZN(n119) );
  MOAI22D1BWP30P140 U185 ( .A1(n130), .A2(n119), .B1(n128), .B2(i_data_bus[23]), .ZN(N310) );
  INVD1BWP30P140 U186 ( .I(i_data_bus[43]), .ZN(n120) );
  MOAI22D1BWP30P140 U187 ( .A1(n123), .A2(n120), .B1(n128), .B2(i_data_bus[11]), .ZN(N298) );
  INVD1BWP30P140 U188 ( .I(i_data_bus[54]), .ZN(n121) );
  MOAI22D1BWP30P140 U189 ( .A1(n130), .A2(n121), .B1(n128), .B2(i_data_bus[22]), .ZN(N309) );
  INVD1BWP30P140 U190 ( .I(i_data_bus[42]), .ZN(n122) );
  MOAI22D1BWP30P140 U191 ( .A1(n123), .A2(n122), .B1(n128), .B2(i_data_bus[10]), .ZN(N297) );
  INVD1BWP30P140 U192 ( .I(i_data_bus[53]), .ZN(n124) );
  MOAI22D1BWP30P140 U193 ( .A1(n130), .A2(n124), .B1(n128), .B2(i_data_bus[21]), .ZN(N308) );
  INVD1BWP30P140 U194 ( .I(i_data_bus[41]), .ZN(n125) );
  INVD1BWP30P140 U195 ( .I(i_data_bus[52]), .ZN(n127) );
  MOAI22D1BWP30P140 U196 ( .A1(n130), .A2(n127), .B1(n128), .B2(i_data_bus[20]), .ZN(N307) );
  INVD1BWP30P140 U197 ( .I(i_data_bus[40]), .ZN(n129) );
  MOAI22D1BWP30P140 U198 ( .A1(n130), .A2(n129), .B1(n128), .B2(i_data_bus[8]), 
        .ZN(N295) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_138 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  ND2OPTIBD1BWP30P140 U3 ( .A1(n75), .A2(i_data_bus[57]), .ZN(n76) );
  ND2OPTPAD4BWP30P140 U4 ( .A1(n6), .A2(n5), .ZN(n126) );
  INVD4BWP30P140 U5 ( .I(n15), .ZN(n95) );
  NR2D3BWP30P140 U6 ( .A1(n95), .A2(n100), .ZN(n19) );
  IOA21D1BWP30P140 U7 ( .A1(n26), .A2(i_data_bus[6]), .B(n27), .ZN(N325) );
  INVD6BWP30P140 U8 ( .I(n26), .ZN(n81) );
  INVD6BWP30P140 U9 ( .I(n26), .ZN(n89) );
  OAI21D2BWP30P140 U10 ( .A1(n89), .A2(n79), .B(n78), .ZN(N347) );
  OAI21D2BWP30P140 U11 ( .A1(n81), .A2(n104), .B(n82), .ZN(N349) );
  OAI21D2BWP30P140 U12 ( .A1(n81), .A2(n91), .B(n83), .ZN(N350) );
  OAI21D2BWP30P140 U13 ( .A1(n89), .A2(n85), .B(n84), .ZN(N343) );
  OAI21D2BWP30P140 U14 ( .A1(n81), .A2(n88), .B(n87), .ZN(N342) );
  OAI21D2BWP30P140 U15 ( .A1(n81), .A2(n34), .B(n33), .ZN(N338) );
  OAI21D2BWP30P140 U16 ( .A1(n81), .A2(n36), .B(n35), .ZN(N336) );
  OAI21D2BWP30P140 U17 ( .A1(n81), .A2(n46), .B(n45), .ZN(N333) );
  OAI21D2BWP30P140 U18 ( .A1(n81), .A2(n50), .B(n49), .ZN(N331) );
  OAI21D2BWP30P140 U19 ( .A1(n89), .A2(n54), .B(n53), .ZN(N329) );
  OAI21D2BWP30P140 U20 ( .A1(n81), .A2(n58), .B(n57), .ZN(N327) );
  OAI21D2BWP30P140 U21 ( .A1(n81), .A2(n60), .B(n59), .ZN(N326) );
  OAI21D2BWP30P140 U22 ( .A1(n81), .A2(n62), .B(n61), .ZN(N324) );
  OAI21D2BWP30P140 U23 ( .A1(n81), .A2(n64), .B(n63), .ZN(N323) );
  OAI21D2BWP30P140 U24 ( .A1(n81), .A2(n66), .B(n65), .ZN(N322) );
  OAI21D2BWP30P140 U25 ( .A1(n81), .A2(n68), .B(n67), .ZN(N321) );
  OAI21D2BWP30P140 U26 ( .A1(n81), .A2(n70), .B(n69), .ZN(N320) );
  OAI21D2BWP30P140 U27 ( .A1(n81), .A2(n72), .B(n71), .ZN(N319) );
  OAI21D2BWP30P140 U28 ( .A1(n81), .A2(n74), .B(n73), .ZN(N337) );
  OAI21D2BWP30P140 U29 ( .A1(n81), .A2(n102), .B(n80), .ZN(N348) );
  INVD6BWP30P140 U30 ( .I(n96), .ZN(n75) );
  INVD2BWP30P140 U31 ( .I(i_valid[1]), .ZN(n16) );
  CKND2D2BWP30P140 U32 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n21) );
  BUFFD4BWP30P140 U33 ( .I(n126), .Z(n1) );
  INVD3BWP30P140 U34 ( .I(n2), .ZN(n94) );
  CKND2D3BWP30P140 U35 ( .A1(i_valid[0]), .A2(n22), .ZN(n2) );
  INVD1BWP30P140 U36 ( .I(i_cmd[0]), .ZN(n3) );
  NR2OPTPAD2BWP30P140 U37 ( .A1(n3), .A2(n100), .ZN(n6) );
  INVD4BWP30P140 U38 ( .I(i_cmd[1]), .ZN(n15) );
  ND2OPTIBD1BWP30P140 U39 ( .A1(n93), .A2(n92), .ZN(N318) );
  OR2D1BWP30P140 U40 ( .A1(n105), .A2(n91), .Z(n92) );
  ND2OPTIBD1BWP30P140 U41 ( .A1(n90), .A2(i_data_bus[63]), .ZN(n93) );
  ND2D1BWP30P140 U42 ( .A1(n75), .A2(i_data_bus[41]), .ZN(n55) );
  ND2D1BWP30P140 U43 ( .A1(n75), .A2(i_data_bus[43]), .ZN(n51) );
  ND2D1BWP30P140 U44 ( .A1(n75), .A2(i_data_bus[45]), .ZN(n47) );
  ND2D1BWP30P140 U45 ( .A1(n75), .A2(i_data_bus[47]), .ZN(n43) );
  ND2D1BWP30P140 U46 ( .A1(n75), .A2(i_data_bus[52]), .ZN(n37) );
  ND2D1BWP30P140 U47 ( .A1(n75), .A2(i_data_bus[53]), .ZN(n39) );
  ND2D1BWP30P140 U48 ( .A1(n75), .A2(i_data_bus[54]), .ZN(n41) );
  ND2D1BWP30P140 U49 ( .A1(n75), .A2(i_data_bus[59]), .ZN(n31) );
  INVD8BWP30P140 U50 ( .I(n90), .ZN(n129) );
  INVD4BWP30P140 U51 ( .I(n20), .ZN(n26) );
  INVD1BWP30P140 U52 ( .I(rst), .ZN(n4) );
  ND2D1BWP30P140 U53 ( .A1(n4), .A2(i_en), .ZN(n100) );
  INVD2BWP30P140 U54 ( .I(i_valid[1]), .ZN(n99) );
  INVD3BWP30P140 U55 ( .I(i_valid[0]), .ZN(n17) );
  MUX2NOPTD4BWP30P140 U56 ( .I0(n99), .I1(n17), .S(n15), .ZN(n5) );
  INVD4BWP30P140 U57 ( .I(n126), .ZN(n90) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[49]), .ZN(n7) );
  INVD1BWP30P140 U59 ( .I(n100), .ZN(n22) );
  INVD2BWP30P140 U60 ( .I(i_cmd[0]), .ZN(n98) );
  ND2OPTPAD8BWP30P140 U61 ( .A1(n94), .A2(n98), .ZN(n105) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[17]), .ZN(n36) );
  OAI22OPTPBD1BWP30P140 U63 ( .A1(n129), .A2(n7), .B1(n105), .B2(n36), .ZN(
        N304) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[50]), .ZN(n8) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[18]), .ZN(n74) );
  OAI22OPTPBD1BWP30P140 U66 ( .A1(n129), .A2(n8), .B1(n105), .B2(n74), .ZN(
        N305) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[51]), .ZN(n9) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[19]), .ZN(n34) );
  OAI22OPTPBD1BWP30P140 U69 ( .A1(n129), .A2(n9), .B1(n105), .B2(n34), .ZN(
        N306) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[39]), .ZN(n10) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[7]), .ZN(n60) );
  OAI22OPTPBD1BWP30P140 U72 ( .A1(n129), .A2(n10), .B1(n105), .B2(n60), .ZN(
        N294) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[38]), .ZN(n11) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[6]), .ZN(n28) );
  OAI22OPTPBD1BWP30P140 U75 ( .A1(n129), .A2(n11), .B1(n105), .B2(n28), .ZN(
        N293) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[37]), .ZN(n12) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[5]), .ZN(n62) );
  OAI22OPTPBD1BWP30P140 U78 ( .A1(n129), .A2(n12), .B1(n105), .B2(n62), .ZN(
        N292) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[36]), .ZN(n13) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[4]), .ZN(n64) );
  OAI22OPTPBD1BWP30P140 U81 ( .A1(n129), .A2(n13), .B1(n105), .B2(n64), .ZN(
        N291) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[35]), .ZN(n14) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[3]), .ZN(n66) );
  OAI22OPTPBD1BWP30P140 U84 ( .A1(n129), .A2(n14), .B1(n105), .B2(n66), .ZN(
        N290) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[16]), .ZN(n25) );
  MUX2NOPTD4BWP30P140 U86 ( .I0(n17), .I1(n16), .S(i_cmd[0]), .ZN(n18) );
  CKND2D4BWP30P140 U87 ( .A1(n19), .A2(n18), .ZN(n20) );
  INVD2BWP30P140 U88 ( .I(n21), .ZN(n23) );
  ND2OPTPAD4BWP30P140 U89 ( .A1(n23), .A2(n22), .ZN(n96) );
  ND2D1BWP30P140 U90 ( .A1(n75), .A2(i_data_bus[48]), .ZN(n24) );
  OAI21D1BWP30P140 U91 ( .A1(n25), .A2(n89), .B(n24), .ZN(N335) );
  ND2D1BWP30P140 U92 ( .A1(n75), .A2(i_data_bus[38]), .ZN(n27) );
  INVD1BWP30P140 U93 ( .I(i_data_bus[26]), .ZN(n30) );
  ND2D1BWP30P140 U94 ( .A1(n75), .A2(i_data_bus[58]), .ZN(n29) );
  OAI21D1BWP30P140 U95 ( .A1(n30), .A2(n89), .B(n29), .ZN(N345) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[27]), .ZN(n32) );
  OAI21D1BWP30P140 U97 ( .A1(n32), .A2(n89), .B(n31), .ZN(N346) );
  INVD12BWP30P140 U98 ( .I(n96), .ZN(n86) );
  ND2OPTIBD4BWP30P140 U99 ( .A1(n86), .A2(i_data_bus[51]), .ZN(n33) );
  ND2OPTIBD4BWP30P140 U100 ( .A1(n86), .A2(i_data_bus[49]), .ZN(n35) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[20]), .ZN(n38) );
  OAI21D1BWP30P140 U102 ( .A1(n89), .A2(n38), .B(n37), .ZN(N339) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[21]), .ZN(n40) );
  OAI21D1BWP30P140 U104 ( .A1(n89), .A2(n40), .B(n39), .ZN(N340) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[22]), .ZN(n42) );
  OAI21D1BWP30P140 U106 ( .A1(n89), .A2(n42), .B(n41), .ZN(N341) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[15]), .ZN(n44) );
  OAI21D1BWP30P140 U108 ( .A1(n89), .A2(n44), .B(n43), .ZN(N334) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[14]), .ZN(n46) );
  ND2OPTIBD4BWP30P140 U110 ( .A1(n86), .A2(i_data_bus[46]), .ZN(n45) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[13]), .ZN(n48) );
  OAI21D1BWP30P140 U112 ( .A1(n89), .A2(n48), .B(n47), .ZN(N332) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[12]), .ZN(n50) );
  ND2OPTIBD4BWP30P140 U114 ( .A1(n86), .A2(i_data_bus[44]), .ZN(n49) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[11]), .ZN(n52) );
  OAI21D1BWP30P140 U116 ( .A1(n89), .A2(n52), .B(n51), .ZN(N330) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[10]), .ZN(n54) );
  ND2OPTIBD4BWP30P140 U118 ( .A1(n86), .A2(i_data_bus[42]), .ZN(n53) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[9]), .ZN(n56) );
  OAI21D1BWP30P140 U120 ( .A1(n89), .A2(n56), .B(n55), .ZN(N328) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[8]), .ZN(n58) );
  ND2OPTIBD4BWP30P140 U122 ( .A1(n86), .A2(i_data_bus[40]), .ZN(n57) );
  ND2OPTIBD4BWP30P140 U123 ( .A1(n86), .A2(i_data_bus[39]), .ZN(n59) );
  ND2OPTIBD4BWP30P140 U124 ( .A1(n86), .A2(i_data_bus[37]), .ZN(n61) );
  ND2OPTIBD4BWP30P140 U125 ( .A1(n86), .A2(i_data_bus[36]), .ZN(n63) );
  ND2OPTIBD4BWP30P140 U126 ( .A1(n86), .A2(i_data_bus[35]), .ZN(n65) );
  INVD1BWP30P140 U127 ( .I(i_data_bus[2]), .ZN(n68) );
  ND2OPTIBD4BWP30P140 U128 ( .A1(n86), .A2(i_data_bus[34]), .ZN(n67) );
  INVD1BWP30P140 U129 ( .I(i_data_bus[1]), .ZN(n70) );
  ND2OPTIBD4BWP30P140 U130 ( .A1(n86), .A2(i_data_bus[33]), .ZN(n69) );
  INVD1BWP30P140 U131 ( .I(i_data_bus[0]), .ZN(n72) );
  ND2OPTIBD4BWP30P140 U132 ( .A1(n86), .A2(i_data_bus[32]), .ZN(n71) );
  ND2OPTIBD4BWP30P140 U133 ( .A1(n86), .A2(i_data_bus[50]), .ZN(n73) );
  INVD1BWP30P140 U134 ( .I(i_data_bus[25]), .ZN(n77) );
  OAI21D1BWP30P140 U135 ( .A1(n89), .A2(n77), .B(n76), .ZN(N344) );
  INVD1BWP30P140 U136 ( .I(i_data_bus[28]), .ZN(n79) );
  ND2OPTIBD4BWP30P140 U137 ( .A1(n86), .A2(i_data_bus[60]), .ZN(n78) );
  INVD1BWP30P140 U138 ( .I(i_data_bus[29]), .ZN(n102) );
  ND2OPTIBD4BWP30P140 U139 ( .A1(n86), .A2(i_data_bus[61]), .ZN(n80) );
  INVD1BWP30P140 U140 ( .I(i_data_bus[30]), .ZN(n104) );
  ND2OPTIBD4BWP30P140 U141 ( .A1(n86), .A2(i_data_bus[62]), .ZN(n82) );
  INVD1BWP30P140 U142 ( .I(i_data_bus[31]), .ZN(n91) );
  ND2OPTIBD4BWP30P140 U143 ( .A1(n86), .A2(i_data_bus[63]), .ZN(n83) );
  INVD1BWP30P140 U144 ( .I(i_data_bus[24]), .ZN(n85) );
  ND2OPTIBD4BWP30P140 U145 ( .A1(n86), .A2(i_data_bus[56]), .ZN(n84) );
  INVD1BWP30P140 U146 ( .I(i_data_bus[23]), .ZN(n88) );
  ND2OPTIBD4BWP30P140 U147 ( .A1(n86), .A2(i_data_bus[55]), .ZN(n87) );
  INVD1BWP30P140 U148 ( .I(n94), .ZN(n97) );
  OAI21D1BWP30P140 U149 ( .A1(n97), .A2(n95), .B(n96), .ZN(N354) );
  OAI31D1BWP30P140 U150 ( .A1(n100), .A2(n99), .A3(n98), .B(n105), .ZN(N353)
         );
  INVD1BWP30P140 U151 ( .I(i_data_bus[61]), .ZN(n101) );
  OAI22D1BWP30P140 U152 ( .A1(n105), .A2(n102), .B1(n126), .B2(n101), .ZN(N316) );
  INVD1BWP30P140 U153 ( .I(i_data_bus[62]), .ZN(n103) );
  OAI22D1BWP30P140 U154 ( .A1(n105), .A2(n104), .B1(n126), .B2(n103), .ZN(N317) );
  INVD1BWP30P140 U155 ( .I(i_data_bus[60]), .ZN(n106) );
  INVD8BWP30P140 U156 ( .I(n105), .ZN(n127) );
  MOAI22D1BWP30P140 U157 ( .A1(n1), .A2(n106), .B1(n127), .B2(i_data_bus[28]), 
        .ZN(N315) );
  INVD1BWP30P140 U158 ( .I(i_data_bus[48]), .ZN(n107) );
  MOAI22D1BWP30P140 U159 ( .A1(n129), .A2(n107), .B1(n127), .B2(i_data_bus[16]), .ZN(N303) );
  INVD1BWP30P140 U160 ( .I(i_data_bus[34]), .ZN(n108) );
  MOAI22D1BWP30P140 U161 ( .A1(n129), .A2(n108), .B1(n127), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140 U162 ( .I(i_data_bus[59]), .ZN(n109) );
  MOAI22D1BWP30P140 U163 ( .A1(n1), .A2(n109), .B1(n127), .B2(i_data_bus[27]), 
        .ZN(N314) );
  INVD1BWP30P140 U164 ( .I(i_data_bus[47]), .ZN(n110) );
  MOAI22D1BWP30P140 U165 ( .A1(n129), .A2(n110), .B1(n127), .B2(i_data_bus[15]), .ZN(N302) );
  INVD1BWP30P140 U166 ( .I(i_data_bus[33]), .ZN(n111) );
  MOAI22D1BWP30P140 U167 ( .A1(n129), .A2(n111), .B1(n127), .B2(i_data_bus[1]), 
        .ZN(N288) );
  INVD1BWP30P140 U168 ( .I(i_data_bus[58]), .ZN(n112) );
  MOAI22D1BWP30P140 U169 ( .A1(n1), .A2(n112), .B1(n127), .B2(i_data_bus[26]), 
        .ZN(N313) );
  INVD1BWP30P140 U170 ( .I(i_data_bus[46]), .ZN(n113) );
  MOAI22D1BWP30P140 U171 ( .A1(n129), .A2(n113), .B1(n127), .B2(i_data_bus[14]), .ZN(N301) );
  INVD1BWP30P140 U172 ( .I(i_data_bus[32]), .ZN(n114) );
  MOAI22D1BWP30P140 U173 ( .A1(n129), .A2(n114), .B1(n127), .B2(i_data_bus[0]), 
        .ZN(N287) );
  INVD1BWP30P140 U174 ( .I(i_data_bus[57]), .ZN(n115) );
  MOAI22D1BWP30P140 U175 ( .A1(n1), .A2(n115), .B1(n127), .B2(i_data_bus[25]), 
        .ZN(N312) );
  INVD1BWP30P140 U176 ( .I(i_data_bus[45]), .ZN(n116) );
  MOAI22D1BWP30P140 U177 ( .A1(n129), .A2(n116), .B1(n127), .B2(i_data_bus[13]), .ZN(N300) );
  INVD1BWP30P140 U178 ( .I(i_data_bus[56]), .ZN(n117) );
  MOAI22D1BWP30P140 U179 ( .A1(n1), .A2(n117), .B1(n127), .B2(i_data_bus[24]), 
        .ZN(N311) );
  INVD1BWP30P140 U180 ( .I(i_data_bus[44]), .ZN(n118) );
  MOAI22D1BWP30P140 U181 ( .A1(n129), .A2(n118), .B1(n127), .B2(i_data_bus[12]), .ZN(N299) );
  INVD1BWP30P140 U182 ( .I(i_data_bus[55]), .ZN(n119) );
  MOAI22D1BWP30P140 U183 ( .A1(n1), .A2(n119), .B1(n127), .B2(i_data_bus[23]), 
        .ZN(N310) );
  INVD1BWP30P140 U184 ( .I(i_data_bus[43]), .ZN(n120) );
  MOAI22D1BWP30P140 U185 ( .A1(n129), .A2(n120), .B1(n127), .B2(i_data_bus[11]), .ZN(N298) );
  INVD1BWP30P140 U186 ( .I(i_data_bus[54]), .ZN(n121) );
  MOAI22D1BWP30P140 U187 ( .A1(n1), .A2(n121), .B1(n127), .B2(i_data_bus[22]), 
        .ZN(N309) );
  INVD1BWP30P140 U188 ( .I(i_data_bus[42]), .ZN(n122) );
  MOAI22D1BWP30P140 U189 ( .A1(n129), .A2(n122), .B1(n127), .B2(i_data_bus[10]), .ZN(N297) );
  INVD1BWP30P140 U190 ( .I(i_data_bus[53]), .ZN(n123) );
  MOAI22D1BWP30P140 U191 ( .A1(n1), .A2(n123), .B1(n127), .B2(i_data_bus[21]), 
        .ZN(N308) );
  INVD1BWP30P140 U192 ( .I(i_data_bus[41]), .ZN(n124) );
  MOAI22D1BWP30P140 U193 ( .A1(n129), .A2(n124), .B1(n127), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140 U194 ( .I(i_data_bus[52]), .ZN(n125) );
  MOAI22D1BWP30P140 U195 ( .A1(n1), .A2(n125), .B1(n127), .B2(i_data_bus[20]), 
        .ZN(N307) );
  INVD1BWP30P140 U196 ( .I(i_data_bus[40]), .ZN(n128) );
  MOAI22D1BWP30P140 U197 ( .A1(n129), .A2(n128), .B1(n127), .B2(i_data_bus[8]), 
        .ZN(N295) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_139 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI21D1BWP30P140 U3 ( .A1(n89), .A2(n33), .B(n32), .ZN(N323) );
  OAI21D1BWP30P140 U4 ( .A1(n89), .A2(n37), .B(n36), .ZN(N326) );
  CKND2D2BWP30P140 U5 ( .A1(n66), .A2(i_data_bus[57]), .ZN(n53) );
  ND2D2BWP30P140 U6 ( .A1(n66), .A2(i_data_bus[61]), .ZN(n61) );
  ND2D2BWP30P140 U7 ( .A1(n66), .A2(i_data_bus[63]), .ZN(n67) );
  CKND2D2BWP30P140 U8 ( .A1(n66), .A2(i_data_bus[33]), .ZN(n24) );
  CKND2D2BWP30P140 U9 ( .A1(n66), .A2(i_data_bus[34]), .ZN(n26) );
  CKND2D2BWP30P140 U10 ( .A1(n66), .A2(i_data_bus[42]), .ZN(n43) );
  CKND2D2BWP30P140 U11 ( .A1(n66), .A2(i_data_bus[53]), .ZN(n45) );
  CKND2D2BWP30P140 U12 ( .A1(n66), .A2(i_data_bus[59]), .ZN(n57) );
  ND2OPTIBD1BWP30P140 U13 ( .A1(n63), .A2(i_data_bus[40]), .ZN(n38) );
  ND2OPTPAD6BWP30P140 U14 ( .A1(n71), .A2(n74), .ZN(n92) );
  INVD3BWP30P140 U15 ( .I(n15), .ZN(n18) );
  INVD6BWP30P140 U16 ( .I(n117), .ZN(n91) );
  CKND2D4BWP30P140 U17 ( .A1(n72), .A2(n14), .ZN(n15) );
  INVD6BWP30P140 U18 ( .I(n19), .ZN(n40) );
  INVD9BWP30P140 U19 ( .I(n79), .ZN(n63) );
  OAI21D1BWP30P140 U20 ( .A1(n89), .A2(n46), .B(n45), .ZN(N340) );
  OAI21D1BWP30P140 U21 ( .A1(n89), .A2(n58), .B(n57), .ZN(N346) );
  ND2OPTPAD4BWP30P140 U22 ( .A1(n5), .A2(n4), .ZN(n117) );
  INVD12BWP30P140 U23 ( .I(n40), .ZN(n89) );
  ND2OPTIBD1BWP30P140 U24 ( .A1(n63), .A2(i_data_bus[38]), .ZN(n34) );
  ND2OPTIBD1BWP30P140 U25 ( .A1(n63), .A2(i_data_bus[35]), .ZN(n22) );
  ND2OPTIBD1BWP30P140 U26 ( .A1(n63), .A2(i_data_bus[60]), .ZN(n59) );
  ND2OPTIBD1BWP30P140 U27 ( .A1(n63), .A2(i_data_bus[58]), .ZN(n55) );
  ND2OPTIBD1BWP30P140 U28 ( .A1(n63), .A2(i_data_bus[56]), .ZN(n51) );
  ND2OPTIBD1BWP30P140 U29 ( .A1(n63), .A2(i_data_bus[54]), .ZN(n47) );
  ND2OPTIBD1BWP30P140 U30 ( .A1(n63), .A2(i_data_bus[41]), .ZN(n41) );
  ND2OPTIBD1BWP30P140 U31 ( .A1(n63), .A2(i_data_bus[62]), .ZN(n64) );
  INVD3BWP30P140 U32 ( .I(i_cmd[0]), .ZN(n74) );
  BUFFD4BWP30P140 U33 ( .I(n117), .Z(n1) );
  ND2OPTPAD4BWP30P140 U34 ( .A1(n18), .A2(n17), .ZN(n19) );
  INVD3BWP30P140 U35 ( .I(n2), .ZN(n71) );
  CKND2D3BWP30P140 U36 ( .A1(i_valid[0]), .A2(n14), .ZN(n2) );
  INVD6BWP30P140 U37 ( .I(n91), .ZN(n96) );
  ND2OPTPAD2BWP30P140 U38 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n20) );
  INVD6BWP30P140 U39 ( .I(n79), .ZN(n66) );
  MUX2NOPTD4BWP30P140 U40 ( .I0(n16), .I1(n75), .S(i_cmd[0]), .ZN(n17) );
  CKND2D3BWP30P140 U41 ( .A1(n66), .A2(i_data_bus[37]), .ZN(n28) );
  OAI21D2BWP30P140 U42 ( .A1(n89), .A2(n29), .B(n28), .ZN(N324) );
  CKND2D3BWP30P140 U43 ( .A1(n66), .A2(i_data_bus[36]), .ZN(n32) );
  CKND2D3BWP30P140 U44 ( .A1(n66), .A2(i_data_bus[39]), .ZN(n36) );
  CKND2D3BWP30P140 U45 ( .A1(n66), .A2(i_data_bus[55]), .ZN(n49) );
  OAI21D2BWP30P140 U46 ( .A1(n89), .A2(n50), .B(n49), .ZN(N342) );
  OAI21D2BWP30P140 U47 ( .A1(n89), .A2(n54), .B(n53), .ZN(N344) );
  OAI21D2BWP30P140 U48 ( .A1(n89), .A2(n62), .B(n61), .ZN(N348) );
  OAI21D2BWP30P140 U49 ( .A1(n89), .A2(n68), .B(n67), .ZN(N350) );
  OAI21D2BWP30P140 U50 ( .A1(n89), .A2(n25), .B(n24), .ZN(N320) );
  OAI21D2BWP30P140 U51 ( .A1(n89), .A2(n27), .B(n26), .ZN(N321) );
  ND2OPTIBD1BWP30P140 U52 ( .A1(n63), .A2(i_data_bus[32]), .ZN(n30) );
  OAI21D2BWP30P140 U53 ( .A1(n89), .A2(n31), .B(n30), .ZN(N319) );
  OAI21D2BWP30P140 U54 ( .A1(n89), .A2(n39), .B(n38), .ZN(N327) );
  OAI21D2BWP30P140 U55 ( .A1(n89), .A2(n44), .B(n43), .ZN(N329) );
  ND2OPTIBD1BWP30P140 U56 ( .A1(n70), .A2(n69), .ZN(N304) );
  OR2D1BWP30P140 U57 ( .A1(n92), .A2(n86), .Z(n69) );
  ND2OPTIBD1BWP30P140 U58 ( .A1(n91), .A2(i_data_bus[49]), .ZN(n70) );
  INVD1BWP30P140 U59 ( .I(n76), .ZN(n14) );
  INVD1BWP30P140 U60 ( .I(rst), .ZN(n3) );
  ND2D1BWP30P140 U61 ( .A1(n3), .A2(i_en), .ZN(n76) );
  INR2D4BWP30P140 U62 ( .A1(i_cmd[0]), .B1(n76), .ZN(n5) );
  INVD2BWP30P140 U63 ( .I(i_valid[0]), .ZN(n16) );
  INVD4BWP30P140 U64 ( .I(i_valid[1]), .ZN(n75) );
  MUX2NOPTD4BWP30P140 U65 ( .I0(n16), .I1(n75), .S(i_cmd[1]), .ZN(n4) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[63]), .ZN(n6) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[31]), .ZN(n68) );
  OAI22OPTPBD1BWP30P140 U68 ( .A1(n96), .A2(n6), .B1(n92), .B2(n68), .ZN(N318)
         );
  INVD1BWP30P140 U69 ( .I(i_data_bus[62]), .ZN(n7) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[30]), .ZN(n65) );
  OAI22OPTPBD1BWP30P140 U71 ( .A1(n96), .A2(n7), .B1(n92), .B2(n65), .ZN(N317)
         );
  INVD1BWP30P140 U72 ( .I(i_data_bus[61]), .ZN(n8) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[29]), .ZN(n62) );
  OAI22OPTPBD1BWP30P140 U74 ( .A1(n96), .A2(n8), .B1(n92), .B2(n62), .ZN(N316)
         );
  INVD1BWP30P140 U75 ( .I(i_data_bus[35]), .ZN(n9) );
  INVD1BWP30P140 U76 ( .I(i_data_bus[3]), .ZN(n23) );
  OAI22OPTPBD1BWP30P140 U77 ( .A1(n96), .A2(n9), .B1(n92), .B2(n23), .ZN(N290)
         );
  INVD1BWP30P140 U78 ( .I(i_data_bus[36]), .ZN(n10) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[4]), .ZN(n33) );
  OAI22OPTPBD1BWP30P140 U80 ( .A1(n96), .A2(n10), .B1(n92), .B2(n33), .ZN(N291) );
  INVD1BWP30P140 U81 ( .I(i_data_bus[38]), .ZN(n11) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[6]), .ZN(n35) );
  OAI22OPTPBD1BWP30P140 U83 ( .A1(n96), .A2(n11), .B1(n92), .B2(n35), .ZN(N293) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[39]), .ZN(n12) );
  INVD1BWP30P140 U85 ( .I(i_data_bus[7]), .ZN(n37) );
  OAI22OPTPBD1BWP30P140 U86 ( .A1(n96), .A2(n12), .B1(n92), .B2(n37), .ZN(N294) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[37]), .ZN(n13) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[5]), .ZN(n29) );
  OAI22OPTPBD1BWP30P140 U89 ( .A1(n96), .A2(n13), .B1(n92), .B2(n29), .ZN(N292) );
  INVD2BWP30P140 U90 ( .I(i_cmd[1]), .ZN(n72) );
  INVD3BWP30P140 U91 ( .I(n20), .ZN(n21) );
  ND2OPTPAD6BWP30P140 U92 ( .A1(n21), .A2(n14), .ZN(n79) );
  OAI21D1BWP30P140 U93 ( .A1(n89), .A2(n23), .B(n22), .ZN(N322) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[1]), .ZN(n25) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[2]), .ZN(n27) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[0]), .ZN(n31) );
  OAI21D1BWP30P140 U97 ( .A1(n89), .A2(n35), .B(n34), .ZN(N325) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[8]), .ZN(n39) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[9]), .ZN(n42) );
  OAI21D1BWP30P140 U100 ( .A1(n89), .A2(n42), .B(n41), .ZN(N328) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[10]), .ZN(n44) );
  INVD1BWP30P140 U102 ( .I(i_data_bus[21]), .ZN(n46) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[22]), .ZN(n48) );
  OAI21D1BWP30P140 U104 ( .A1(n89), .A2(n48), .B(n47), .ZN(N341) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[23]), .ZN(n50) );
  INVD1BWP30P140 U106 ( .I(i_data_bus[24]), .ZN(n52) );
  OAI21D1BWP30P140 U107 ( .A1(n89), .A2(n52), .B(n51), .ZN(N343) );
  INVD1BWP30P140 U108 ( .I(i_data_bus[25]), .ZN(n54) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[26]), .ZN(n56) );
  OAI21D1BWP30P140 U110 ( .A1(n89), .A2(n56), .B(n55), .ZN(N345) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[27]), .ZN(n58) );
  INVD1BWP30P140 U112 ( .I(i_data_bus[28]), .ZN(n60) );
  OAI21D1BWP30P140 U113 ( .A1(n89), .A2(n60), .B(n59), .ZN(N347) );
  OAI21D1BWP30P140 U114 ( .A1(n89), .A2(n65), .B(n64), .ZN(N349) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[17]), .ZN(n86) );
  INVD1BWP30P140 U116 ( .I(n71), .ZN(n73) );
  OAI21D1BWP30P140 U117 ( .A1(n73), .A2(i_cmd[1]), .B(n79), .ZN(N354) );
  OAI31D1BWP30P140 U118 ( .A1(n76), .A2(n75), .A3(n74), .B(n92), .ZN(N353) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[19]), .ZN(n88) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[51]), .ZN(n77) );
  OAI22D1BWP30P140 U121 ( .A1(n92), .A2(n88), .B1(n117), .B2(n77), .ZN(N306)
         );
  INVD1BWP30P140 U122 ( .I(i_data_bus[18]), .ZN(n87) );
  INVD1BWP30P140 U123 ( .I(i_data_bus[50]), .ZN(n78) );
  OAI22D1BWP30P140 U124 ( .A1(n92), .A2(n87), .B1(n117), .B2(n78), .ZN(N305)
         );
  INVD1BWP30P140 U125 ( .I(i_data_bus[11]), .ZN(n80) );
  MOAI22D1BWP30P140 U126 ( .A1(n80), .A2(n89), .B1(i_data_bus[43]), .B2(n63), 
        .ZN(N330) );
  INVD1BWP30P140 U127 ( .I(i_data_bus[12]), .ZN(n81) );
  MOAI22D1BWP30P140 U128 ( .A1(n81), .A2(n89), .B1(i_data_bus[44]), .B2(n63), 
        .ZN(N331) );
  INVD1BWP30P140 U129 ( .I(i_data_bus[13]), .ZN(n82) );
  MOAI22D1BWP30P140 U130 ( .A1(n82), .A2(n89), .B1(i_data_bus[45]), .B2(n63), 
        .ZN(N332) );
  INVD1BWP30P140 U131 ( .I(i_data_bus[14]), .ZN(n83) );
  MOAI22D1BWP30P140 U132 ( .A1(n83), .A2(n89), .B1(i_data_bus[46]), .B2(n63), 
        .ZN(N333) );
  INVD1BWP30P140 U133 ( .I(i_data_bus[15]), .ZN(n84) );
  MOAI22D1BWP30P140 U134 ( .A1(n84), .A2(n89), .B1(i_data_bus[47]), .B2(n63), 
        .ZN(N334) );
  INVD1BWP30P140 U135 ( .I(i_data_bus[16]), .ZN(n85) );
  MOAI22D1BWP30P140 U136 ( .A1(n85), .A2(n89), .B1(i_data_bus[48]), .B2(n63), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U137 ( .A1(n86), .A2(n89), .B1(i_data_bus[49]), .B2(n63), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U138 ( .A1(n87), .A2(n89), .B1(i_data_bus[50]), .B2(n63), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U139 ( .A1(n88), .A2(n89), .B1(i_data_bus[51]), .B2(n63), 
        .ZN(N338) );
  INVD1BWP30P140 U140 ( .I(i_data_bus[20]), .ZN(n90) );
  MOAI22D1BWP30P140 U141 ( .A1(n90), .A2(n89), .B1(i_data_bus[52]), .B2(n63), 
        .ZN(N339) );
  INVD6BWP30P140 U142 ( .I(n91), .ZN(n114) );
  INVD1BWP30P140 U143 ( .I(i_data_bus[60]), .ZN(n93) );
  INVD8BWP30P140 U144 ( .I(n92), .ZN(n115) );
  MOAI22D1BWP30P140 U145 ( .A1(n114), .A2(n93), .B1(n115), .B2(i_data_bus[28]), 
        .ZN(N315) );
  INVD1BWP30P140 U146 ( .I(i_data_bus[48]), .ZN(n94) );
  MOAI22D1BWP30P140 U147 ( .A1(n1), .A2(n94), .B1(n115), .B2(i_data_bus[16]), 
        .ZN(N303) );
  INVD1BWP30P140 U148 ( .I(i_data_bus[34]), .ZN(n95) );
  MOAI22D1BWP30P140 U149 ( .A1(n114), .A2(n95), .B1(n115), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140 U150 ( .I(i_data_bus[59]), .ZN(n97) );
  MOAI22D1BWP30P140 U151 ( .A1(n96), .A2(n97), .B1(n115), .B2(i_data_bus[27]), 
        .ZN(N314) );
  INVD1BWP30P140 U152 ( .I(i_data_bus[47]), .ZN(n98) );
  MOAI22D1BWP30P140 U153 ( .A1(n1), .A2(n98), .B1(n115), .B2(i_data_bus[15]), 
        .ZN(N302) );
  INVD1BWP30P140 U154 ( .I(i_data_bus[33]), .ZN(n99) );
  MOAI22D1BWP30P140 U155 ( .A1(n114), .A2(n99), .B1(n115), .B2(i_data_bus[1]), 
        .ZN(N288) );
  INVD1BWP30P140 U156 ( .I(i_data_bus[58]), .ZN(n100) );
  MOAI22D1BWP30P140 U157 ( .A1(n114), .A2(n100), .B1(n115), .B2(i_data_bus[26]), .ZN(N313) );
  INVD1BWP30P140 U158 ( .I(i_data_bus[46]), .ZN(n101) );
  MOAI22D1BWP30P140 U159 ( .A1(n1), .A2(n101), .B1(n115), .B2(i_data_bus[14]), 
        .ZN(N301) );
  INVD1BWP30P140 U160 ( .I(i_data_bus[32]), .ZN(n102) );
  MOAI22D1BWP30P140 U161 ( .A1(n114), .A2(n102), .B1(n115), .B2(i_data_bus[0]), 
        .ZN(N287) );
  INVD1BWP30P140 U162 ( .I(i_data_bus[57]), .ZN(n103) );
  MOAI22D1BWP30P140 U163 ( .A1(n114), .A2(n103), .B1(n115), .B2(i_data_bus[25]), .ZN(N312) );
  INVD1BWP30P140 U164 ( .I(i_data_bus[45]), .ZN(n104) );
  MOAI22D1BWP30P140 U165 ( .A1(n1), .A2(n104), .B1(n115), .B2(i_data_bus[13]), 
        .ZN(N300) );
  INVD1BWP30P140 U166 ( .I(i_data_bus[56]), .ZN(n105) );
  MOAI22D1BWP30P140 U167 ( .A1(n114), .A2(n105), .B1(n115), .B2(i_data_bus[24]), .ZN(N311) );
  INVD1BWP30P140 U168 ( .I(i_data_bus[44]), .ZN(n106) );
  MOAI22D1BWP30P140 U169 ( .A1(n1), .A2(n106), .B1(n115), .B2(i_data_bus[12]), 
        .ZN(N299) );
  INVD1BWP30P140 U170 ( .I(i_data_bus[55]), .ZN(n107) );
  MOAI22D1BWP30P140 U171 ( .A1(n114), .A2(n107), .B1(n115), .B2(i_data_bus[23]), .ZN(N310) );
  INVD1BWP30P140 U172 ( .I(i_data_bus[43]), .ZN(n108) );
  MOAI22D1BWP30P140 U173 ( .A1(n1), .A2(n108), .B1(n115), .B2(i_data_bus[11]), 
        .ZN(N298) );
  INVD1BWP30P140 U174 ( .I(i_data_bus[54]), .ZN(n109) );
  MOAI22D1BWP30P140 U175 ( .A1(n114), .A2(n109), .B1(n115), .B2(i_data_bus[22]), .ZN(N309) );
  INVD1BWP30P140 U176 ( .I(i_data_bus[42]), .ZN(n110) );
  MOAI22D1BWP30P140 U177 ( .A1(n1), .A2(n110), .B1(n115), .B2(i_data_bus[10]), 
        .ZN(N297) );
  INVD1BWP30P140 U178 ( .I(i_data_bus[53]), .ZN(n111) );
  MOAI22D1BWP30P140 U179 ( .A1(n114), .A2(n111), .B1(n115), .B2(i_data_bus[21]), .ZN(N308) );
  INVD1BWP30P140 U180 ( .I(i_data_bus[41]), .ZN(n112) );
  MOAI22D1BWP30P140 U181 ( .A1(n1), .A2(n112), .B1(n115), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140 U182 ( .I(i_data_bus[52]), .ZN(n113) );
  MOAI22D1BWP30P140 U183 ( .A1(n114), .A2(n113), .B1(n115), .B2(i_data_bus[20]), .ZN(N307) );
  INVD1BWP30P140 U184 ( .I(i_data_bus[40]), .ZN(n116) );
  MOAI22D1BWP30P140 U185 ( .A1(n1), .A2(n116), .B1(n115), .B2(i_data_bus[8]), 
        .ZN(N295) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_140 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1P5BWP30P140 U3 ( .A1(n2), .A2(n13), .B1(n47), .B2(n74), .ZN(N305) );
  OAI22D1P5BWP30P140 U4 ( .A1(n2), .A2(n21), .B1(n47), .B2(n59), .ZN(N290) );
  INVD6BWP30P140 U5 ( .I(n55), .ZN(n86) );
  BUFFD6BWP30P140 U6 ( .I(n17), .Z(n27) );
  INR2D8BWP30P140 U7 ( .A1(i_valid[1]), .B1(n32), .ZN(n85) );
  INVD2BWP30P140 U8 ( .I(i_cmd[0]), .ZN(n11) );
  CKND2D2BWP30P140 U9 ( .A1(i_cmd[0]), .A2(n4), .ZN(n7) );
  INVD8BWP30P140 U10 ( .I(n101), .ZN(n1) );
  INVD15BWP30P140 U11 ( .I(n1), .ZN(n2) );
  IND2D1BWP30P140 U12 ( .A1(n48), .B1(n47), .ZN(N353) );
  INVD4BWP30P140 U13 ( .I(i_cmd[1]), .ZN(n5) );
  NR2D4BWP30P140 U14 ( .A1(n5), .A2(i_valid[1]), .ZN(n6) );
  OAI22OPTPBD2BWP30P140 U15 ( .A1(n2), .A2(n22), .B1(n27), .B2(n60), .ZN(N291)
         );
  OAI22OPTPBD2BWP30P140 U16 ( .A1(n2), .A2(n23), .B1(n27), .B2(n61), .ZN(N292)
         );
  OAI22OPTPBD2BWP30P140 U17 ( .A1(n2), .A2(n24), .B1(n27), .B2(n62), .ZN(N293)
         );
  OAI22OPTPBD2BWP30P140 U18 ( .A1(n2), .A2(n25), .B1(n27), .B2(n63), .ZN(N294)
         );
  OAI22OPTPBD2BWP30P140 U19 ( .A1(n2), .A2(n26), .B1(n27), .B2(n73), .ZN(N304)
         );
  OAI22OPTPBD2BWP30P140 U20 ( .A1(n2), .A2(n28), .B1(n27), .B2(n30), .ZN(N306)
         );
  INVD1BWP30P140 U21 ( .I(n43), .ZN(n45) );
  NR2OPTPAD2BWP30P140 U22 ( .A1(n7), .A2(n6), .ZN(n10) );
  NR3D0BWP30P140 U23 ( .A1(n46), .A2(n45), .A3(n44), .ZN(n48) );
  INVD2BWP30P140 U24 ( .I(n8), .ZN(n9) );
  ND2OPTPAD4BWP30P140 U25 ( .A1(n12), .A2(n11), .ZN(n17) );
  INVD4BWP30P140 U26 ( .I(n17), .ZN(n107) );
  CKND2D4BWP30P140 U27 ( .A1(i_valid[0]), .A2(n4), .ZN(n35) );
  ND2D1BWP30P140 U28 ( .A1(n16), .A2(n15), .ZN(N295) );
  OR2D1BWP30P140 U29 ( .A1(n101), .A2(n14), .Z(n16) );
  ND2D1BWP30P140 U30 ( .A1(n107), .A2(i_data_bus[8]), .ZN(n15) );
  INVD1BWP30P140 U31 ( .I(i_data_bus[40]), .ZN(n14) );
  ND2D1BWP30P140 U32 ( .A1(n34), .A2(n33), .ZN(N338) );
  ND2D1BWP30P140 U33 ( .A1(n85), .A2(i_data_bus[51]), .ZN(n33) );
  IND2D1BWP30P140 U34 ( .A1(n54), .B1(n31), .ZN(n34) );
  INR2D1BWP30P140 U35 ( .A1(i_data_bus[19]), .B1(n53), .ZN(n31) );
  ND2D1BWP30P140 U36 ( .A1(n42), .A2(n41), .ZN(N350) );
  ND2D1BWP30P140 U37 ( .A1(n85), .A2(i_data_bus[63]), .ZN(n41) );
  IND2D1BWP30P140 U38 ( .A1(n54), .B1(n40), .ZN(n42) );
  INR2D1BWP30P140 U39 ( .A1(i_data_bus[31]), .B1(n53), .ZN(n40) );
  CKND2D4BWP30P140 U40 ( .A1(i_cmd[1]), .A2(n4), .ZN(n32) );
  INVD1BWP30P140 U41 ( .I(n50), .ZN(n51) );
  INVD1BWP30P140 U42 ( .I(n36), .ZN(n49) );
  INVD1BWP30P140 U43 ( .I(n44), .ZN(n4) );
  INVD1BWP30P140 U44 ( .I(rst), .ZN(n3) );
  ND2D1BWP30P140 U45 ( .A1(n3), .A2(i_en), .ZN(n44) );
  NR2OPTPAD1BWP30P140 U46 ( .A1(i_cmd[1]), .A2(i_valid[0]), .ZN(n8) );
  ND2OPTPAD4BWP30P140 U47 ( .A1(n10), .A2(n9), .ZN(n101) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[50]), .ZN(n13) );
  INVD2BWP30P140 U49 ( .I(n35), .ZN(n12) );
  BUFFD2BWP30P140 U50 ( .I(n17), .Z(n47) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[18]), .ZN(n74) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[63]), .ZN(n18) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[31]), .ZN(n39) );
  OAI22OPTPBD2BWP30P140 U54 ( .A1(n2), .A2(n18), .B1(n27), .B2(n39), .ZN(N318)
         );
  INVD1BWP30P140 U55 ( .I(i_data_bus[62]), .ZN(n19) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[30]), .ZN(n87) );
  OAI22OPTPBD2BWP30P140 U57 ( .A1(n2), .A2(n19), .B1(n27), .B2(n87), .ZN(N317)
         );
  INVD1BWP30P140 U58 ( .I(i_data_bus[61]), .ZN(n20) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[29]), .ZN(n84) );
  OAI22OPTPBD2BWP30P140 U60 ( .A1(n2), .A2(n20), .B1(n27), .B2(n84), .ZN(N316)
         );
  INVD1BWP30P140 U61 ( .I(i_data_bus[35]), .ZN(n21) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[3]), .ZN(n59) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[36]), .ZN(n22) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[4]), .ZN(n60) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[37]), .ZN(n23) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[5]), .ZN(n61) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[38]), .ZN(n24) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[6]), .ZN(n62) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[39]), .ZN(n25) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[7]), .ZN(n63) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[49]), .ZN(n26) );
  INVD1BWP30P140 U72 ( .I(i_data_bus[17]), .ZN(n73) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[51]), .ZN(n28) );
  INVD1BWP30P140 U74 ( .I(i_data_bus[19]), .ZN(n30) );
  IND2D4BWP30P140 U75 ( .A1(i_valid[1]), .B1(i_cmd[0]), .ZN(n29) );
  INVD2BWP30P140 U76 ( .I(i_cmd[1]), .ZN(n50) );
  ND2OPTPAD4BWP30P140 U77 ( .A1(n29), .A2(n50), .ZN(n54) );
  OAI21OPTREPBD2BWP30P140 U78 ( .A1(i_cmd[0]), .A2(i_valid[0]), .B(n4), .ZN(
        n53) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[32]), .ZN(n38) );
  CKBD1BWP30P140 U80 ( .I(n35), .Z(n36) );
  CKBD1BWP30P140 U81 ( .I(i_cmd[0]), .Z(n43) );
  ND3D1BWP30P140 U82 ( .A1(n49), .A2(n45), .A3(i_data_bus[0]), .ZN(n37) );
  OAI21D2BWP30P140 U83 ( .A1(n2), .A2(n38), .B(n37), .ZN(N287) );
  INVD1BWP30P140 U84 ( .I(i_valid[1]), .ZN(n46) );
  INVD1BWP30P140 U85 ( .I(n85), .ZN(n52) );
  OAI21D1BWP30P140 U86 ( .A1(n36), .A2(n51), .B(n52), .ZN(N354) );
  INVD1BWP30P140 U87 ( .I(i_data_bus[0]), .ZN(n56) );
  NR2OPTPAD4BWP30P140 U88 ( .A1(n54), .A2(n53), .ZN(n55) );
  MOAI22D1BWP30P140 U89 ( .A1(n56), .A2(n86), .B1(i_data_bus[32]), .B2(n85), 
        .ZN(N319) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[1]), .ZN(n57) );
  MOAI22D1BWP30P140 U91 ( .A1(n57), .A2(n86), .B1(i_data_bus[33]), .B2(n85), 
        .ZN(N320) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[2]), .ZN(n58) );
  MOAI22D1BWP30P140 U93 ( .A1(n58), .A2(n86), .B1(i_data_bus[34]), .B2(n85), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U94 ( .A1(n59), .A2(n86), .B1(i_data_bus[35]), .B2(n85), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U95 ( .A1(n60), .A2(n86), .B1(i_data_bus[36]), .B2(n85), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U96 ( .A1(n61), .A2(n86), .B1(i_data_bus[37]), .B2(n85), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U97 ( .A1(n62), .A2(n86), .B1(i_data_bus[38]), .B2(n85), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U98 ( .A1(n63), .A2(n86), .B1(i_data_bus[39]), .B2(n85), 
        .ZN(N326) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[8]), .ZN(n64) );
  MOAI22D1BWP30P140 U100 ( .A1(n64), .A2(n86), .B1(i_data_bus[40]), .B2(n85), 
        .ZN(N327) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[9]), .ZN(n65) );
  MOAI22D1BWP30P140 U102 ( .A1(n65), .A2(n86), .B1(i_data_bus[41]), .B2(n85), 
        .ZN(N328) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[10]), .ZN(n66) );
  MOAI22D1BWP30P140 U104 ( .A1(n66), .A2(n86), .B1(i_data_bus[42]), .B2(n85), 
        .ZN(N329) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[11]), .ZN(n67) );
  MOAI22D1BWP30P140 U106 ( .A1(n67), .A2(n86), .B1(i_data_bus[43]), .B2(n85), 
        .ZN(N330) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[12]), .ZN(n68) );
  MOAI22D1BWP30P140 U108 ( .A1(n68), .A2(n86), .B1(i_data_bus[44]), .B2(n85), 
        .ZN(N331) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[13]), .ZN(n69) );
  MOAI22D1BWP30P140 U110 ( .A1(n69), .A2(n86), .B1(i_data_bus[45]), .B2(n85), 
        .ZN(N332) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[14]), .ZN(n70) );
  MOAI22D1BWP30P140 U112 ( .A1(n70), .A2(n86), .B1(i_data_bus[46]), .B2(n85), 
        .ZN(N333) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[15]), .ZN(n71) );
  MOAI22D1BWP30P140 U114 ( .A1(n71), .A2(n86), .B1(i_data_bus[47]), .B2(n85), 
        .ZN(N334) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[16]), .ZN(n72) );
  MOAI22D1BWP30P140 U116 ( .A1(n72), .A2(n86), .B1(i_data_bus[48]), .B2(n85), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U117 ( .A1(n73), .A2(n86), .B1(i_data_bus[49]), .B2(n85), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U118 ( .A1(n74), .A2(n86), .B1(i_data_bus[50]), .B2(n85), 
        .ZN(N337) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[20]), .ZN(n75) );
  MOAI22D1BWP30P140 U120 ( .A1(n75), .A2(n86), .B1(i_data_bus[52]), .B2(n85), 
        .ZN(N339) );
  INVD1BWP30P140 U121 ( .I(i_data_bus[21]), .ZN(n76) );
  MOAI22D1BWP30P140 U122 ( .A1(n76), .A2(n86), .B1(i_data_bus[53]), .B2(n85), 
        .ZN(N340) );
  INVD1BWP30P140 U123 ( .I(i_data_bus[22]), .ZN(n77) );
  MOAI22D1BWP30P140 U124 ( .A1(n77), .A2(n86), .B1(i_data_bus[54]), .B2(n85), 
        .ZN(N341) );
  INVD1BWP30P140 U125 ( .I(i_data_bus[23]), .ZN(n78) );
  MOAI22D1BWP30P140 U126 ( .A1(n78), .A2(n86), .B1(i_data_bus[55]), .B2(n85), 
        .ZN(N342) );
  INVD1BWP30P140 U127 ( .I(i_data_bus[24]), .ZN(n79) );
  MOAI22D1BWP30P140 U128 ( .A1(n79), .A2(n86), .B1(i_data_bus[56]), .B2(n85), 
        .ZN(N343) );
  INVD1BWP30P140 U129 ( .I(i_data_bus[25]), .ZN(n80) );
  MOAI22D1BWP30P140 U130 ( .A1(n80), .A2(n86), .B1(i_data_bus[57]), .B2(n85), 
        .ZN(N344) );
  INVD1BWP30P140 U131 ( .I(i_data_bus[26]), .ZN(n81) );
  MOAI22D1BWP30P140 U132 ( .A1(n81), .A2(n86), .B1(i_data_bus[58]), .B2(n85), 
        .ZN(N345) );
  INVD1BWP30P140 U133 ( .I(i_data_bus[27]), .ZN(n82) );
  MOAI22D1BWP30P140 U134 ( .A1(n82), .A2(n86), .B1(i_data_bus[59]), .B2(n85), 
        .ZN(N346) );
  INVD1BWP30P140 U135 ( .I(i_data_bus[28]), .ZN(n83) );
  MOAI22D1BWP30P140 U136 ( .A1(n83), .A2(n86), .B1(i_data_bus[60]), .B2(n85), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U137 ( .A1(n84), .A2(n86), .B1(i_data_bus[61]), .B2(n85), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U138 ( .A1(n87), .A2(n86), .B1(i_data_bus[62]), .B2(n85), 
        .ZN(N349) );
  INVD1BWP30P140 U139 ( .I(i_data_bus[60]), .ZN(n88) );
  MOAI22D1BWP30P140 U140 ( .A1(n2), .A2(n88), .B1(n107), .B2(i_data_bus[28]), 
        .ZN(N315) );
  INVD1BWP30P140 U141 ( .I(i_data_bus[48]), .ZN(n89) );
  MOAI22D1BWP30P140 U142 ( .A1(n2), .A2(n89), .B1(n107), .B2(i_data_bus[16]), 
        .ZN(N303) );
  INVD1BWP30P140 U143 ( .I(i_data_bus[34]), .ZN(n90) );
  MOAI22D1BWP30P140 U144 ( .A1(n2), .A2(n90), .B1(n107), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140 U145 ( .I(i_data_bus[59]), .ZN(n91) );
  MOAI22D1BWP30P140 U146 ( .A1(n2), .A2(n91), .B1(n107), .B2(i_data_bus[27]), 
        .ZN(N314) );
  INVD1BWP30P140 U147 ( .I(i_data_bus[47]), .ZN(n92) );
  MOAI22D1BWP30P140 U148 ( .A1(n2), .A2(n92), .B1(n107), .B2(i_data_bus[15]), 
        .ZN(N302) );
  INVD1BWP30P140 U149 ( .I(i_data_bus[33]), .ZN(n93) );
  MOAI22D1BWP30P140 U150 ( .A1(n2), .A2(n93), .B1(n107), .B2(i_data_bus[1]), 
        .ZN(N288) );
  INVD1BWP30P140 U151 ( .I(i_data_bus[58]), .ZN(n94) );
  MOAI22D1BWP30P140 U152 ( .A1(n2), .A2(n94), .B1(n107), .B2(i_data_bus[26]), 
        .ZN(N313) );
  INVD1BWP30P140 U153 ( .I(i_data_bus[46]), .ZN(n95) );
  MOAI22D1BWP30P140 U154 ( .A1(n2), .A2(n95), .B1(n107), .B2(i_data_bus[14]), 
        .ZN(N301) );
  INVD1BWP30P140 U155 ( .I(i_data_bus[57]), .ZN(n96) );
  MOAI22D1BWP30P140 U156 ( .A1(n2), .A2(n96), .B1(n107), .B2(i_data_bus[25]), 
        .ZN(N312) );
  INVD1BWP30P140 U157 ( .I(i_data_bus[45]), .ZN(n97) );
  MOAI22D1BWP30P140 U158 ( .A1(n2), .A2(n97), .B1(n107), .B2(i_data_bus[13]), 
        .ZN(N300) );
  INVD1BWP30P140 U159 ( .I(i_data_bus[56]), .ZN(n98) );
  MOAI22D1BWP30P140 U160 ( .A1(n2), .A2(n98), .B1(n107), .B2(i_data_bus[24]), 
        .ZN(N311) );
  INVD1BWP30P140 U161 ( .I(i_data_bus[44]), .ZN(n99) );
  MOAI22D1BWP30P140 U162 ( .A1(n2), .A2(n99), .B1(n107), .B2(i_data_bus[12]), 
        .ZN(N299) );
  INVD1BWP30P140 U163 ( .I(i_data_bus[55]), .ZN(n100) );
  MOAI22D1BWP30P140 U164 ( .A1(n101), .A2(n100), .B1(n107), .B2(i_data_bus[23]), .ZN(N310) );
  INVD1BWP30P140 U165 ( .I(i_data_bus[43]), .ZN(n102) );
  MOAI22D1BWP30P140 U166 ( .A1(n2), .A2(n102), .B1(n107), .B2(i_data_bus[11]), 
        .ZN(N298) );
  INVD1BWP30P140 U167 ( .I(i_data_bus[54]), .ZN(n103) );
  MOAI22D1BWP30P140 U168 ( .A1(n2), .A2(n103), .B1(n107), .B2(i_data_bus[22]), 
        .ZN(N309) );
  INVD1BWP30P140 U169 ( .I(i_data_bus[42]), .ZN(n104) );
  MOAI22D1BWP30P140 U170 ( .A1(n2), .A2(n104), .B1(n107), .B2(i_data_bus[10]), 
        .ZN(N297) );
  INVD1BWP30P140 U171 ( .I(i_data_bus[53]), .ZN(n105) );
  MOAI22D1BWP30P140 U172 ( .A1(n2), .A2(n105), .B1(n107), .B2(i_data_bus[21]), 
        .ZN(N308) );
  INVD1BWP30P140 U173 ( .I(i_data_bus[41]), .ZN(n106) );
  MOAI22D1BWP30P140 U174 ( .A1(n2), .A2(n106), .B1(n107), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140 U175 ( .I(i_data_bus[52]), .ZN(n108) );
  MOAI22D1BWP30P140 U176 ( .A1(n2), .A2(n108), .B1(n107), .B2(i_data_bus[20]), 
        .ZN(N307) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_141 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  ND2OPTPAD6BWP30P140 U3 ( .A1(n24), .A2(n15), .ZN(n73) );
  CKND2D3BWP30P140 U4 ( .A1(i_cmd[1]), .A2(n6), .ZN(n21) );
  INVD1BWP30P140 U5 ( .I(i_cmd[1]), .ZN(n25) );
  INVD6BWP30P140 U6 ( .I(n44), .ZN(n1) );
  ND2D1BWP30P140 U7 ( .A1(n11), .A2(n10), .ZN(n2) );
  CKND2D4BWP30P140 U8 ( .A1(n11), .A2(n10), .ZN(n3) );
  IND2D1BWP30P140 U9 ( .A1(n17), .B1(n73), .ZN(N353) );
  NR3D0BWP30P140 U10 ( .A1(n16), .A2(n15), .A3(n18), .ZN(n17) );
  INVD1BWP30P140 U11 ( .I(n71), .ZN(n26) );
  IND2D1BWP30P140 U12 ( .A1(n14), .B1(n13), .ZN(N295) );
  NR2D1BWP30P140 U13 ( .A1(n73), .A2(n49), .ZN(n14) );
  OR2D1BWP30P140 U14 ( .A1(n12), .A2(n2), .Z(n13) );
  ND2D1BWP30P140 U15 ( .A1(n23), .A2(n22), .ZN(N350) );
  ND2D1BWP30P140 U16 ( .A1(n44), .A2(i_data_bus[31]), .ZN(n23) );
  ND2D1BWP30P140 U17 ( .A1(n71), .A2(i_data_bus[63]), .ZN(n22) );
  ND2OPTIBD4BWP30P140 U18 ( .A1(n11), .A2(n10), .ZN(n95) );
  INVD1BWP30P140 U19 ( .I(n18), .ZN(n6) );
  INVD1BWP30P140 U20 ( .I(rst), .ZN(n4) );
  ND2D1BWP30P140 U21 ( .A1(n4), .A2(i_en), .ZN(n18) );
  CKND2D2BWP30P140 U22 ( .A1(i_valid[0]), .A2(n6), .ZN(n5) );
  INVD3BWP30P140 U23 ( .I(n5), .ZN(n24) );
  INVD2BWP30P140 U24 ( .I(i_cmd[0]), .ZN(n15) );
  INVD1BWP30P140 U25 ( .I(i_data_bus[40]), .ZN(n12) );
  NR2D1BWP30P140 U26 ( .A1(i_cmd[1]), .A2(i_valid[0]), .ZN(n8) );
  ND2OPTIBD4BWP30P140 U27 ( .A1(i_cmd[0]), .A2(n6), .ZN(n7) );
  NR2OPTPAD4BWP30P140 U28 ( .A1(n8), .A2(n7), .ZN(n11) );
  INVD1BWP30P140 U29 ( .I(i_valid[1]), .ZN(n9) );
  ND2OPTIBD2BWP30P140 U30 ( .A1(n9), .A2(i_cmd[1]), .ZN(n10) );
  INVD1BWP30P140 U31 ( .I(i_valid[1]), .ZN(n16) );
  CKND2D3BWP30P140 U32 ( .A1(n25), .A2(n6), .ZN(n20) );
  MUX2NOPTD2BWP30P140 U33 ( .I0(i_valid[0]), .I1(i_valid[1]), .S(i_cmd[0]), 
        .ZN(n19) );
  NR2OPTPAD4BWP30P140 U34 ( .A1(n19), .A2(n20), .ZN(n44) );
  INVD1BWP30P140 U35 ( .I(i_data_bus[31]), .ZN(n34) );
  INR2D8BWP30P140 U36 ( .A1(i_valid[1]), .B1(n21), .ZN(n71) );
  INVD1BWP30P140 U37 ( .I(n24), .ZN(n27) );
  OAI21D1BWP30P140 U38 ( .A1(n27), .A2(i_cmd[1]), .B(n26), .ZN(N354) );
  INVD1BWP30P140 U39 ( .I(i_data_bus[17]), .ZN(n58) );
  INVD1BWP30P140 U40 ( .I(i_data_bus[49]), .ZN(n28) );
  OAI22D1BWP30P140 U41 ( .A1(n73), .A2(n58), .B1(n3), .B2(n28), .ZN(N304) );
  INVD1BWP30P140 U42 ( .I(i_data_bus[18]), .ZN(n59) );
  INVD1BWP30P140 U43 ( .I(i_data_bus[50]), .ZN(n29) );
  OAI22D1BWP30P140 U44 ( .A1(n73), .A2(n59), .B1(n95), .B2(n29), .ZN(N305) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[19]), .ZN(n60) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[51]), .ZN(n30) );
  OAI22D1BWP30P140 U47 ( .A1(n73), .A2(n60), .B1(n3), .B2(n30), .ZN(N306) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[29]), .ZN(n70) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[61]), .ZN(n31) );
  OAI22D1BWP30P140 U50 ( .A1(n73), .A2(n70), .B1(n95), .B2(n31), .ZN(N316) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[30]), .ZN(n72) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[62]), .ZN(n32) );
  OAI22D1BWP30P140 U53 ( .A1(n73), .A2(n72), .B1(n3), .B2(n32), .ZN(N317) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[63]), .ZN(n33) );
  OAI22D1BWP30P140 U55 ( .A1(n73), .A2(n34), .B1(n95), .B2(n33), .ZN(N318) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[3]), .ZN(n43) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[35]), .ZN(n35) );
  OAI22D1BWP30P140 U58 ( .A1(n73), .A2(n43), .B1(n3), .B2(n35), .ZN(N290) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[7]), .ZN(n48) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[39]), .ZN(n36) );
  OAI22D1BWP30P140 U61 ( .A1(n73), .A2(n48), .B1(n95), .B2(n36), .ZN(N294) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[6]), .ZN(n47) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[38]), .ZN(n37) );
  OAI22D1BWP30P140 U64 ( .A1(n73), .A2(n47), .B1(n3), .B2(n37), .ZN(N293) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[5]), .ZN(n46) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[37]), .ZN(n38) );
  OAI22D1BWP30P140 U67 ( .A1(n73), .A2(n46), .B1(n95), .B2(n38), .ZN(N292) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[4]), .ZN(n45) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[36]), .ZN(n39) );
  OAI22D1BWP30P140 U70 ( .A1(n73), .A2(n45), .B1(n95), .B2(n39), .ZN(N291) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[0]), .ZN(n40) );
  MOAI22D1BWP30P140 U72 ( .A1(n40), .A2(n1), .B1(i_data_bus[32]), .B2(n71), 
        .ZN(N319) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[1]), .ZN(n41) );
  MOAI22D1BWP30P140 U74 ( .A1(n41), .A2(n1), .B1(i_data_bus[33]), .B2(n71), 
        .ZN(N320) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[2]), .ZN(n42) );
  MOAI22D1BWP30P140 U76 ( .A1(n42), .A2(n1), .B1(i_data_bus[34]), .B2(n71), 
        .ZN(N321) );
  MOAI22D1BWP30P140 U77 ( .A1(n43), .A2(n1), .B1(i_data_bus[35]), .B2(n71), 
        .ZN(N322) );
  MOAI22D1BWP30P140 U78 ( .A1(n45), .A2(n1), .B1(i_data_bus[36]), .B2(n71), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U79 ( .A1(n46), .A2(n1), .B1(i_data_bus[37]), .B2(n71), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U80 ( .A1(n47), .A2(n1), .B1(i_data_bus[38]), .B2(n71), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U81 ( .A1(n48), .A2(n1), .B1(i_data_bus[39]), .B2(n71), 
        .ZN(N326) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[8]), .ZN(n49) );
  MOAI22D1BWP30P140 U83 ( .A1(n49), .A2(n1), .B1(i_data_bus[40]), .B2(n71), 
        .ZN(N327) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[9]), .ZN(n50) );
  MOAI22D1BWP30P140 U85 ( .A1(n50), .A2(n1), .B1(i_data_bus[41]), .B2(n71), 
        .ZN(N328) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[10]), .ZN(n51) );
  MOAI22D1BWP30P140 U87 ( .A1(n51), .A2(n1), .B1(i_data_bus[42]), .B2(n71), 
        .ZN(N329) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[11]), .ZN(n52) );
  MOAI22D1BWP30P140 U89 ( .A1(n52), .A2(n1), .B1(i_data_bus[43]), .B2(n71), 
        .ZN(N330) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[12]), .ZN(n53) );
  MOAI22D1BWP30P140 U91 ( .A1(n53), .A2(n1), .B1(i_data_bus[44]), .B2(n71), 
        .ZN(N331) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[13]), .ZN(n54) );
  MOAI22D1BWP30P140 U93 ( .A1(n54), .A2(n1), .B1(i_data_bus[45]), .B2(n71), 
        .ZN(N332) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[14]), .ZN(n55) );
  MOAI22D1BWP30P140 U95 ( .A1(n55), .A2(n1), .B1(i_data_bus[46]), .B2(n71), 
        .ZN(N333) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[15]), .ZN(n56) );
  MOAI22D1BWP30P140 U97 ( .A1(n56), .A2(n1), .B1(i_data_bus[47]), .B2(n71), 
        .ZN(N334) );
  INVD1BWP30P140 U98 ( .I(i_data_bus[16]), .ZN(n57) );
  MOAI22D1BWP30P140 U99 ( .A1(n57), .A2(n1), .B1(i_data_bus[48]), .B2(n71), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U100 ( .A1(n58), .A2(n1), .B1(i_data_bus[49]), .B2(n71), 
        .ZN(N336) );
  MOAI22D1BWP30P140 U101 ( .A1(n59), .A2(n1), .B1(i_data_bus[50]), .B2(n71), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U102 ( .A1(n60), .A2(n1), .B1(i_data_bus[51]), .B2(n71), 
        .ZN(N338) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[20]), .ZN(n61) );
  MOAI22D1BWP30P140 U104 ( .A1(n61), .A2(n1), .B1(i_data_bus[52]), .B2(n71), 
        .ZN(N339) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[21]), .ZN(n62) );
  MOAI22D1BWP30P140 U106 ( .A1(n62), .A2(n1), .B1(i_data_bus[53]), .B2(n71), 
        .ZN(N340) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[22]), .ZN(n63) );
  MOAI22D1BWP30P140 U108 ( .A1(n63), .A2(n1), .B1(i_data_bus[54]), .B2(n71), 
        .ZN(N341) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[23]), .ZN(n64) );
  MOAI22D1BWP30P140 U110 ( .A1(n64), .A2(n1), .B1(i_data_bus[55]), .B2(n71), 
        .ZN(N342) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[24]), .ZN(n65) );
  MOAI22D1BWP30P140 U112 ( .A1(n65), .A2(n1), .B1(i_data_bus[56]), .B2(n71), 
        .ZN(N343) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[25]), .ZN(n66) );
  MOAI22D1BWP30P140 U114 ( .A1(n66), .A2(n1), .B1(i_data_bus[57]), .B2(n71), 
        .ZN(N344) );
  INVD1BWP30P140 U115 ( .I(i_data_bus[26]), .ZN(n67) );
  MOAI22D1BWP30P140 U116 ( .A1(n67), .A2(n1), .B1(i_data_bus[58]), .B2(n71), 
        .ZN(N345) );
  INVD1BWP30P140 U117 ( .I(i_data_bus[27]), .ZN(n68) );
  MOAI22D1BWP30P140 U118 ( .A1(n68), .A2(n1), .B1(i_data_bus[59]), .B2(n71), 
        .ZN(N346) );
  INVD1BWP30P140 U119 ( .I(i_data_bus[28]), .ZN(n69) );
  MOAI22D1BWP30P140 U120 ( .A1(n69), .A2(n1), .B1(i_data_bus[60]), .B2(n71), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U121 ( .A1(n70), .A2(n1), .B1(i_data_bus[61]), .B2(n71), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U122 ( .A1(n72), .A2(n1), .B1(i_data_bus[62]), .B2(n71), 
        .ZN(N349) );
  INVD1BWP30P140 U123 ( .I(i_data_bus[60]), .ZN(n74) );
  INVD8BWP30P140 U124 ( .I(n73), .ZN(n93) );
  MOAI22D1BWP30P140 U125 ( .A1(n3), .A2(n74), .B1(n93), .B2(i_data_bus[28]), 
        .ZN(N315) );
  INVD1BWP30P140 U126 ( .I(i_data_bus[48]), .ZN(n75) );
  MOAI22D1BWP30P140 U127 ( .A1(n3), .A2(n75), .B1(n93), .B2(i_data_bus[16]), 
        .ZN(N303) );
  INVD1BWP30P140 U128 ( .I(i_data_bus[34]), .ZN(n76) );
  MOAI22D1BWP30P140 U129 ( .A1(n95), .A2(n76), .B1(n93), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140 U130 ( .I(i_data_bus[59]), .ZN(n77) );
  MOAI22D1BWP30P140 U131 ( .A1(n3), .A2(n77), .B1(n93), .B2(i_data_bus[27]), 
        .ZN(N314) );
  INVD1BWP30P140 U132 ( .I(i_data_bus[47]), .ZN(n78) );
  MOAI22D1BWP30P140 U133 ( .A1(n95), .A2(n78), .B1(n93), .B2(i_data_bus[15]), 
        .ZN(N302) );
  INVD1BWP30P140 U134 ( .I(i_data_bus[33]), .ZN(n79) );
  MOAI22D1BWP30P140 U135 ( .A1(n3), .A2(n79), .B1(n93), .B2(i_data_bus[1]), 
        .ZN(N288) );
  INVD1BWP30P140 U136 ( .I(i_data_bus[58]), .ZN(n80) );
  MOAI22D1BWP30P140 U137 ( .A1(n95), .A2(n80), .B1(n93), .B2(i_data_bus[26]), 
        .ZN(N313) );
  INVD1BWP30P140 U138 ( .I(i_data_bus[46]), .ZN(n81) );
  MOAI22D1BWP30P140 U139 ( .A1(n3), .A2(n81), .B1(n93), .B2(i_data_bus[14]), 
        .ZN(N301) );
  INVD1BWP30P140 U140 ( .I(i_data_bus[32]), .ZN(n82) );
  MOAI22D1BWP30P140 U141 ( .A1(n95), .A2(n82), .B1(n93), .B2(i_data_bus[0]), 
        .ZN(N287) );
  INVD1BWP30P140 U142 ( .I(i_data_bus[57]), .ZN(n83) );
  MOAI22D1BWP30P140 U143 ( .A1(n3), .A2(n83), .B1(n93), .B2(i_data_bus[25]), 
        .ZN(N312) );
  INVD1BWP30P140 U144 ( .I(i_data_bus[45]), .ZN(n84) );
  MOAI22D1BWP30P140 U145 ( .A1(n95), .A2(n84), .B1(n93), .B2(i_data_bus[13]), 
        .ZN(N300) );
  INVD1BWP30P140 U146 ( .I(i_data_bus[56]), .ZN(n85) );
  MOAI22D1BWP30P140 U147 ( .A1(n3), .A2(n85), .B1(n93), .B2(i_data_bus[24]), 
        .ZN(N311) );
  INVD1BWP30P140 U148 ( .I(i_data_bus[44]), .ZN(n86) );
  MOAI22D1BWP30P140 U149 ( .A1(n95), .A2(n86), .B1(n93), .B2(i_data_bus[12]), 
        .ZN(N299) );
  INVD1BWP30P140 U150 ( .I(i_data_bus[55]), .ZN(n87) );
  MOAI22D1BWP30P140 U151 ( .A1(n3), .A2(n87), .B1(n93), .B2(i_data_bus[23]), 
        .ZN(N310) );
  INVD1BWP30P140 U152 ( .I(i_data_bus[43]), .ZN(n88) );
  MOAI22D1BWP30P140 U153 ( .A1(n95), .A2(n88), .B1(n93), .B2(i_data_bus[11]), 
        .ZN(N298) );
  INVD1BWP30P140 U154 ( .I(i_data_bus[54]), .ZN(n89) );
  MOAI22D1BWP30P140 U155 ( .A1(n3), .A2(n89), .B1(n93), .B2(i_data_bus[22]), 
        .ZN(N309) );
  INVD1BWP30P140 U156 ( .I(i_data_bus[42]), .ZN(n90) );
  MOAI22D1BWP30P140 U157 ( .A1(n95), .A2(n90), .B1(n93), .B2(i_data_bus[10]), 
        .ZN(N297) );
  INVD1BWP30P140 U158 ( .I(i_data_bus[53]), .ZN(n91) );
  MOAI22D1BWP30P140 U159 ( .A1(n3), .A2(n91), .B1(n93), .B2(i_data_bus[21]), 
        .ZN(N308) );
  INVD1BWP30P140 U160 ( .I(i_data_bus[41]), .ZN(n92) );
  MOAI22D1BWP30P140 U161 ( .A1(n95), .A2(n92), .B1(n93), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140 U162 ( .I(i_data_bus[52]), .ZN(n94) );
  MOAI22D1BWP30P140 U163 ( .A1(n3), .A2(n94), .B1(n93), .B2(i_data_bus[20]), 
        .ZN(N307) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_142 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  CKND2D3BWP30P140 U3 ( .A1(n11), .A2(n10), .ZN(n3) );
  NR2OPTPAD2BWP30P140 U4 ( .A1(n19), .A2(n20), .ZN(n44) );
  INVD1P5BWP30P140 U5 ( .I(i_cmd[0]), .ZN(n15) );
  ND2OPTIBD2BWP30P140 U6 ( .A1(n9), .A2(i_cmd[1]), .ZN(n10) );
  CKND2D2BWP30P140 U7 ( .A1(n25), .A2(n6), .ZN(n20) );
  ND2OPTPAD6BWP30P140 U8 ( .A1(n24), .A2(n15), .ZN(n73) );
  INVD6BWP30P140 U9 ( .I(n44), .ZN(n1) );
  INVD3BWP30P140 U10 ( .I(n5), .ZN(n24) );
  INVD8BWP30P140 U11 ( .I(n73), .ZN(n93) );
  OAI22D1BWP30P140 U12 ( .A1(n3), .A2(n29), .B1(n73), .B2(n45), .ZN(N318) );
  OAI22D1BWP30P140 U13 ( .A1(n3), .A2(n31), .B1(n73), .B2(n42), .ZN(N316) );
  OAI22D1BWP30P140 U14 ( .A1(n3), .A2(n33), .B1(n73), .B2(n53), .ZN(N305) );
  OAI22D1BWP30P140 U15 ( .A1(n3), .A2(n35), .B1(n73), .B2(n69), .ZN(N290) );
  OAI22D1BWP30P140 U16 ( .A1(n3), .A2(n37), .B1(n73), .B2(n67), .ZN(N292) );
  NR2D1BWP30P140 U17 ( .A1(i_cmd[1]), .A2(i_valid[0]), .ZN(n8) );
  MUX2NOPTD2BWP30P140 U18 ( .I0(i_valid[0]), .I1(i_valid[1]), .S(i_cmd[0]), 
        .ZN(n19) );
  CKND2D4BWP30P140 U19 ( .A1(n11), .A2(n10), .ZN(n95) );
  INVD1BWP30P140 U20 ( .I(i_valid[1]), .ZN(n9) );
  ND2OPTIBD1BWP30P140 U21 ( .A1(n11), .A2(n10), .ZN(n2) );
  IND2D1BWP30P140 U22 ( .A1(n17), .B1(n73), .ZN(N353) );
  NR3D0BWP30P140 U23 ( .A1(n16), .A2(n15), .A3(n18), .ZN(n17) );
  INVD1BWP30P140 U24 ( .I(n71), .ZN(n27) );
  IND2D1BWP30P140 U25 ( .A1(n14), .B1(n13), .ZN(N307) );
  NR2D1BWP30P140 U26 ( .A1(n73), .A2(n51), .ZN(n14) );
  OR2D1BWP30P140 U27 ( .A1(n12), .A2(n2), .Z(n13) );
  ND2D1BWP30P140 U28 ( .A1(n23), .A2(n22), .ZN(N319) );
  ND2D1BWP30P140 U29 ( .A1(n44), .A2(i_data_bus[0]), .ZN(n23) );
  ND2D1BWP30P140 U30 ( .A1(n71), .A2(i_data_bus[32]), .ZN(n22) );
  INVD1BWP30P140 U31 ( .I(n18), .ZN(n6) );
  INVD1BWP30P140 U32 ( .I(n25), .ZN(n26) );
  INVD1BWP30P140 U33 ( .I(rst), .ZN(n4) );
  ND2D1BWP30P140 U34 ( .A1(n4), .A2(i_en), .ZN(n18) );
  CKND2D2BWP30P140 U35 ( .A1(i_valid[0]), .A2(n6), .ZN(n5) );
  INVD1BWP30P140 U36 ( .I(i_data_bus[52]), .ZN(n12) );
  ND2OPTPAD2BWP30P140 U37 ( .A1(i_cmd[0]), .A2(n6), .ZN(n7) );
  NR2OPTPAD2BWP30P140 U38 ( .A1(n8), .A2(n7), .ZN(n11) );
  INVD1BWP30P140 U39 ( .I(i_valid[1]), .ZN(n16) );
  INVD2BWP30P140 U40 ( .I(i_cmd[1]), .ZN(n25) );
  ND2OPTPAD2BWP30P140 U41 ( .A1(i_cmd[1]), .A2(n6), .ZN(n21) );
  INR2D8BWP30P140 U42 ( .A1(i_valid[1]), .B1(n21), .ZN(n71) );
  INVD1BWP30P140 U43 ( .I(n24), .ZN(n28) );
  OAI21D1BWP30P140 U44 ( .A1(n28), .A2(n26), .B(n27), .ZN(N354) );
  INVD1BWP30P140 U45 ( .I(i_data_bus[31]), .ZN(n45) );
  INVD1BWP30P140 U46 ( .I(i_data_bus[63]), .ZN(n29) );
  INVD1BWP30P140 U47 ( .I(i_data_bus[30]), .ZN(n43) );
  INVD1BWP30P140 U48 ( .I(i_data_bus[62]), .ZN(n30) );
  OAI22D1BWP30P140 U49 ( .A1(n73), .A2(n43), .B1(n95), .B2(n30), .ZN(N317) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[29]), .ZN(n42) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[61]), .ZN(n31) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[19]), .ZN(n52) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[51]), .ZN(n32) );
  OAI22D1BWP30P140 U54 ( .A1(n73), .A2(n52), .B1(n95), .B2(n32), .ZN(N306) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[18]), .ZN(n53) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[50]), .ZN(n33) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[17]), .ZN(n54) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[49]), .ZN(n34) );
  OAI22D1BWP30P140 U59 ( .A1(n73), .A2(n54), .B1(n95), .B2(n34), .ZN(N304) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[3]), .ZN(n69) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[35]), .ZN(n35) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[4]), .ZN(n68) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[36]), .ZN(n36) );
  OAI22D1BWP30P140 U64 ( .A1(n73), .A2(n68), .B1(n95), .B2(n36), .ZN(N291) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[5]), .ZN(n67) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[37]), .ZN(n37) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[6]), .ZN(n66) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[38]), .ZN(n38) );
  OAI22D1BWP30P140 U69 ( .A1(n73), .A2(n66), .B1(n95), .B2(n38), .ZN(N293) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[7]), .ZN(n65) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[39]), .ZN(n39) );
  OAI22D1BWP30P140 U72 ( .A1(n73), .A2(n65), .B1(n95), .B2(n39), .ZN(N294) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[26]), .ZN(n40) );
  MOAI22D1BWP30P140 U74 ( .A1(n40), .A2(n1), .B1(i_data_bus[58]), .B2(n71), 
        .ZN(N345) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[28]), .ZN(n41) );
  MOAI22D1BWP30P140 U76 ( .A1(n41), .A2(n1), .B1(i_data_bus[60]), .B2(n71), 
        .ZN(N347) );
  MOAI22D1BWP30P140 U77 ( .A1(n42), .A2(n1), .B1(i_data_bus[61]), .B2(n71), 
        .ZN(N348) );
  MOAI22D1BWP30P140 U78 ( .A1(n43), .A2(n1), .B1(i_data_bus[62]), .B2(n71), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U79 ( .A1(n45), .A2(n1), .B1(i_data_bus[63]), .B2(n71), 
        .ZN(N350) );
  INVD1BWP30P140 U80 ( .I(i_data_bus[25]), .ZN(n46) );
  MOAI22D1BWP30P140 U81 ( .A1(n46), .A2(n1), .B1(i_data_bus[57]), .B2(n71), 
        .ZN(N344) );
  INVD1BWP30P140 U82 ( .I(i_data_bus[24]), .ZN(n47) );
  MOAI22D1BWP30P140 U83 ( .A1(n47), .A2(n1), .B1(i_data_bus[56]), .B2(n71), 
        .ZN(N343) );
  INVD1BWP30P140 U84 ( .I(i_data_bus[23]), .ZN(n48) );
  MOAI22D1BWP30P140 U85 ( .A1(n48), .A2(n1), .B1(i_data_bus[55]), .B2(n71), 
        .ZN(N342) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[22]), .ZN(n49) );
  MOAI22D1BWP30P140 U87 ( .A1(n49), .A2(n1), .B1(i_data_bus[54]), .B2(n71), 
        .ZN(N341) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[21]), .ZN(n50) );
  MOAI22D1BWP30P140 U89 ( .A1(n50), .A2(n1), .B1(i_data_bus[53]), .B2(n71), 
        .ZN(N340) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[20]), .ZN(n51) );
  MOAI22D1BWP30P140 U91 ( .A1(n51), .A2(n1), .B1(i_data_bus[52]), .B2(n71), 
        .ZN(N339) );
  MOAI22D1BWP30P140 U92 ( .A1(n52), .A2(n1), .B1(i_data_bus[51]), .B2(n71), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U93 ( .A1(n53), .A2(n1), .B1(i_data_bus[50]), .B2(n71), 
        .ZN(N337) );
  MOAI22D1BWP30P140 U94 ( .A1(n54), .A2(n1), .B1(i_data_bus[49]), .B2(n71), 
        .ZN(N336) );
  INVD1BWP30P140 U95 ( .I(i_data_bus[16]), .ZN(n55) );
  MOAI22D1BWP30P140 U96 ( .A1(n55), .A2(n1), .B1(i_data_bus[48]), .B2(n71), 
        .ZN(N335) );
  INVD1BWP30P140 U97 ( .I(i_data_bus[15]), .ZN(n56) );
  MOAI22D1BWP30P140 U98 ( .A1(n56), .A2(n1), .B1(i_data_bus[47]), .B2(n71), 
        .ZN(N334) );
  INVD1BWP30P140 U99 ( .I(i_data_bus[14]), .ZN(n57) );
  MOAI22D1BWP30P140 U100 ( .A1(n57), .A2(n1), .B1(i_data_bus[46]), .B2(n71), 
        .ZN(N333) );
  INVD1BWP30P140 U101 ( .I(i_data_bus[13]), .ZN(n58) );
  MOAI22D1BWP30P140 U102 ( .A1(n58), .A2(n1), .B1(i_data_bus[45]), .B2(n71), 
        .ZN(N332) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[12]), .ZN(n59) );
  MOAI22D1BWP30P140 U104 ( .A1(n59), .A2(n1), .B1(i_data_bus[44]), .B2(n71), 
        .ZN(N331) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[11]), .ZN(n60) );
  MOAI22D1BWP30P140 U106 ( .A1(n60), .A2(n1), .B1(i_data_bus[43]), .B2(n71), 
        .ZN(N330) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[10]), .ZN(n61) );
  MOAI22D1BWP30P140 U108 ( .A1(n61), .A2(n1), .B1(i_data_bus[42]), .B2(n71), 
        .ZN(N329) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[27]), .ZN(n62) );
  MOAI22D1BWP30P140 U110 ( .A1(n62), .A2(n1), .B1(i_data_bus[59]), .B2(n71), 
        .ZN(N346) );
  INVD1BWP30P140 U111 ( .I(i_data_bus[9]), .ZN(n63) );
  MOAI22D1BWP30P140 U112 ( .A1(n63), .A2(n1), .B1(i_data_bus[41]), .B2(n71), 
        .ZN(N328) );
  INVD1BWP30P140 U113 ( .I(i_data_bus[8]), .ZN(n64) );
  MOAI22D1BWP30P140 U114 ( .A1(n64), .A2(n1), .B1(i_data_bus[40]), .B2(n71), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U115 ( .A1(n65), .A2(n1), .B1(i_data_bus[39]), .B2(n71), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U116 ( .A1(n66), .A2(n1), .B1(i_data_bus[38]), .B2(n71), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U117 ( .A1(n67), .A2(n1), .B1(i_data_bus[37]), .B2(n71), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U118 ( .A1(n68), .A2(n1), .B1(i_data_bus[36]), .B2(n71), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U119 ( .A1(n69), .A2(n1), .B1(i_data_bus[35]), .B2(n71), 
        .ZN(N322) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[2]), .ZN(n70) );
  MOAI22D1BWP30P140 U121 ( .A1(n70), .A2(n1), .B1(i_data_bus[34]), .B2(n71), 
        .ZN(N321) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[1]), .ZN(n72) );
  MOAI22D1BWP30P140 U123 ( .A1(n72), .A2(n1), .B1(i_data_bus[33]), .B2(n71), 
        .ZN(N320) );
  INVD1BWP30P140 U124 ( .I(i_data_bus[60]), .ZN(n74) );
  MOAI22D1BWP30P140 U125 ( .A1(n3), .A2(n74), .B1(n93), .B2(i_data_bus[28]), 
        .ZN(N315) );
  INVD1BWP30P140 U126 ( .I(i_data_bus[48]), .ZN(n75) );
  MOAI22D1BWP30P140 U127 ( .A1(n3), .A2(n75), .B1(n93), .B2(i_data_bus[16]), 
        .ZN(N303) );
  INVD1BWP30P140 U128 ( .I(i_data_bus[34]), .ZN(n76) );
  MOAI22D1BWP30P140 U129 ( .A1(n95), .A2(n76), .B1(n93), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140 U130 ( .I(i_data_bus[59]), .ZN(n77) );
  MOAI22D1BWP30P140 U131 ( .A1(n3), .A2(n77), .B1(n93), .B2(i_data_bus[27]), 
        .ZN(N314) );
  INVD1BWP30P140 U132 ( .I(i_data_bus[47]), .ZN(n78) );
  MOAI22D1BWP30P140 U133 ( .A1(n95), .A2(n78), .B1(n93), .B2(i_data_bus[15]), 
        .ZN(N302) );
  INVD1BWP30P140 U134 ( .I(i_data_bus[33]), .ZN(n79) );
  MOAI22D1BWP30P140 U135 ( .A1(n3), .A2(n79), .B1(n93), .B2(i_data_bus[1]), 
        .ZN(N288) );
  INVD1BWP30P140 U136 ( .I(i_data_bus[58]), .ZN(n80) );
  MOAI22D1BWP30P140 U137 ( .A1(n95), .A2(n80), .B1(n93), .B2(i_data_bus[26]), 
        .ZN(N313) );
  INVD1BWP30P140 U138 ( .I(i_data_bus[46]), .ZN(n81) );
  MOAI22D1BWP30P140 U139 ( .A1(n3), .A2(n81), .B1(n93), .B2(i_data_bus[14]), 
        .ZN(N301) );
  INVD1BWP30P140 U140 ( .I(i_data_bus[32]), .ZN(n82) );
  MOAI22D1BWP30P140 U141 ( .A1(n95), .A2(n82), .B1(n93), .B2(i_data_bus[0]), 
        .ZN(N287) );
  INVD1BWP30P140 U142 ( .I(i_data_bus[57]), .ZN(n83) );
  MOAI22D1BWP30P140 U143 ( .A1(n3), .A2(n83), .B1(n93), .B2(i_data_bus[25]), 
        .ZN(N312) );
  INVD1BWP30P140 U144 ( .I(i_data_bus[45]), .ZN(n84) );
  MOAI22D1BWP30P140 U145 ( .A1(n95), .A2(n84), .B1(n93), .B2(i_data_bus[13]), 
        .ZN(N300) );
  INVD1BWP30P140 U146 ( .I(i_data_bus[56]), .ZN(n85) );
  MOAI22D1BWP30P140 U147 ( .A1(n3), .A2(n85), .B1(n93), .B2(i_data_bus[24]), 
        .ZN(N311) );
  INVD1BWP30P140 U148 ( .I(i_data_bus[44]), .ZN(n86) );
  MOAI22D1BWP30P140 U149 ( .A1(n95), .A2(n86), .B1(n93), .B2(i_data_bus[12]), 
        .ZN(N299) );
  INVD1BWP30P140 U150 ( .I(i_data_bus[55]), .ZN(n87) );
  MOAI22D1BWP30P140 U151 ( .A1(n3), .A2(n87), .B1(n93), .B2(i_data_bus[23]), 
        .ZN(N310) );
  INVD1BWP30P140 U152 ( .I(i_data_bus[43]), .ZN(n88) );
  MOAI22D1BWP30P140 U153 ( .A1(n95), .A2(n88), .B1(n93), .B2(i_data_bus[11]), 
        .ZN(N298) );
  INVD1BWP30P140 U154 ( .I(i_data_bus[54]), .ZN(n89) );
  MOAI22D1BWP30P140 U155 ( .A1(n3), .A2(n89), .B1(n93), .B2(i_data_bus[22]), 
        .ZN(N309) );
  INVD1BWP30P140 U156 ( .I(i_data_bus[42]), .ZN(n90) );
  MOAI22D1BWP30P140 U157 ( .A1(n95), .A2(n90), .B1(n93), .B2(i_data_bus[10]), 
        .ZN(N297) );
  INVD1BWP30P140 U158 ( .I(i_data_bus[53]), .ZN(n91) );
  MOAI22D1BWP30P140 U159 ( .A1(n3), .A2(n91), .B1(n93), .B2(i_data_bus[21]), 
        .ZN(N308) );
  INVD1BWP30P140 U160 ( .I(i_data_bus[41]), .ZN(n92) );
  MOAI22D1BWP30P140 U161 ( .A1(n95), .A2(n92), .B1(n93), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140 U162 ( .I(i_data_bus[40]), .ZN(n94) );
  MOAI22D1BWP30P140 U163 ( .A1(n3), .A2(n94), .B1(n93), .B2(i_data_bus[8]), 
        .ZN(N295) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_143 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  DFQD1BWP30P140 o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140 o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140 o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140 o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0]) );
  OAI22D1BWP30P140 U3 ( .A1(n93), .A2(n28), .B1(n2), .B2(n45), .ZN(N305) );
  OAI22D1BWP30P140 U4 ( .A1(n93), .A2(n32), .B1(n2), .B2(n63), .ZN(N318) );
  OAI22D1BWP30P140 U5 ( .A1(n93), .A2(n34), .B1(n2), .B2(n57), .ZN(N291) );
  OAI22D1BWP30P140 U6 ( .A1(n93), .A2(n36), .B1(n2), .B2(n55), .ZN(N293) );
  OAI22D1BWP30P140 U7 ( .A1(n93), .A2(n37), .B1(n2), .B2(n54), .ZN(N294) );
  ND2OPTIBD6BWP30P140 U8 ( .A1(n11), .A2(n10), .ZN(n6) );
  ND2D2BWP30P140 U9 ( .A1(n3), .A2(i_cmd[1]), .ZN(n10) );
  CKND2D4BWP30P140 U10 ( .A1(n22), .A2(n14), .ZN(n71) );
  INVD1BWP30P140 U11 ( .I(i_cmd[0]), .ZN(n14) );
  CKND2D3BWP30P140 U12 ( .A1(n23), .A2(n9), .ZN(n18) );
  CKND2D3BWP30P140 U13 ( .A1(i_cmd[0]), .A2(n9), .ZN(n4) );
  NR2D1P5BWP30P140 U14 ( .A1(i_cmd[1]), .A2(i_valid[0]), .ZN(n5) );
  INVD6BWP30P140 U15 ( .I(n71), .ZN(n91) );
  OAI22D1BWP30P140 U16 ( .A1(n6), .A2(n27), .B1(n2), .B2(n47), .ZN(N304) );
  OAI22D1BWP30P140 U17 ( .A1(n93), .A2(n30), .B1(n2), .B2(n65), .ZN(N316) );
  BUFFD12BWP30P140 U18 ( .I(n71), .Z(n2) );
  INVD2BWP30P140 U19 ( .I(n8), .ZN(n22) );
  INVD6BWP30P140 U20 ( .I(n41), .ZN(n1) );
  OAI22OPTPBD1BWP30P140 U21 ( .A1(n6), .A2(n29), .B1(n2), .B2(n44), .ZN(N306)
         );
  OAI22OPTPBD1BWP30P140 U22 ( .A1(n6), .A2(n31), .B1(n2), .B2(n64), .ZN(N317)
         );
  OAI22OPTPBD1BWP30P140 U23 ( .A1(n6), .A2(n33), .B1(n2), .B2(n58), .ZN(N290)
         );
  NR2D3BWP30P140 U24 ( .A1(n5), .A2(n4), .ZN(n11) );
  ND3D1BWP30P140 U25 ( .A1(n10), .A2(n11), .A3(i_data_bus[40]), .ZN(n12) );
  INVD1BWP30P140 U26 ( .I(i_valid[1]), .ZN(n3) );
  OAI22OPTPBD1BWP30P140 U27 ( .A1(n2), .A2(n56), .B1(n6), .B2(n35), .ZN(N292)
         );
  ND2OPTIBD4BWP30P140 U28 ( .A1(n11), .A2(n10), .ZN(n93) );
  NR2D1BWP30P140 U29 ( .A1(n71), .A2(n53), .ZN(n13) );
  ND2D1BWP30P140 U30 ( .A1(n21), .A2(n20), .ZN(N343) );
  ND2D1BWP30P140 U31 ( .A1(n41), .A2(i_data_bus[24]), .ZN(n21) );
  ND2D1BWP30P140 U32 ( .A1(n69), .A2(i_data_bus[56]), .ZN(n20) );
  IND2D1BWP30P140 U33 ( .A1(n15), .B1(n2), .ZN(N353) );
  NR3D0BWP30P140 U34 ( .A1(n3), .A2(n14), .A3(n16), .ZN(n15) );
  INVD1BWP30P140 U35 ( .I(n69), .ZN(n25) );
  INVD1BWP30P140 U36 ( .I(n16), .ZN(n9) );
  INVD1BWP30P140 U37 ( .I(n23), .ZN(n24) );
  INVD1BWP30P140 U38 ( .I(rst), .ZN(n7) );
  ND2D1BWP30P140 U39 ( .A1(n7), .A2(i_en), .ZN(n16) );
  CKND2D2BWP30P140 U40 ( .A1(i_valid[0]), .A2(n9), .ZN(n8) );
  IND2D1BWP30P140 U41 ( .A1(n13), .B1(n12), .ZN(N295) );
  INVD2BWP30P140 U42 ( .I(i_cmd[1]), .ZN(n23) );
  MUX2NOPTD2BWP30P140 U43 ( .I0(i_valid[0]), .I1(i_valid[1]), .S(i_cmd[0]), 
        .ZN(n17) );
  NR2OPTPAD4BWP30P140 U44 ( .A1(n17), .A2(n18), .ZN(n41) );
  ND2OPTIBD4BWP30P140 U45 ( .A1(i_cmd[1]), .A2(n9), .ZN(n19) );
  INR2D8BWP30P140 U46 ( .A1(i_valid[1]), .B1(n19), .ZN(n69) );
  INVD1BWP30P140 U47 ( .I(n22), .ZN(n26) );
  OAI21D1BWP30P140 U48 ( .A1(n26), .A2(n24), .B(n25), .ZN(N354) );
  INVD1BWP30P140 U49 ( .I(i_data_bus[17]), .ZN(n47) );
  INVD1BWP30P140 U50 ( .I(i_data_bus[49]), .ZN(n27) );
  INVD1BWP30P140 U51 ( .I(i_data_bus[18]), .ZN(n45) );
  INVD1BWP30P140 U52 ( .I(i_data_bus[50]), .ZN(n28) );
  INVD1BWP30P140 U53 ( .I(i_data_bus[19]), .ZN(n44) );
  INVD1BWP30P140 U54 ( .I(i_data_bus[51]), .ZN(n29) );
  INVD1BWP30P140 U55 ( .I(i_data_bus[29]), .ZN(n65) );
  INVD1BWP30P140 U56 ( .I(i_data_bus[61]), .ZN(n30) );
  INVD1BWP30P140 U57 ( .I(i_data_bus[30]), .ZN(n64) );
  INVD1BWP30P140 U58 ( .I(i_data_bus[62]), .ZN(n31) );
  INVD1BWP30P140 U59 ( .I(i_data_bus[31]), .ZN(n63) );
  INVD1BWP30P140 U60 ( .I(i_data_bus[63]), .ZN(n32) );
  INVD1BWP30P140 U61 ( .I(i_data_bus[3]), .ZN(n58) );
  INVD1BWP30P140 U62 ( .I(i_data_bus[35]), .ZN(n33) );
  INVD1BWP30P140 U63 ( .I(i_data_bus[4]), .ZN(n57) );
  INVD1BWP30P140 U64 ( .I(i_data_bus[36]), .ZN(n34) );
  INVD1BWP30P140 U65 ( .I(i_data_bus[5]), .ZN(n56) );
  INVD1BWP30P140 U66 ( .I(i_data_bus[37]), .ZN(n35) );
  INVD1BWP30P140 U67 ( .I(i_data_bus[6]), .ZN(n55) );
  INVD1BWP30P140 U68 ( .I(i_data_bus[38]), .ZN(n36) );
  INVD1BWP30P140 U69 ( .I(i_data_bus[7]), .ZN(n54) );
  INVD1BWP30P140 U70 ( .I(i_data_bus[39]), .ZN(n37) );
  INVD1BWP30P140 U71 ( .I(i_data_bus[20]), .ZN(n38) );
  MOAI22D1BWP30P140 U72 ( .A1(n38), .A2(n1), .B1(i_data_bus[52]), .B2(n69), 
        .ZN(N339) );
  INVD1BWP30P140 U73 ( .I(i_data_bus[21]), .ZN(n39) );
  MOAI22D1BWP30P140 U74 ( .A1(n39), .A2(n1), .B1(i_data_bus[53]), .B2(n69), 
        .ZN(N340) );
  INVD1BWP30P140 U75 ( .I(i_data_bus[15]), .ZN(n40) );
  MOAI22D1BWP30P140 U76 ( .A1(n40), .A2(n1), .B1(i_data_bus[47]), .B2(n69), 
        .ZN(N334) );
  INVD1BWP30P140 U77 ( .I(i_data_bus[14]), .ZN(n42) );
  MOAI22D1BWP30P140 U78 ( .A1(n42), .A2(n1), .B1(i_data_bus[46]), .B2(n69), 
        .ZN(N333) );
  INVD1BWP30P140 U79 ( .I(i_data_bus[16]), .ZN(n43) );
  MOAI22D1BWP30P140 U80 ( .A1(n43), .A2(n1), .B1(i_data_bus[48]), .B2(n69), 
        .ZN(N335) );
  MOAI22D1BWP30P140 U81 ( .A1(n44), .A2(n1), .B1(i_data_bus[51]), .B2(n69), 
        .ZN(N338) );
  MOAI22D1BWP30P140 U82 ( .A1(n45), .A2(n1), .B1(i_data_bus[50]), .B2(n69), 
        .ZN(N337) );
  INVD1BWP30P140 U83 ( .I(i_data_bus[22]), .ZN(n46) );
  MOAI22D1BWP30P140 U84 ( .A1(n46), .A2(n1), .B1(i_data_bus[54]), .B2(n69), 
        .ZN(N341) );
  MOAI22D1BWP30P140 U85 ( .A1(n47), .A2(n1), .B1(i_data_bus[49]), .B2(n69), 
        .ZN(N336) );
  INVD1BWP30P140 U86 ( .I(i_data_bus[23]), .ZN(n48) );
  MOAI22D1BWP30P140 U87 ( .A1(n48), .A2(n1), .B1(i_data_bus[55]), .B2(n69), 
        .ZN(N342) );
  INVD1BWP30P140 U88 ( .I(i_data_bus[13]), .ZN(n49) );
  MOAI22D1BWP30P140 U89 ( .A1(n49), .A2(n1), .B1(i_data_bus[45]), .B2(n69), 
        .ZN(N332) );
  INVD1BWP30P140 U90 ( .I(i_data_bus[11]), .ZN(n50) );
  MOAI22D1BWP30P140 U91 ( .A1(n50), .A2(n1), .B1(i_data_bus[43]), .B2(n69), 
        .ZN(N330) );
  INVD1BWP30P140 U92 ( .I(i_data_bus[10]), .ZN(n51) );
  MOAI22D1BWP30P140 U93 ( .A1(n51), .A2(n1), .B1(i_data_bus[42]), .B2(n69), 
        .ZN(N329) );
  INVD1BWP30P140 U94 ( .I(i_data_bus[9]), .ZN(n52) );
  MOAI22D1BWP30P140 U95 ( .A1(n52), .A2(n1), .B1(i_data_bus[41]), .B2(n69), 
        .ZN(N328) );
  INVD1BWP30P140 U96 ( .I(i_data_bus[8]), .ZN(n53) );
  MOAI22D1BWP30P140 U97 ( .A1(n53), .A2(n1), .B1(i_data_bus[40]), .B2(n69), 
        .ZN(N327) );
  MOAI22D1BWP30P140 U98 ( .A1(n54), .A2(n1), .B1(i_data_bus[39]), .B2(n69), 
        .ZN(N326) );
  MOAI22D1BWP30P140 U99 ( .A1(n55), .A2(n1), .B1(i_data_bus[38]), .B2(n69), 
        .ZN(N325) );
  MOAI22D1BWP30P140 U100 ( .A1(n56), .A2(n1), .B1(i_data_bus[37]), .B2(n69), 
        .ZN(N324) );
  MOAI22D1BWP30P140 U101 ( .A1(n57), .A2(n1), .B1(i_data_bus[36]), .B2(n69), 
        .ZN(N323) );
  MOAI22D1BWP30P140 U102 ( .A1(n58), .A2(n1), .B1(i_data_bus[35]), .B2(n69), 
        .ZN(N322) );
  INVD1BWP30P140 U103 ( .I(i_data_bus[2]), .ZN(n59) );
  MOAI22D1BWP30P140 U104 ( .A1(n59), .A2(n1), .B1(i_data_bus[34]), .B2(n69), 
        .ZN(N321) );
  INVD1BWP30P140 U105 ( .I(i_data_bus[1]), .ZN(n60) );
  MOAI22D1BWP30P140 U106 ( .A1(n60), .A2(n1), .B1(i_data_bus[33]), .B2(n69), 
        .ZN(N320) );
  INVD1BWP30P140 U107 ( .I(i_data_bus[0]), .ZN(n61) );
  MOAI22D1BWP30P140 U108 ( .A1(n61), .A2(n1), .B1(i_data_bus[32]), .B2(n69), 
        .ZN(N319) );
  INVD1BWP30P140 U109 ( .I(i_data_bus[12]), .ZN(n62) );
  MOAI22D1BWP30P140 U110 ( .A1(n62), .A2(n1), .B1(i_data_bus[44]), .B2(n69), 
        .ZN(N331) );
  MOAI22D1BWP30P140 U111 ( .A1(n63), .A2(n1), .B1(i_data_bus[63]), .B2(n69), 
        .ZN(N350) );
  MOAI22D1BWP30P140 U112 ( .A1(n64), .A2(n1), .B1(i_data_bus[62]), .B2(n69), 
        .ZN(N349) );
  MOAI22D1BWP30P140 U113 ( .A1(n65), .A2(n1), .B1(i_data_bus[61]), .B2(n69), 
        .ZN(N348) );
  INVD1BWP30P140 U114 ( .I(i_data_bus[28]), .ZN(n66) );
  MOAI22D1BWP30P140 U115 ( .A1(n66), .A2(n1), .B1(i_data_bus[60]), .B2(n69), 
        .ZN(N347) );
  INVD1BWP30P140 U116 ( .I(i_data_bus[27]), .ZN(n67) );
  MOAI22D1BWP30P140 U117 ( .A1(n67), .A2(n1), .B1(i_data_bus[59]), .B2(n69), 
        .ZN(N346) );
  INVD1BWP30P140 U118 ( .I(i_data_bus[26]), .ZN(n68) );
  MOAI22D1BWP30P140 U119 ( .A1(n68), .A2(n1), .B1(i_data_bus[58]), .B2(n69), 
        .ZN(N345) );
  INVD1BWP30P140 U120 ( .I(i_data_bus[25]), .ZN(n70) );
  MOAI22D1BWP30P140 U121 ( .A1(n70), .A2(n1), .B1(i_data_bus[57]), .B2(n69), 
        .ZN(N344) );
  INVD1BWP30P140 U122 ( .I(i_data_bus[60]), .ZN(n72) );
  MOAI22D1BWP30P140 U123 ( .A1(n6), .A2(n72), .B1(n91), .B2(i_data_bus[28]), 
        .ZN(N315) );
  INVD1BWP30P140 U124 ( .I(i_data_bus[48]), .ZN(n73) );
  MOAI22D1BWP30P140 U125 ( .A1(n6), .A2(n73), .B1(n91), .B2(i_data_bus[16]), 
        .ZN(N303) );
  INVD1BWP30P140 U126 ( .I(i_data_bus[34]), .ZN(n74) );
  MOAI22D1BWP30P140 U127 ( .A1(n93), .A2(n74), .B1(n91), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140 U128 ( .I(i_data_bus[59]), .ZN(n75) );
  MOAI22D1BWP30P140 U129 ( .A1(n6), .A2(n75), .B1(n91), .B2(i_data_bus[27]), 
        .ZN(N314) );
  INVD1BWP30P140 U130 ( .I(i_data_bus[47]), .ZN(n76) );
  MOAI22D1BWP30P140 U131 ( .A1(n93), .A2(n76), .B1(n91), .B2(i_data_bus[15]), 
        .ZN(N302) );
  INVD1BWP30P140 U132 ( .I(i_data_bus[33]), .ZN(n77) );
  MOAI22D1BWP30P140 U133 ( .A1(n6), .A2(n77), .B1(n91), .B2(i_data_bus[1]), 
        .ZN(N288) );
  INVD1BWP30P140 U134 ( .I(i_data_bus[58]), .ZN(n78) );
  MOAI22D1BWP30P140 U135 ( .A1(n93), .A2(n78), .B1(n91), .B2(i_data_bus[26]), 
        .ZN(N313) );
  INVD1BWP30P140 U136 ( .I(i_data_bus[46]), .ZN(n79) );
  MOAI22D1BWP30P140 U137 ( .A1(n93), .A2(n79), .B1(n91), .B2(i_data_bus[14]), 
        .ZN(N301) );
  INVD1BWP30P140 U138 ( .I(i_data_bus[32]), .ZN(n80) );
  MOAI22D1BWP30P140 U139 ( .A1(n93), .A2(n80), .B1(n91), .B2(i_data_bus[0]), 
        .ZN(N287) );
  INVD1BWP30P140 U140 ( .I(i_data_bus[57]), .ZN(n81) );
  MOAI22D1BWP30P140 U141 ( .A1(n6), .A2(n81), .B1(n91), .B2(i_data_bus[25]), 
        .ZN(N312) );
  INVD1BWP30P140 U142 ( .I(i_data_bus[45]), .ZN(n82) );
  MOAI22D1BWP30P140 U143 ( .A1(n93), .A2(n82), .B1(n91), .B2(i_data_bus[13]), 
        .ZN(N300) );
  INVD1BWP30P140 U144 ( .I(i_data_bus[56]), .ZN(n83) );
  MOAI22D1BWP30P140 U145 ( .A1(n6), .A2(n83), .B1(n91), .B2(i_data_bus[24]), 
        .ZN(N311) );
  INVD1BWP30P140 U146 ( .I(i_data_bus[44]), .ZN(n84) );
  MOAI22D1BWP30P140 U147 ( .A1(n93), .A2(n84), .B1(n91), .B2(i_data_bus[12]), 
        .ZN(N299) );
  INVD1BWP30P140 U148 ( .I(i_data_bus[55]), .ZN(n85) );
  MOAI22D1BWP30P140 U149 ( .A1(n6), .A2(n85), .B1(n91), .B2(i_data_bus[23]), 
        .ZN(N310) );
  INVD1BWP30P140 U150 ( .I(i_data_bus[43]), .ZN(n86) );
  MOAI22D1BWP30P140 U151 ( .A1(n93), .A2(n86), .B1(n91), .B2(i_data_bus[11]), 
        .ZN(N298) );
  INVD1BWP30P140 U152 ( .I(i_data_bus[54]), .ZN(n87) );
  MOAI22D1BWP30P140 U153 ( .A1(n6), .A2(n87), .B1(n91), .B2(i_data_bus[22]), 
        .ZN(N309) );
  INVD1BWP30P140 U154 ( .I(i_data_bus[42]), .ZN(n88) );
  MOAI22D1BWP30P140 U155 ( .A1(n93), .A2(n88), .B1(n91), .B2(i_data_bus[10]), 
        .ZN(N297) );
  INVD1BWP30P140 U156 ( .I(i_data_bus[53]), .ZN(n89) );
  MOAI22D1BWP30P140 U157 ( .A1(n6), .A2(n89), .B1(n91), .B2(i_data_bus[21]), 
        .ZN(N308) );
  INVD1BWP30P140 U158 ( .I(i_data_bus[41]), .ZN(n90) );
  MOAI22D1BWP30P140 U159 ( .A1(n93), .A2(n90), .B1(n91), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140 U160 ( .I(i_data_bus[52]), .ZN(n92) );
  MOAI22D1BWP30P140 U161 ( .A1(n6), .A2(n92), .B1(n91), .B2(i_data_bus[20]), 
        .ZN(N307) );
endmodule


module benes_simple_seq ( clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, 
        i_en, i_cmd );
  input [31:0] i_valid;
  input [1023:0] i_data_bus;
  output [31:0] o_valid;
  output [1023:0] o_data_bus;
  input [287:0] i_cmd;
  input clk, rst, i_en;
  wire   n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, connection_0__0__31_,
         connection_0__0__30_, connection_0__0__29_, connection_0__0__28_,
         connection_0__0__27_, connection_0__0__26_, connection_0__0__25_,
         connection_0__0__24_, connection_0__0__23_, connection_0__0__22_,
         connection_0__0__21_, connection_0__0__20_, connection_0__0__19_,
         connection_0__0__18_, connection_0__0__17_, connection_0__0__16_,
         connection_0__0__15_, connection_0__0__14_, connection_0__0__13_,
         connection_0__0__12_, connection_0__0__11_, connection_0__0__10_,
         connection_0__0__9_, connection_0__0__8_, connection_0__0__7_,
         connection_0__0__6_, connection_0__0__5_, connection_0__0__4_,
         connection_0__0__3_, connection_0__0__2_, connection_0__0__1_,
         connection_0__0__0_, connection_0__1__31_, connection_0__1__30_,
         connection_0__1__29_, connection_0__1__28_, connection_0__1__27_,
         connection_0__1__26_, connection_0__1__25_, connection_0__1__24_,
         connection_0__1__23_, connection_0__1__22_, connection_0__1__21_,
         connection_0__1__20_, connection_0__1__19_, connection_0__1__18_,
         connection_0__1__17_, connection_0__1__16_, connection_0__1__15_,
         connection_0__1__14_, connection_0__1__13_, connection_0__1__12_,
         connection_0__1__11_, connection_0__1__10_, connection_0__1__9_,
         connection_0__1__8_, connection_0__1__7_, connection_0__1__6_,
         connection_0__1__5_, connection_0__1__4_, connection_0__1__3_,
         connection_0__1__2_, connection_0__1__1_, connection_0__1__0_,
         connection_0__2__31_, connection_0__2__30_, connection_0__2__29_,
         connection_0__2__28_, connection_0__2__27_, connection_0__2__26_,
         connection_0__2__25_, connection_0__2__24_, connection_0__2__23_,
         connection_0__2__22_, connection_0__2__21_, connection_0__2__20_,
         connection_0__2__19_, connection_0__2__18_, connection_0__2__17_,
         connection_0__2__16_, connection_0__2__15_, connection_0__2__14_,
         connection_0__2__13_, connection_0__2__12_, connection_0__2__11_,
         connection_0__2__10_, connection_0__2__9_, connection_0__2__8_,
         connection_0__2__7_, connection_0__2__6_, connection_0__2__5_,
         connection_0__2__4_, connection_0__2__3_, connection_0__2__2_,
         connection_0__2__1_, connection_0__2__0_, connection_0__3__31_,
         connection_0__3__30_, connection_0__3__29_, connection_0__3__28_,
         connection_0__3__27_, connection_0__3__26_, connection_0__3__25_,
         connection_0__3__24_, connection_0__3__23_, connection_0__3__22_,
         connection_0__3__21_, connection_0__3__20_, connection_0__3__19_,
         connection_0__3__18_, connection_0__3__17_, connection_0__3__16_,
         connection_0__3__15_, connection_0__3__14_, connection_0__3__13_,
         connection_0__3__12_, connection_0__3__11_, connection_0__3__10_,
         connection_0__3__9_, connection_0__3__8_, connection_0__3__7_,
         connection_0__3__6_, connection_0__3__5_, connection_0__3__4_,
         connection_0__3__3_, connection_0__3__2_, connection_0__3__1_,
         connection_0__3__0_, connection_0__4__31_, connection_0__4__30_,
         connection_0__4__29_, connection_0__4__28_, connection_0__4__27_,
         connection_0__4__26_, connection_0__4__25_, connection_0__4__24_,
         connection_0__4__23_, connection_0__4__22_, connection_0__4__21_,
         connection_0__4__20_, connection_0__4__19_, connection_0__4__18_,
         connection_0__4__17_, connection_0__4__16_, connection_0__4__15_,
         connection_0__4__14_, connection_0__4__13_, connection_0__4__12_,
         connection_0__4__11_, connection_0__4__10_, connection_0__4__9_,
         connection_0__4__8_, connection_0__4__7_, connection_0__4__6_,
         connection_0__4__5_, connection_0__4__4_, connection_0__4__3_,
         connection_0__4__2_, connection_0__4__1_, connection_0__4__0_,
         connection_0__5__31_, connection_0__5__30_, connection_0__5__29_,
         connection_0__5__28_, connection_0__5__27_, connection_0__5__26_,
         connection_0__5__25_, connection_0__5__24_, connection_0__5__23_,
         connection_0__5__22_, connection_0__5__21_, connection_0__5__20_,
         connection_0__5__19_, connection_0__5__18_, connection_0__5__17_,
         connection_0__5__16_, connection_0__5__15_, connection_0__5__14_,
         connection_0__5__13_, connection_0__5__12_, connection_0__5__11_,
         connection_0__5__10_, connection_0__5__9_, connection_0__5__8_,
         connection_0__5__7_, connection_0__5__6_, connection_0__5__5_,
         connection_0__5__4_, connection_0__5__3_, connection_0__5__2_,
         connection_0__5__1_, connection_0__5__0_, connection_0__6__31_,
         connection_0__6__30_, connection_0__6__29_, connection_0__6__28_,
         connection_0__6__27_, connection_0__6__26_, connection_0__6__25_,
         connection_0__6__24_, connection_0__6__23_, connection_0__6__22_,
         connection_0__6__21_, connection_0__6__20_, connection_0__6__19_,
         connection_0__6__18_, connection_0__6__17_, connection_0__6__16_,
         connection_0__6__15_, connection_0__6__14_, connection_0__6__13_,
         connection_0__6__12_, connection_0__6__11_, connection_0__6__10_,
         connection_0__6__9_, connection_0__6__8_, connection_0__6__7_,
         connection_0__6__6_, connection_0__6__5_, connection_0__6__4_,
         connection_0__6__3_, connection_0__6__2_, connection_0__6__1_,
         connection_0__6__0_, connection_0__7__31_, connection_0__7__30_,
         connection_0__7__29_, connection_0__7__28_, connection_0__7__27_,
         connection_0__7__26_, connection_0__7__25_, connection_0__7__24_,
         connection_0__7__23_, connection_0__7__22_, connection_0__7__21_,
         connection_0__7__20_, connection_0__7__19_, connection_0__7__18_,
         connection_0__7__17_, connection_0__7__16_, connection_0__7__15_,
         connection_0__7__14_, connection_0__7__13_, connection_0__7__12_,
         connection_0__7__11_, connection_0__7__10_, connection_0__7__9_,
         connection_0__7__8_, connection_0__7__7_, connection_0__7__6_,
         connection_0__7__5_, connection_0__7__4_, connection_0__7__3_,
         connection_0__7__2_, connection_0__7__1_, connection_0__7__0_,
         connection_0__8__31_, connection_0__8__30_, connection_0__8__29_,
         connection_0__8__28_, connection_0__8__27_, connection_0__8__26_,
         connection_0__8__25_, connection_0__8__24_, connection_0__8__23_,
         connection_0__8__22_, connection_0__8__21_, connection_0__8__20_,
         connection_0__8__19_, connection_0__8__18_, connection_0__8__17_,
         connection_0__8__16_, connection_0__8__15_, connection_0__8__14_,
         connection_0__8__13_, connection_0__8__12_, connection_0__8__11_,
         connection_0__8__10_, connection_0__8__9_, connection_0__8__8_,
         connection_0__8__7_, connection_0__8__6_, connection_0__8__5_,
         connection_0__8__4_, connection_0__8__3_, connection_0__8__2_,
         connection_0__8__1_, connection_0__8__0_, connection_0__9__31_,
         connection_0__9__30_, connection_0__9__29_, connection_0__9__28_,
         connection_0__9__27_, connection_0__9__26_, connection_0__9__25_,
         connection_0__9__24_, connection_0__9__23_, connection_0__9__22_,
         connection_0__9__21_, connection_0__9__20_, connection_0__9__19_,
         connection_0__9__18_, connection_0__9__17_, connection_0__9__16_,
         connection_0__9__15_, connection_0__9__14_, connection_0__9__13_,
         connection_0__9__12_, connection_0__9__11_, connection_0__9__10_,
         connection_0__9__9_, connection_0__9__8_, connection_0__9__7_,
         connection_0__9__6_, connection_0__9__5_, connection_0__9__4_,
         connection_0__9__3_, connection_0__9__2_, connection_0__9__1_,
         connection_0__9__0_, connection_0__10__31_, connection_0__10__30_,
         connection_0__10__29_, connection_0__10__28_, connection_0__10__27_,
         connection_0__10__26_, connection_0__10__25_, connection_0__10__24_,
         connection_0__10__23_, connection_0__10__22_, connection_0__10__21_,
         connection_0__10__20_, connection_0__10__19_, connection_0__10__18_,
         connection_0__10__17_, connection_0__10__16_, connection_0__10__15_,
         connection_0__10__14_, connection_0__10__13_, connection_0__10__12_,
         connection_0__10__11_, connection_0__10__10_, connection_0__10__9_,
         connection_0__10__8_, connection_0__10__7_, connection_0__10__6_,
         connection_0__10__5_, connection_0__10__4_, connection_0__10__3_,
         connection_0__10__2_, connection_0__10__1_, connection_0__10__0_,
         connection_0__11__31_, connection_0__11__30_, connection_0__11__29_,
         connection_0__11__28_, connection_0__11__27_, connection_0__11__26_,
         connection_0__11__25_, connection_0__11__24_, connection_0__11__23_,
         connection_0__11__22_, connection_0__11__21_, connection_0__11__20_,
         connection_0__11__19_, connection_0__11__18_, connection_0__11__17_,
         connection_0__11__16_, connection_0__11__15_, connection_0__11__14_,
         connection_0__11__13_, connection_0__11__12_, connection_0__11__11_,
         connection_0__11__10_, connection_0__11__9_, connection_0__11__8_,
         connection_0__11__7_, connection_0__11__6_, connection_0__11__5_,
         connection_0__11__4_, connection_0__11__3_, connection_0__11__2_,
         connection_0__11__1_, connection_0__11__0_, connection_0__12__31_,
         connection_0__12__30_, connection_0__12__29_, connection_0__12__28_,
         connection_0__12__27_, connection_0__12__26_, connection_0__12__25_,
         connection_0__12__24_, connection_0__12__23_, connection_0__12__22_,
         connection_0__12__21_, connection_0__12__20_, connection_0__12__19_,
         connection_0__12__18_, connection_0__12__17_, connection_0__12__16_,
         connection_0__12__15_, connection_0__12__14_, connection_0__12__13_,
         connection_0__12__12_, connection_0__12__11_, connection_0__12__10_,
         connection_0__12__9_, connection_0__12__8_, connection_0__12__7_,
         connection_0__12__6_, connection_0__12__5_, connection_0__12__4_,
         connection_0__12__3_, connection_0__12__2_, connection_0__12__1_,
         connection_0__12__0_, connection_0__13__31_, connection_0__13__30_,
         connection_0__13__29_, connection_0__13__28_, connection_0__13__27_,
         connection_0__13__26_, connection_0__13__25_, connection_0__13__24_,
         connection_0__13__23_, connection_0__13__22_, connection_0__13__21_,
         connection_0__13__20_, connection_0__13__19_, connection_0__13__18_,
         connection_0__13__17_, connection_0__13__16_, connection_0__13__15_,
         connection_0__13__14_, connection_0__13__13_, connection_0__13__12_,
         connection_0__13__11_, connection_0__13__10_, connection_0__13__9_,
         connection_0__13__8_, connection_0__13__7_, connection_0__13__6_,
         connection_0__13__5_, connection_0__13__4_, connection_0__13__3_,
         connection_0__13__2_, connection_0__13__1_, connection_0__13__0_,
         connection_0__14__31_, connection_0__14__30_, connection_0__14__29_,
         connection_0__14__28_, connection_0__14__27_, connection_0__14__26_,
         connection_0__14__25_, connection_0__14__24_, connection_0__14__23_,
         connection_0__14__22_, connection_0__14__21_, connection_0__14__20_,
         connection_0__14__19_, connection_0__14__18_, connection_0__14__17_,
         connection_0__14__16_, connection_0__14__15_, connection_0__14__14_,
         connection_0__14__13_, connection_0__14__12_, connection_0__14__11_,
         connection_0__14__10_, connection_0__14__9_, connection_0__14__8_,
         connection_0__14__7_, connection_0__14__6_, connection_0__14__5_,
         connection_0__14__4_, connection_0__14__3_, connection_0__14__2_,
         connection_0__14__1_, connection_0__14__0_, connection_0__15__31_,
         connection_0__15__30_, connection_0__15__29_, connection_0__15__28_,
         connection_0__15__27_, connection_0__15__26_, connection_0__15__25_,
         connection_0__15__24_, connection_0__15__23_, connection_0__15__22_,
         connection_0__15__21_, connection_0__15__20_, connection_0__15__19_,
         connection_0__15__18_, connection_0__15__17_, connection_0__15__16_,
         connection_0__15__15_, connection_0__15__14_, connection_0__15__13_,
         connection_0__15__12_, connection_0__15__11_, connection_0__15__10_,
         connection_0__15__9_, connection_0__15__8_, connection_0__15__7_,
         connection_0__15__6_, connection_0__15__5_, connection_0__15__4_,
         connection_0__15__3_, connection_0__15__2_, connection_0__15__1_,
         connection_0__15__0_, connection_0__16__31_, connection_0__16__30_,
         connection_0__16__29_, connection_0__16__28_, connection_0__16__27_,
         connection_0__16__26_, connection_0__16__25_, connection_0__16__24_,
         connection_0__16__23_, connection_0__16__22_, connection_0__16__21_,
         connection_0__16__20_, connection_0__16__19_, connection_0__16__18_,
         connection_0__16__17_, connection_0__16__16_, connection_0__16__15_,
         connection_0__16__14_, connection_0__16__13_, connection_0__16__12_,
         connection_0__16__11_, connection_0__16__10_, connection_0__16__9_,
         connection_0__16__8_, connection_0__16__7_, connection_0__16__6_,
         connection_0__16__5_, connection_0__16__4_, connection_0__16__3_,
         connection_0__16__2_, connection_0__16__1_, connection_0__16__0_,
         connection_0__17__31_, connection_0__17__30_, connection_0__17__29_,
         connection_0__17__28_, connection_0__17__27_, connection_0__17__26_,
         connection_0__17__25_, connection_0__17__24_, connection_0__17__23_,
         connection_0__17__22_, connection_0__17__21_, connection_0__17__20_,
         connection_0__17__19_, connection_0__17__18_, connection_0__17__17_,
         connection_0__17__16_, connection_0__17__15_, connection_0__17__14_,
         connection_0__17__13_, connection_0__17__12_, connection_0__17__11_,
         connection_0__17__10_, connection_0__17__9_, connection_0__17__8_,
         connection_0__17__7_, connection_0__17__6_, connection_0__17__5_,
         connection_0__17__4_, connection_0__17__3_, connection_0__17__2_,
         connection_0__17__1_, connection_0__17__0_, connection_0__18__31_,
         connection_0__18__30_, connection_0__18__29_, connection_0__18__28_,
         connection_0__18__27_, connection_0__18__26_, connection_0__18__25_,
         connection_0__18__24_, connection_0__18__23_, connection_0__18__22_,
         connection_0__18__21_, connection_0__18__20_, connection_0__18__19_,
         connection_0__18__18_, connection_0__18__17_, connection_0__18__16_,
         connection_0__18__15_, connection_0__18__14_, connection_0__18__13_,
         connection_0__18__12_, connection_0__18__11_, connection_0__18__10_,
         connection_0__18__9_, connection_0__18__8_, connection_0__18__7_,
         connection_0__18__6_, connection_0__18__5_, connection_0__18__4_,
         connection_0__18__3_, connection_0__18__2_, connection_0__18__1_,
         connection_0__18__0_, connection_0__19__31_, connection_0__19__30_,
         connection_0__19__29_, connection_0__19__28_, connection_0__19__27_,
         connection_0__19__26_, connection_0__19__25_, connection_0__19__24_,
         connection_0__19__23_, connection_0__19__22_, connection_0__19__21_,
         connection_0__19__20_, connection_0__19__19_, connection_0__19__18_,
         connection_0__19__17_, connection_0__19__16_, connection_0__19__15_,
         connection_0__19__14_, connection_0__19__13_, connection_0__19__12_,
         connection_0__19__11_, connection_0__19__10_, connection_0__19__9_,
         connection_0__19__8_, connection_0__19__7_, connection_0__19__6_,
         connection_0__19__5_, connection_0__19__4_, connection_0__19__3_,
         connection_0__19__2_, connection_0__19__1_, connection_0__19__0_,
         connection_0__20__31_, connection_0__20__30_, connection_0__20__29_,
         connection_0__20__28_, connection_0__20__27_, connection_0__20__26_,
         connection_0__20__25_, connection_0__20__24_, connection_0__20__23_,
         connection_0__20__22_, connection_0__20__21_, connection_0__20__20_,
         connection_0__20__19_, connection_0__20__18_, connection_0__20__17_,
         connection_0__20__16_, connection_0__20__15_, connection_0__20__14_,
         connection_0__20__13_, connection_0__20__12_, connection_0__20__11_,
         connection_0__20__10_, connection_0__20__9_, connection_0__20__8_,
         connection_0__20__7_, connection_0__20__6_, connection_0__20__5_,
         connection_0__20__4_, connection_0__20__3_, connection_0__20__2_,
         connection_0__20__1_, connection_0__20__0_, connection_0__21__31_,
         connection_0__21__30_, connection_0__21__29_, connection_0__21__28_,
         connection_0__21__27_, connection_0__21__26_, connection_0__21__25_,
         connection_0__21__24_, connection_0__21__23_, connection_0__21__22_,
         connection_0__21__21_, connection_0__21__20_, connection_0__21__19_,
         connection_0__21__18_, connection_0__21__17_, connection_0__21__16_,
         connection_0__21__15_, connection_0__21__14_, connection_0__21__13_,
         connection_0__21__12_, connection_0__21__11_, connection_0__21__10_,
         connection_0__21__9_, connection_0__21__8_, connection_0__21__7_,
         connection_0__21__6_, connection_0__21__5_, connection_0__21__4_,
         connection_0__21__3_, connection_0__21__2_, connection_0__21__1_,
         connection_0__21__0_, connection_0__22__31_, connection_0__22__30_,
         connection_0__22__29_, connection_0__22__28_, connection_0__22__27_,
         connection_0__22__26_, connection_0__22__25_, connection_0__22__24_,
         connection_0__22__23_, connection_0__22__22_, connection_0__22__21_,
         connection_0__22__20_, connection_0__22__19_, connection_0__22__18_,
         connection_0__22__17_, connection_0__22__16_, connection_0__22__15_,
         connection_0__22__14_, connection_0__22__13_, connection_0__22__12_,
         connection_0__22__11_, connection_0__22__10_, connection_0__22__9_,
         connection_0__22__8_, connection_0__22__7_, connection_0__22__6_,
         connection_0__22__5_, connection_0__22__4_, connection_0__22__3_,
         connection_0__22__2_, connection_0__22__1_, connection_0__22__0_,
         connection_0__23__31_, connection_0__23__30_, connection_0__23__29_,
         connection_0__23__28_, connection_0__23__27_, connection_0__23__26_,
         connection_0__23__25_, connection_0__23__24_, connection_0__23__23_,
         connection_0__23__22_, connection_0__23__21_, connection_0__23__20_,
         connection_0__23__19_, connection_0__23__18_, connection_0__23__17_,
         connection_0__23__16_, connection_0__23__15_, connection_0__23__14_,
         connection_0__23__13_, connection_0__23__12_, connection_0__23__11_,
         connection_0__23__10_, connection_0__23__9_, connection_0__23__8_,
         connection_0__23__7_, connection_0__23__6_, connection_0__23__5_,
         connection_0__23__4_, connection_0__23__3_, connection_0__23__2_,
         connection_0__23__1_, connection_0__23__0_, connection_0__24__31_,
         connection_0__24__30_, connection_0__24__29_, connection_0__24__28_,
         connection_0__24__27_, connection_0__24__26_, connection_0__24__25_,
         connection_0__24__24_, connection_0__24__23_, connection_0__24__22_,
         connection_0__24__21_, connection_0__24__20_, connection_0__24__19_,
         connection_0__24__18_, connection_0__24__17_, connection_0__24__16_,
         connection_0__24__15_, connection_0__24__14_, connection_0__24__13_,
         connection_0__24__12_, connection_0__24__11_, connection_0__24__10_,
         connection_0__24__9_, connection_0__24__8_, connection_0__24__7_,
         connection_0__24__6_, connection_0__24__5_, connection_0__24__4_,
         connection_0__24__3_, connection_0__24__2_, connection_0__24__1_,
         connection_0__24__0_, connection_0__25__31_, connection_0__25__30_,
         connection_0__25__29_, connection_0__25__28_, connection_0__25__27_,
         connection_0__25__26_, connection_0__25__25_, connection_0__25__24_,
         connection_0__25__23_, connection_0__25__22_, connection_0__25__21_,
         connection_0__25__20_, connection_0__25__19_, connection_0__25__18_,
         connection_0__25__17_, connection_0__25__16_, connection_0__25__15_,
         connection_0__25__14_, connection_0__25__13_, connection_0__25__12_,
         connection_0__25__11_, connection_0__25__10_, connection_0__25__9_,
         connection_0__25__8_, connection_0__25__7_, connection_0__25__6_,
         connection_0__25__5_, connection_0__25__4_, connection_0__25__3_,
         connection_0__25__2_, connection_0__25__1_, connection_0__25__0_,
         connection_0__26__31_, connection_0__26__30_, connection_0__26__29_,
         connection_0__26__28_, connection_0__26__27_, connection_0__26__26_,
         connection_0__26__25_, connection_0__26__24_, connection_0__26__23_,
         connection_0__26__22_, connection_0__26__21_, connection_0__26__20_,
         connection_0__26__19_, connection_0__26__18_, connection_0__26__17_,
         connection_0__26__16_, connection_0__26__15_, connection_0__26__14_,
         connection_0__26__13_, connection_0__26__12_, connection_0__26__11_,
         connection_0__26__10_, connection_0__26__9_, connection_0__26__8_,
         connection_0__26__7_, connection_0__26__6_, connection_0__26__5_,
         connection_0__26__4_, connection_0__26__3_, connection_0__26__2_,
         connection_0__26__1_, connection_0__26__0_, connection_0__27__31_,
         connection_0__27__30_, connection_0__27__29_, connection_0__27__28_,
         connection_0__27__27_, connection_0__27__26_, connection_0__27__25_,
         connection_0__27__24_, connection_0__27__23_, connection_0__27__22_,
         connection_0__27__21_, connection_0__27__20_, connection_0__27__19_,
         connection_0__27__18_, connection_0__27__17_, connection_0__27__16_,
         connection_0__27__15_, connection_0__27__14_, connection_0__27__13_,
         connection_0__27__12_, connection_0__27__11_, connection_0__27__10_,
         connection_0__27__9_, connection_0__27__8_, connection_0__27__7_,
         connection_0__27__6_, connection_0__27__5_, connection_0__27__4_,
         connection_0__27__3_, connection_0__27__2_, connection_0__27__1_,
         connection_0__27__0_, connection_0__28__31_, connection_0__28__30_,
         connection_0__28__29_, connection_0__28__28_, connection_0__28__27_,
         connection_0__28__26_, connection_0__28__25_, connection_0__28__24_,
         connection_0__28__23_, connection_0__28__22_, connection_0__28__21_,
         connection_0__28__20_, connection_0__28__19_, connection_0__28__18_,
         connection_0__28__17_, connection_0__28__16_, connection_0__28__15_,
         connection_0__28__14_, connection_0__28__13_, connection_0__28__12_,
         connection_0__28__11_, connection_0__28__10_, connection_0__28__9_,
         connection_0__28__8_, connection_0__28__7_, connection_0__28__6_,
         connection_0__28__5_, connection_0__28__4_, connection_0__28__3_,
         connection_0__28__2_, connection_0__28__1_, connection_0__28__0_,
         connection_0__29__31_, connection_0__29__30_, connection_0__29__29_,
         connection_0__29__28_, connection_0__29__27_, connection_0__29__26_,
         connection_0__29__25_, connection_0__29__24_, connection_0__29__23_,
         connection_0__29__22_, connection_0__29__21_, connection_0__29__20_,
         connection_0__29__19_, connection_0__29__18_, connection_0__29__17_,
         connection_0__29__16_, connection_0__29__15_, connection_0__29__14_,
         connection_0__29__13_, connection_0__29__12_, connection_0__29__11_,
         connection_0__29__10_, connection_0__29__9_, connection_0__29__8_,
         connection_0__29__7_, connection_0__29__6_, connection_0__29__5_,
         connection_0__29__4_, connection_0__29__3_, connection_0__29__2_,
         connection_0__29__1_, connection_0__29__0_, connection_0__30__31_,
         connection_0__30__30_, connection_0__30__29_, connection_0__30__28_,
         connection_0__30__27_, connection_0__30__26_, connection_0__30__25_,
         connection_0__30__24_, connection_0__30__23_, connection_0__30__22_,
         connection_0__30__21_, connection_0__30__20_, connection_0__30__19_,
         connection_0__30__18_, connection_0__30__17_, connection_0__30__16_,
         connection_0__30__15_, connection_0__30__14_, connection_0__30__13_,
         connection_0__30__12_, connection_0__30__11_, connection_0__30__10_,
         connection_0__30__9_, connection_0__30__8_, connection_0__30__7_,
         connection_0__30__6_, connection_0__30__5_, connection_0__30__4_,
         connection_0__30__3_, connection_0__30__2_, connection_0__30__1_,
         connection_0__30__0_, connection_0__31__31_, connection_0__31__30_,
         connection_0__31__29_, connection_0__31__28_, connection_0__31__27_,
         connection_0__31__26_, connection_0__31__25_, connection_0__31__24_,
         connection_0__31__23_, connection_0__31__22_, connection_0__31__21_,
         connection_0__31__20_, connection_0__31__19_, connection_0__31__18_,
         connection_0__31__17_, connection_0__31__16_, connection_0__31__15_,
         connection_0__31__14_, connection_0__31__13_, connection_0__31__12_,
         connection_0__31__11_, connection_0__31__10_, connection_0__31__9_,
         connection_0__31__8_, connection_0__31__7_, connection_0__31__6_,
         connection_0__31__5_, connection_0__31__4_, connection_0__31__3_,
         connection_0__31__2_, connection_0__31__1_, connection_0__31__0_,
         connection_valid_0__0_, connection_valid_0__1_,
         connection_valid_0__2_, connection_valid_0__3_,
         connection_valid_0__4_, connection_valid_0__5_,
         connection_valid_0__6_, connection_valid_0__7_,
         connection_valid_0__8_, connection_valid_0__9_,
         connection_valid_0__10_, connection_valid_0__11_,
         connection_valid_0__12_, connection_valid_0__13_,
         connection_valid_0__14_, connection_valid_0__15_,
         connection_valid_0__16_, connection_valid_0__17_,
         connection_valid_0__18_, connection_valid_0__19_,
         connection_valid_0__20_, connection_valid_0__21_,
         connection_valid_0__22_, connection_valid_0__23_,
         connection_valid_0__24_, connection_valid_0__25_,
         connection_valid_0__26_, connection_valid_0__27_,
         connection_valid_0__28_, connection_valid_0__29_,
         connection_valid_0__30_, connection_valid_0__31_,
         connection_valid_1__0_, connection_valid_1__1_,
         connection_valid_1__2_, connection_valid_1__3_,
         connection_valid_1__4_, connection_valid_1__5_,
         connection_valid_1__6_, connection_valid_1__7_,
         connection_valid_1__8_, connection_valid_1__9_,
         connection_valid_1__10_, connection_valid_1__11_,
         connection_valid_1__12_, connection_valid_1__13_,
         connection_valid_1__14_, connection_valid_1__15_,
         connection_valid_1__16_, connection_valid_1__17_,
         connection_valid_1__18_, connection_valid_1__19_,
         connection_valid_1__20_, connection_valid_1__21_,
         connection_valid_1__22_, connection_valid_1__23_,
         connection_valid_1__24_, connection_valid_1__25_,
         connection_valid_1__26_, connection_valid_1__27_,
         connection_valid_1__28_, connection_valid_1__29_,
         connection_valid_1__30_, connection_valid_1__31_,
         connection_valid_2__0_, connection_valid_2__1_,
         connection_valid_2__2_, connection_valid_2__3_,
         connection_valid_2__4_, connection_valid_2__5_,
         connection_valid_2__6_, connection_valid_2__7_,
         connection_valid_2__8_, connection_valid_2__9_,
         connection_valid_2__10_, connection_valid_2__11_,
         connection_valid_2__12_, connection_valid_2__13_,
         connection_valid_2__14_, connection_valid_2__15_,
         connection_valid_2__16_, connection_valid_2__17_,
         connection_valid_2__18_, connection_valid_2__19_,
         connection_valid_2__20_, connection_valid_2__21_,
         connection_valid_2__22_, connection_valid_2__23_,
         connection_valid_2__24_, connection_valid_2__25_,
         connection_valid_2__26_, connection_valid_2__27_,
         connection_valid_2__28_, connection_valid_2__29_,
         connection_valid_2__30_, connection_valid_2__31_,
         connection_valid_3__0_, connection_valid_3__1_,
         connection_valid_3__2_, connection_valid_3__3_,
         connection_valid_3__4_, connection_valid_3__5_,
         connection_valid_3__6_, connection_valid_3__7_,
         connection_valid_3__8_, connection_valid_3__9_,
         connection_valid_3__10_, connection_valid_3__11_,
         connection_valid_3__12_, connection_valid_3__13_,
         connection_valid_3__14_, connection_valid_3__15_,
         connection_valid_3__16_, connection_valid_3__17_,
         connection_valid_3__18_, connection_valid_3__19_,
         connection_valid_3__20_, connection_valid_3__21_,
         connection_valid_3__22_, connection_valid_3__23_,
         connection_valid_3__24_, connection_valid_3__25_,
         connection_valid_3__26_, connection_valid_3__27_,
         connection_valid_3__28_, connection_valid_3__29_,
         connection_valid_3__30_, connection_valid_3__31_,
         connection_valid_4__0_, connection_valid_4__1_,
         connection_valid_4__2_, connection_valid_4__3_,
         connection_valid_4__4_, connection_valid_4__5_,
         connection_valid_4__6_, connection_valid_4__7_,
         connection_valid_4__8_, connection_valid_4__9_,
         connection_valid_4__10_, connection_valid_4__11_,
         connection_valid_4__12_, connection_valid_4__13_,
         connection_valid_4__14_, connection_valid_4__15_,
         connection_valid_4__16_, connection_valid_4__17_,
         connection_valid_4__18_, connection_valid_4__19_,
         connection_valid_4__20_, connection_valid_4__21_,
         connection_valid_4__22_, connection_valid_4__23_,
         connection_valid_4__24_, connection_valid_4__25_,
         connection_valid_4__26_, connection_valid_4__27_,
         connection_valid_4__28_, connection_valid_4__29_,
         connection_valid_4__30_, connection_valid_4__31_,
         connection_valid_5__0_, connection_valid_5__1_,
         connection_valid_5__2_, connection_valid_5__3_,
         connection_valid_5__4_, connection_valid_5__5_,
         connection_valid_5__6_, connection_valid_5__7_,
         connection_valid_5__8_, connection_valid_5__9_,
         connection_valid_5__10_, connection_valid_5__11_,
         connection_valid_5__12_, connection_valid_5__13_,
         connection_valid_5__14_, connection_valid_5__15_,
         connection_valid_5__16_, connection_valid_5__17_,
         connection_valid_5__18_, connection_valid_5__19_,
         connection_valid_5__20_, connection_valid_5__21_,
         connection_valid_5__22_, connection_valid_5__23_,
         connection_valid_5__24_, connection_valid_5__25_,
         connection_valid_5__26_, connection_valid_5__27_,
         connection_valid_5__28_, connection_valid_5__29_,
         connection_valid_5__30_, connection_valid_5__31_,
         connection_valid_6__0_, connection_valid_6__1_,
         connection_valid_6__2_, connection_valid_6__3_,
         connection_valid_6__4_, connection_valid_6__5_,
         connection_valid_6__6_, connection_valid_6__7_,
         connection_valid_6__8_, connection_valid_6__9_,
         connection_valid_6__10_, connection_valid_6__11_,
         connection_valid_6__12_, connection_valid_6__13_,
         connection_valid_6__14_, connection_valid_6__15_,
         connection_valid_6__16_, connection_valid_6__17_,
         connection_valid_6__18_, connection_valid_6__19_,
         connection_valid_6__20_, connection_valid_6__21_,
         connection_valid_6__22_, connection_valid_6__23_,
         connection_valid_6__24_, connection_valid_6__25_,
         connection_valid_6__26_, connection_valid_6__27_,
         connection_valid_6__28_, connection_valid_6__29_,
         connection_valid_6__30_, connection_valid_6__31_,
         connection_valid_7__0_, connection_valid_7__1_,
         connection_valid_7__2_, connection_valid_7__3_,
         connection_valid_7__4_, connection_valid_7__5_,
         connection_valid_7__6_, connection_valid_7__7_,
         connection_valid_7__8_, connection_valid_7__9_,
         connection_valid_7__10_, connection_valid_7__11_,
         connection_valid_7__12_, connection_valid_7__13_,
         connection_valid_7__14_, connection_valid_7__15_,
         connection_valid_7__16_, connection_valid_7__17_,
         connection_valid_7__18_, connection_valid_7__19_,
         connection_valid_7__20_, connection_valid_7__21_,
         connection_valid_7__22_, connection_valid_7__23_,
         connection_valid_7__24_, connection_valid_7__25_,
         connection_valid_7__26_, connection_valid_7__27_,
         connection_valid_7__28_, connection_valid_7__29_,
         connection_valid_7__30_, connection_valid_7__31_,
         connection_1__0__31_, connection_1__0__30_, connection_1__0__29_,
         connection_1__0__28_, connection_1__0__27_, connection_1__0__26_,
         connection_1__0__25_, connection_1__0__24_, connection_1__0__23_,
         connection_1__0__22_, connection_1__0__21_, connection_1__0__20_,
         connection_1__0__19_, connection_1__0__18_, connection_1__0__17_,
         connection_1__0__16_, connection_1__0__15_, connection_1__0__14_,
         connection_1__0__13_, connection_1__0__12_, connection_1__0__11_,
         connection_1__0__10_, connection_1__0__9_, connection_1__0__8_,
         connection_1__0__7_, connection_1__0__6_, connection_1__0__5_,
         connection_1__0__4_, connection_1__0__3_, connection_1__0__2_,
         connection_1__0__1_, connection_1__0__0_, connection_1__1__31_,
         connection_1__1__30_, connection_1__1__29_, connection_1__1__28_,
         connection_1__1__27_, connection_1__1__26_, connection_1__1__25_,
         connection_1__1__24_, connection_1__1__23_, connection_1__1__22_,
         connection_1__1__21_, connection_1__1__20_, connection_1__1__19_,
         connection_1__1__18_, connection_1__1__17_, connection_1__1__16_,
         connection_1__1__15_, connection_1__1__14_, connection_1__1__13_,
         connection_1__1__12_, connection_1__1__11_, connection_1__1__10_,
         connection_1__1__9_, connection_1__1__8_, connection_1__1__7_,
         connection_1__1__6_, connection_1__1__5_, connection_1__1__4_,
         connection_1__1__3_, connection_1__1__2_, connection_1__1__1_,
         connection_1__1__0_, connection_1__2__31_, connection_1__2__30_,
         connection_1__2__29_, connection_1__2__28_, connection_1__2__27_,
         connection_1__2__26_, connection_1__2__25_, connection_1__2__24_,
         connection_1__2__23_, connection_1__2__22_, connection_1__2__21_,
         connection_1__2__20_, connection_1__2__19_, connection_1__2__18_,
         connection_1__2__17_, connection_1__2__16_, connection_1__2__15_,
         connection_1__2__14_, connection_1__2__13_, connection_1__2__12_,
         connection_1__2__11_, connection_1__2__10_, connection_1__2__9_,
         connection_1__2__8_, connection_1__2__7_, connection_1__2__6_,
         connection_1__2__5_, connection_1__2__4_, connection_1__2__3_,
         connection_1__2__2_, connection_1__2__1_, connection_1__2__0_,
         connection_1__3__31_, connection_1__3__30_, connection_1__3__29_,
         connection_1__3__28_, connection_1__3__27_, connection_1__3__26_,
         connection_1__3__25_, connection_1__3__24_, connection_1__3__23_,
         connection_1__3__22_, connection_1__3__21_, connection_1__3__20_,
         connection_1__3__19_, connection_1__3__18_, connection_1__3__17_,
         connection_1__3__16_, connection_1__3__15_, connection_1__3__14_,
         connection_1__3__13_, connection_1__3__12_, connection_1__3__11_,
         connection_1__3__10_, connection_1__3__9_, connection_1__3__8_,
         connection_1__3__7_, connection_1__3__6_, connection_1__3__5_,
         connection_1__3__4_, connection_1__3__3_, connection_1__3__2_,
         connection_1__3__1_, connection_1__3__0_, connection_1__4__31_,
         connection_1__4__30_, connection_1__4__29_, connection_1__4__28_,
         connection_1__4__27_, connection_1__4__26_, connection_1__4__25_,
         connection_1__4__24_, connection_1__4__23_, connection_1__4__22_,
         connection_1__4__21_, connection_1__4__20_, connection_1__4__19_,
         connection_1__4__18_, connection_1__4__17_, connection_1__4__16_,
         connection_1__4__15_, connection_1__4__14_, connection_1__4__13_,
         connection_1__4__12_, connection_1__4__11_, connection_1__4__10_,
         connection_1__4__9_, connection_1__4__8_, connection_1__4__7_,
         connection_1__4__6_, connection_1__4__5_, connection_1__4__4_,
         connection_1__4__3_, connection_1__4__2_, connection_1__4__1_,
         connection_1__4__0_, connection_1__5__31_, connection_1__5__30_,
         connection_1__5__29_, connection_1__5__28_, connection_1__5__27_,
         connection_1__5__26_, connection_1__5__25_, connection_1__5__24_,
         connection_1__5__23_, connection_1__5__22_, connection_1__5__21_,
         connection_1__5__20_, connection_1__5__19_, connection_1__5__18_,
         connection_1__5__17_, connection_1__5__16_, connection_1__5__15_,
         connection_1__5__14_, connection_1__5__13_, connection_1__5__12_,
         connection_1__5__11_, connection_1__5__10_, connection_1__5__9_,
         connection_1__5__8_, connection_1__5__7_, connection_1__5__6_,
         connection_1__5__5_, connection_1__5__4_, connection_1__5__3_,
         connection_1__5__2_, connection_1__5__1_, connection_1__5__0_,
         connection_1__6__31_, connection_1__6__30_, connection_1__6__29_,
         connection_1__6__28_, connection_1__6__27_, connection_1__6__26_,
         connection_1__6__25_, connection_1__6__24_, connection_1__6__23_,
         connection_1__6__22_, connection_1__6__21_, connection_1__6__20_,
         connection_1__6__19_, connection_1__6__18_, connection_1__6__17_,
         connection_1__6__16_, connection_1__6__15_, connection_1__6__14_,
         connection_1__6__13_, connection_1__6__12_, connection_1__6__11_,
         connection_1__6__10_, connection_1__6__9_, connection_1__6__8_,
         connection_1__6__7_, connection_1__6__6_, connection_1__6__5_,
         connection_1__6__4_, connection_1__6__3_, connection_1__6__2_,
         connection_1__6__1_, connection_1__6__0_, connection_1__7__31_,
         connection_1__7__30_, connection_1__7__29_, connection_1__7__28_,
         connection_1__7__27_, connection_1__7__26_, connection_1__7__25_,
         connection_1__7__24_, connection_1__7__23_, connection_1__7__22_,
         connection_1__7__21_, connection_1__7__20_, connection_1__7__19_,
         connection_1__7__18_, connection_1__7__17_, connection_1__7__16_,
         connection_1__7__15_, connection_1__7__14_, connection_1__7__13_,
         connection_1__7__12_, connection_1__7__11_, connection_1__7__10_,
         connection_1__7__9_, connection_1__7__8_, connection_1__7__7_,
         connection_1__7__6_, connection_1__7__5_, connection_1__7__4_,
         connection_1__7__3_, connection_1__7__2_, connection_1__7__1_,
         connection_1__7__0_, connection_1__8__31_, connection_1__8__30_,
         connection_1__8__29_, connection_1__8__28_, connection_1__8__27_,
         connection_1__8__26_, connection_1__8__25_, connection_1__8__24_,
         connection_1__8__23_, connection_1__8__22_, connection_1__8__21_,
         connection_1__8__20_, connection_1__8__19_, connection_1__8__18_,
         connection_1__8__17_, connection_1__8__16_, connection_1__8__15_,
         connection_1__8__14_, connection_1__8__13_, connection_1__8__12_,
         connection_1__8__11_, connection_1__8__10_, connection_1__8__9_,
         connection_1__8__8_, connection_1__8__7_, connection_1__8__6_,
         connection_1__8__5_, connection_1__8__4_, connection_1__8__3_,
         connection_1__8__2_, connection_1__8__1_, connection_1__8__0_,
         connection_1__9__31_, connection_1__9__30_, connection_1__9__29_,
         connection_1__9__28_, connection_1__9__27_, connection_1__9__26_,
         connection_1__9__25_, connection_1__9__24_, connection_1__9__23_,
         connection_1__9__22_, connection_1__9__21_, connection_1__9__20_,
         connection_1__9__19_, connection_1__9__18_, connection_1__9__17_,
         connection_1__9__16_, connection_1__9__15_, connection_1__9__14_,
         connection_1__9__13_, connection_1__9__12_, connection_1__9__11_,
         connection_1__9__10_, connection_1__9__9_, connection_1__9__8_,
         connection_1__9__7_, connection_1__9__6_, connection_1__9__5_,
         connection_1__9__4_, connection_1__9__3_, connection_1__9__2_,
         connection_1__9__1_, connection_1__9__0_, connection_1__10__31_,
         connection_1__10__30_, connection_1__10__29_, connection_1__10__28_,
         connection_1__10__27_, connection_1__10__26_, connection_1__10__25_,
         connection_1__10__24_, connection_1__10__23_, connection_1__10__22_,
         connection_1__10__21_, connection_1__10__20_, connection_1__10__19_,
         connection_1__10__18_, connection_1__10__17_, connection_1__10__16_,
         connection_1__10__15_, connection_1__10__14_, connection_1__10__13_,
         connection_1__10__12_, connection_1__10__11_, connection_1__10__10_,
         connection_1__10__9_, connection_1__10__8_, connection_1__10__7_,
         connection_1__10__6_, connection_1__10__5_, connection_1__10__4_,
         connection_1__10__3_, connection_1__10__2_, connection_1__10__1_,
         connection_1__10__0_, connection_1__11__31_, connection_1__11__30_,
         connection_1__11__29_, connection_1__11__28_, connection_1__11__27_,
         connection_1__11__26_, connection_1__11__25_, connection_1__11__24_,
         connection_1__11__23_, connection_1__11__22_, connection_1__11__21_,
         connection_1__11__20_, connection_1__11__19_, connection_1__11__18_,
         connection_1__11__17_, connection_1__11__16_, connection_1__11__15_,
         connection_1__11__14_, connection_1__11__13_, connection_1__11__12_,
         connection_1__11__11_, connection_1__11__10_, connection_1__11__9_,
         connection_1__11__8_, connection_1__11__7_, connection_1__11__6_,
         connection_1__11__5_, connection_1__11__4_, connection_1__11__3_,
         connection_1__11__2_, connection_1__11__1_, connection_1__11__0_,
         connection_1__12__31_, connection_1__12__30_, connection_1__12__29_,
         connection_1__12__28_, connection_1__12__27_, connection_1__12__26_,
         connection_1__12__25_, connection_1__12__24_, connection_1__12__23_,
         connection_1__12__22_, connection_1__12__21_, connection_1__12__20_,
         connection_1__12__19_, connection_1__12__18_, connection_1__12__17_,
         connection_1__12__16_, connection_1__12__15_, connection_1__12__14_,
         connection_1__12__13_, connection_1__12__12_, connection_1__12__11_,
         connection_1__12__10_, connection_1__12__9_, connection_1__12__8_,
         connection_1__12__7_, connection_1__12__6_, connection_1__12__5_,
         connection_1__12__4_, connection_1__12__3_, connection_1__12__2_,
         connection_1__12__1_, connection_1__12__0_, connection_1__13__31_,
         connection_1__13__30_, connection_1__13__29_, connection_1__13__28_,
         connection_1__13__27_, connection_1__13__26_, connection_1__13__25_,
         connection_1__13__24_, connection_1__13__23_, connection_1__13__22_,
         connection_1__13__21_, connection_1__13__20_, connection_1__13__19_,
         connection_1__13__18_, connection_1__13__17_, connection_1__13__16_,
         connection_1__13__15_, connection_1__13__14_, connection_1__13__13_,
         connection_1__13__12_, connection_1__13__11_, connection_1__13__10_,
         connection_1__13__9_, connection_1__13__8_, connection_1__13__7_,
         connection_1__13__6_, connection_1__13__5_, connection_1__13__4_,
         connection_1__13__3_, connection_1__13__2_, connection_1__13__1_,
         connection_1__13__0_, connection_1__14__31_, connection_1__14__30_,
         connection_1__14__29_, connection_1__14__28_, connection_1__14__27_,
         connection_1__14__26_, connection_1__14__25_, connection_1__14__24_,
         connection_1__14__23_, connection_1__14__22_, connection_1__14__21_,
         connection_1__14__20_, connection_1__14__19_, connection_1__14__18_,
         connection_1__14__17_, connection_1__14__16_, connection_1__14__15_,
         connection_1__14__14_, connection_1__14__13_, connection_1__14__12_,
         connection_1__14__11_, connection_1__14__10_, connection_1__14__9_,
         connection_1__14__8_, connection_1__14__7_, connection_1__14__6_,
         connection_1__14__5_, connection_1__14__4_, connection_1__14__3_,
         connection_1__14__2_, connection_1__14__1_, connection_1__14__0_,
         connection_1__15__31_, connection_1__15__30_, connection_1__15__29_,
         connection_1__15__28_, connection_1__15__27_, connection_1__15__26_,
         connection_1__15__25_, connection_1__15__24_, connection_1__15__23_,
         connection_1__15__22_, connection_1__15__21_, connection_1__15__20_,
         connection_1__15__19_, connection_1__15__18_, connection_1__15__17_,
         connection_1__15__16_, connection_1__15__15_, connection_1__15__14_,
         connection_1__15__13_, connection_1__15__12_, connection_1__15__11_,
         connection_1__15__10_, connection_1__15__9_, connection_1__15__8_,
         connection_1__15__7_, connection_1__15__6_, connection_1__15__5_,
         connection_1__15__4_, connection_1__15__3_, connection_1__15__2_,
         connection_1__15__1_, connection_1__15__0_, connection_1__16__31_,
         connection_1__16__30_, connection_1__16__29_, connection_1__16__28_,
         connection_1__16__27_, connection_1__16__26_, connection_1__16__25_,
         connection_1__16__24_, connection_1__16__23_, connection_1__16__22_,
         connection_1__16__21_, connection_1__16__20_, connection_1__16__19_,
         connection_1__16__18_, connection_1__16__17_, connection_1__16__16_,
         connection_1__16__15_, connection_1__16__14_, connection_1__16__13_,
         connection_1__16__12_, connection_1__16__11_, connection_1__16__10_,
         connection_1__16__9_, connection_1__16__8_, connection_1__16__7_,
         connection_1__16__6_, connection_1__16__5_, connection_1__16__4_,
         connection_1__16__3_, connection_1__16__2_, connection_1__16__1_,
         connection_1__16__0_, connection_1__17__31_, connection_1__17__30_,
         connection_1__17__29_, connection_1__17__28_, connection_1__17__27_,
         connection_1__17__26_, connection_1__17__25_, connection_1__17__24_,
         connection_1__17__23_, connection_1__17__22_, connection_1__17__21_,
         connection_1__17__20_, connection_1__17__19_, connection_1__17__18_,
         connection_1__17__17_, connection_1__17__16_, connection_1__17__15_,
         connection_1__17__14_, connection_1__17__13_, connection_1__17__12_,
         connection_1__17__11_, connection_1__17__10_, connection_1__17__9_,
         connection_1__17__8_, connection_1__17__7_, connection_1__17__6_,
         connection_1__17__5_, connection_1__17__4_, connection_1__17__3_,
         connection_1__17__2_, connection_1__17__1_, connection_1__17__0_,
         connection_1__18__31_, connection_1__18__30_, connection_1__18__29_,
         connection_1__18__28_, connection_1__18__27_, connection_1__18__26_,
         connection_1__18__25_, connection_1__18__24_, connection_1__18__23_,
         connection_1__18__22_, connection_1__18__21_, connection_1__18__20_,
         connection_1__18__19_, connection_1__18__18_, connection_1__18__17_,
         connection_1__18__16_, connection_1__18__15_, connection_1__18__14_,
         connection_1__18__13_, connection_1__18__12_, connection_1__18__11_,
         connection_1__18__10_, connection_1__18__9_, connection_1__18__8_,
         connection_1__18__7_, connection_1__18__6_, connection_1__18__5_,
         connection_1__18__4_, connection_1__18__3_, connection_1__18__2_,
         connection_1__18__1_, connection_1__18__0_, connection_1__19__31_,
         connection_1__19__30_, connection_1__19__29_, connection_1__19__28_,
         connection_1__19__27_, connection_1__19__26_, connection_1__19__25_,
         connection_1__19__24_, connection_1__19__23_, connection_1__19__22_,
         connection_1__19__21_, connection_1__19__20_, connection_1__19__19_,
         connection_1__19__18_, connection_1__19__17_, connection_1__19__16_,
         connection_1__19__15_, connection_1__19__14_, connection_1__19__13_,
         connection_1__19__12_, connection_1__19__11_, connection_1__19__10_,
         connection_1__19__9_, connection_1__19__8_, connection_1__19__7_,
         connection_1__19__6_, connection_1__19__5_, connection_1__19__4_,
         connection_1__19__3_, connection_1__19__2_, connection_1__19__1_,
         connection_1__19__0_, connection_1__20__31_, connection_1__20__30_,
         connection_1__20__29_, connection_1__20__28_, connection_1__20__27_,
         connection_1__20__26_, connection_1__20__25_, connection_1__20__24_,
         connection_1__20__23_, connection_1__20__22_, connection_1__20__21_,
         connection_1__20__20_, connection_1__20__19_, connection_1__20__18_,
         connection_1__20__17_, connection_1__20__16_, connection_1__20__15_,
         connection_1__20__14_, connection_1__20__13_, connection_1__20__12_,
         connection_1__20__11_, connection_1__20__10_, connection_1__20__9_,
         connection_1__20__8_, connection_1__20__7_, connection_1__20__6_,
         connection_1__20__5_, connection_1__20__4_, connection_1__20__3_,
         connection_1__20__2_, connection_1__20__1_, connection_1__20__0_,
         connection_1__21__31_, connection_1__21__30_, connection_1__21__29_,
         connection_1__21__28_, connection_1__21__27_, connection_1__21__26_,
         connection_1__21__25_, connection_1__21__24_, connection_1__21__23_,
         connection_1__21__22_, connection_1__21__21_, connection_1__21__20_,
         connection_1__21__19_, connection_1__21__18_, connection_1__21__17_,
         connection_1__21__16_, connection_1__21__15_, connection_1__21__14_,
         connection_1__21__13_, connection_1__21__12_, connection_1__21__11_,
         connection_1__21__10_, connection_1__21__9_, connection_1__21__8_,
         connection_1__21__7_, connection_1__21__6_, connection_1__21__5_,
         connection_1__21__4_, connection_1__21__3_, connection_1__21__2_,
         connection_1__21__1_, connection_1__21__0_, connection_1__22__31_,
         connection_1__22__30_, connection_1__22__29_, connection_1__22__28_,
         connection_1__22__27_, connection_1__22__26_, connection_1__22__25_,
         connection_1__22__24_, connection_1__22__23_, connection_1__22__22_,
         connection_1__22__21_, connection_1__22__20_, connection_1__22__19_,
         connection_1__22__18_, connection_1__22__17_, connection_1__22__16_,
         connection_1__22__15_, connection_1__22__14_, connection_1__22__13_,
         connection_1__22__12_, connection_1__22__11_, connection_1__22__10_,
         connection_1__22__9_, connection_1__22__8_, connection_1__22__7_,
         connection_1__22__6_, connection_1__22__5_, connection_1__22__4_,
         connection_1__22__3_, connection_1__22__2_, connection_1__22__1_,
         connection_1__22__0_, connection_1__23__31_, connection_1__23__30_,
         connection_1__23__29_, connection_1__23__28_, connection_1__23__27_,
         connection_1__23__26_, connection_1__23__25_, connection_1__23__24_,
         connection_1__23__23_, connection_1__23__22_, connection_1__23__21_,
         connection_1__23__20_, connection_1__23__19_, connection_1__23__18_,
         connection_1__23__17_, connection_1__23__16_, connection_1__23__15_,
         connection_1__23__14_, connection_1__23__13_, connection_1__23__12_,
         connection_1__23__11_, connection_1__23__10_, connection_1__23__9_,
         connection_1__23__8_, connection_1__23__7_, connection_1__23__6_,
         connection_1__23__5_, connection_1__23__4_, connection_1__23__3_,
         connection_1__23__2_, connection_1__23__1_, connection_1__23__0_,
         connection_1__24__31_, connection_1__24__30_, connection_1__24__29_,
         connection_1__24__28_, connection_1__24__27_, connection_1__24__26_,
         connection_1__24__25_, connection_1__24__24_, connection_1__24__23_,
         connection_1__24__22_, connection_1__24__21_, connection_1__24__20_,
         connection_1__24__19_, connection_1__24__18_, connection_1__24__17_,
         connection_1__24__16_, connection_1__24__15_, connection_1__24__14_,
         connection_1__24__13_, connection_1__24__12_, connection_1__24__11_,
         connection_1__24__10_, connection_1__24__9_, connection_1__24__8_,
         connection_1__24__7_, connection_1__24__6_, connection_1__24__5_,
         connection_1__24__4_, connection_1__24__3_, connection_1__24__2_,
         connection_1__24__1_, connection_1__24__0_, connection_1__25__31_,
         connection_1__25__30_, connection_1__25__29_, connection_1__25__28_,
         connection_1__25__27_, connection_1__25__26_, connection_1__25__25_,
         connection_1__25__24_, connection_1__25__23_, connection_1__25__22_,
         connection_1__25__21_, connection_1__25__20_, connection_1__25__19_,
         connection_1__25__18_, connection_1__25__17_, connection_1__25__16_,
         connection_1__25__15_, connection_1__25__14_, connection_1__25__13_,
         connection_1__25__12_, connection_1__25__11_, connection_1__25__10_,
         connection_1__25__9_, connection_1__25__8_, connection_1__25__7_,
         connection_1__25__6_, connection_1__25__5_, connection_1__25__4_,
         connection_1__25__3_, connection_1__25__2_, connection_1__25__1_,
         connection_1__25__0_, connection_1__26__31_, connection_1__26__30_,
         connection_1__26__29_, connection_1__26__28_, connection_1__26__27_,
         connection_1__26__26_, connection_1__26__25_, connection_1__26__24_,
         connection_1__26__23_, connection_1__26__22_, connection_1__26__21_,
         connection_1__26__20_, connection_1__26__19_, connection_1__26__18_,
         connection_1__26__17_, connection_1__26__16_, connection_1__26__15_,
         connection_1__26__14_, connection_1__26__13_, connection_1__26__12_,
         connection_1__26__11_, connection_1__26__10_, connection_1__26__9_,
         connection_1__26__8_, connection_1__26__7_, connection_1__26__6_,
         connection_1__26__5_, connection_1__26__4_, connection_1__26__3_,
         connection_1__26__2_, connection_1__26__1_, connection_1__26__0_,
         connection_1__27__31_, connection_1__27__30_, connection_1__27__29_,
         connection_1__27__28_, connection_1__27__27_, connection_1__27__26_,
         connection_1__27__25_, connection_1__27__24_, connection_1__27__23_,
         connection_1__27__22_, connection_1__27__21_, connection_1__27__20_,
         connection_1__27__19_, connection_1__27__18_, connection_1__27__17_,
         connection_1__27__16_, connection_1__27__15_, connection_1__27__14_,
         connection_1__27__13_, connection_1__27__12_, connection_1__27__11_,
         connection_1__27__10_, connection_1__27__9_, connection_1__27__8_,
         connection_1__27__7_, connection_1__27__6_, connection_1__27__5_,
         connection_1__27__4_, connection_1__27__3_, connection_1__27__2_,
         connection_1__27__1_, connection_1__27__0_, connection_1__28__31_,
         connection_1__28__30_, connection_1__28__29_, connection_1__28__28_,
         connection_1__28__27_, connection_1__28__26_, connection_1__28__25_,
         connection_1__28__24_, connection_1__28__23_, connection_1__28__22_,
         connection_1__28__21_, connection_1__28__20_, connection_1__28__19_,
         connection_1__28__18_, connection_1__28__17_, connection_1__28__16_,
         connection_1__28__15_, connection_1__28__14_, connection_1__28__13_,
         connection_1__28__12_, connection_1__28__11_, connection_1__28__10_,
         connection_1__28__9_, connection_1__28__8_, connection_1__28__7_,
         connection_1__28__6_, connection_1__28__5_, connection_1__28__4_,
         connection_1__28__3_, connection_1__28__2_, connection_1__28__1_,
         connection_1__28__0_, connection_1__29__31_, connection_1__29__30_,
         connection_1__29__29_, connection_1__29__28_, connection_1__29__27_,
         connection_1__29__26_, connection_1__29__25_, connection_1__29__24_,
         connection_1__29__23_, connection_1__29__22_, connection_1__29__21_,
         connection_1__29__20_, connection_1__29__19_, connection_1__29__18_,
         connection_1__29__17_, connection_1__29__16_, connection_1__29__15_,
         connection_1__29__14_, connection_1__29__13_, connection_1__29__12_,
         connection_1__29__11_, connection_1__29__10_, connection_1__29__9_,
         connection_1__29__8_, connection_1__29__7_, connection_1__29__6_,
         connection_1__29__5_, connection_1__29__4_, connection_1__29__3_,
         connection_1__29__2_, connection_1__29__1_, connection_1__29__0_,
         connection_1__30__31_, connection_1__30__30_, connection_1__30__29_,
         connection_1__30__28_, connection_1__30__27_, connection_1__30__26_,
         connection_1__30__25_, connection_1__30__24_, connection_1__30__23_,
         connection_1__30__22_, connection_1__30__21_, connection_1__30__20_,
         connection_1__30__19_, connection_1__30__18_, connection_1__30__17_,
         connection_1__30__16_, connection_1__30__15_, connection_1__30__14_,
         connection_1__30__13_, connection_1__30__12_, connection_1__30__11_,
         connection_1__30__10_, connection_1__30__9_, connection_1__30__8_,
         connection_1__30__7_, connection_1__30__6_, connection_1__30__5_,
         connection_1__30__4_, connection_1__30__3_, connection_1__30__2_,
         connection_1__30__1_, connection_1__30__0_, connection_1__31__31_,
         connection_1__31__30_, connection_1__31__29_, connection_1__31__28_,
         connection_1__31__27_, connection_1__31__26_, connection_1__31__25_,
         connection_1__31__24_, connection_1__31__23_, connection_1__31__22_,
         connection_1__31__21_, connection_1__31__20_, connection_1__31__19_,
         connection_1__31__18_, connection_1__31__17_, connection_1__31__16_,
         connection_1__31__15_, connection_1__31__14_, connection_1__31__13_,
         connection_1__31__12_, connection_1__31__11_, connection_1__31__10_,
         connection_1__31__9_, connection_1__31__8_, connection_1__31__7_,
         connection_1__31__6_, connection_1__31__5_, connection_1__31__4_,
         connection_1__31__3_, connection_1__31__2_, connection_1__31__1_,
         connection_1__31__0_, connection_2__0__31_, connection_2__0__30_,
         connection_2__0__29_, connection_2__0__28_, connection_2__0__27_,
         connection_2__0__26_, connection_2__0__25_, connection_2__0__24_,
         connection_2__0__23_, connection_2__0__22_, connection_2__0__21_,
         connection_2__0__20_, connection_2__0__19_, connection_2__0__18_,
         connection_2__0__17_, connection_2__0__16_, connection_2__0__15_,
         connection_2__0__14_, connection_2__0__13_, connection_2__0__12_,
         connection_2__0__11_, connection_2__0__10_, connection_2__0__9_,
         connection_2__0__8_, connection_2__0__7_, connection_2__0__6_,
         connection_2__0__5_, connection_2__0__4_, connection_2__0__3_,
         connection_2__0__2_, connection_2__0__1_, connection_2__0__0_,
         connection_2__1__31_, connection_2__1__30_, connection_2__1__29_,
         connection_2__1__28_, connection_2__1__27_, connection_2__1__26_,
         connection_2__1__25_, connection_2__1__24_, connection_2__1__23_,
         connection_2__1__22_, connection_2__1__21_, connection_2__1__20_,
         connection_2__1__19_, connection_2__1__18_, connection_2__1__17_,
         connection_2__1__16_, connection_2__1__15_, connection_2__1__14_,
         connection_2__1__13_, connection_2__1__12_, connection_2__1__11_,
         connection_2__1__10_, connection_2__1__9_, connection_2__1__8_,
         connection_2__1__7_, connection_2__1__6_, connection_2__1__5_,
         connection_2__1__4_, connection_2__1__3_, connection_2__1__2_,
         connection_2__1__1_, connection_2__1__0_, connection_2__2__31_,
         connection_2__2__30_, connection_2__2__29_, connection_2__2__28_,
         connection_2__2__27_, connection_2__2__26_, connection_2__2__25_,
         connection_2__2__24_, connection_2__2__23_, connection_2__2__22_,
         connection_2__2__21_, connection_2__2__20_, connection_2__2__19_,
         connection_2__2__18_, connection_2__2__17_, connection_2__2__16_,
         connection_2__2__15_, connection_2__2__14_, connection_2__2__13_,
         connection_2__2__12_, connection_2__2__11_, connection_2__2__10_,
         connection_2__2__9_, connection_2__2__8_, connection_2__2__7_,
         connection_2__2__6_, connection_2__2__5_, connection_2__2__4_,
         connection_2__2__3_, connection_2__2__2_, connection_2__2__1_,
         connection_2__2__0_, connection_2__3__31_, connection_2__3__30_,
         connection_2__3__29_, connection_2__3__28_, connection_2__3__27_,
         connection_2__3__26_, connection_2__3__25_, connection_2__3__24_,
         connection_2__3__23_, connection_2__3__22_, connection_2__3__21_,
         connection_2__3__20_, connection_2__3__19_, connection_2__3__18_,
         connection_2__3__17_, connection_2__3__16_, connection_2__3__15_,
         connection_2__3__14_, connection_2__3__13_, connection_2__3__12_,
         connection_2__3__11_, connection_2__3__10_, connection_2__3__9_,
         connection_2__3__8_, connection_2__3__7_, connection_2__3__6_,
         connection_2__3__5_, connection_2__3__4_, connection_2__3__3_,
         connection_2__3__2_, connection_2__3__1_, connection_2__3__0_,
         connection_2__4__31_, connection_2__4__30_, connection_2__4__29_,
         connection_2__4__28_, connection_2__4__27_, connection_2__4__26_,
         connection_2__4__25_, connection_2__4__24_, connection_2__4__23_,
         connection_2__4__22_, connection_2__4__21_, connection_2__4__20_,
         connection_2__4__19_, connection_2__4__18_, connection_2__4__17_,
         connection_2__4__16_, connection_2__4__15_, connection_2__4__14_,
         connection_2__4__13_, connection_2__4__12_, connection_2__4__11_,
         connection_2__4__10_, connection_2__4__9_, connection_2__4__8_,
         connection_2__4__7_, connection_2__4__6_, connection_2__4__5_,
         connection_2__4__4_, connection_2__4__3_, connection_2__4__2_,
         connection_2__4__1_, connection_2__4__0_, connection_2__5__31_,
         connection_2__5__30_, connection_2__5__29_, connection_2__5__28_,
         connection_2__5__27_, connection_2__5__26_, connection_2__5__25_,
         connection_2__5__24_, connection_2__5__23_, connection_2__5__22_,
         connection_2__5__21_, connection_2__5__20_, connection_2__5__19_,
         connection_2__5__18_, connection_2__5__17_, connection_2__5__16_,
         connection_2__5__15_, connection_2__5__14_, connection_2__5__13_,
         connection_2__5__12_, connection_2__5__11_, connection_2__5__10_,
         connection_2__5__9_, connection_2__5__8_, connection_2__5__7_,
         connection_2__5__6_, connection_2__5__5_, connection_2__5__4_,
         connection_2__5__3_, connection_2__5__2_, connection_2__5__1_,
         connection_2__5__0_, connection_2__6__31_, connection_2__6__30_,
         connection_2__6__29_, connection_2__6__28_, connection_2__6__27_,
         connection_2__6__26_, connection_2__6__25_, connection_2__6__24_,
         connection_2__6__23_, connection_2__6__22_, connection_2__6__21_,
         connection_2__6__20_, connection_2__6__19_, connection_2__6__18_,
         connection_2__6__17_, connection_2__6__16_, connection_2__6__15_,
         connection_2__6__14_, connection_2__6__13_, connection_2__6__12_,
         connection_2__6__11_, connection_2__6__10_, connection_2__6__9_,
         connection_2__6__8_, connection_2__6__7_, connection_2__6__6_,
         connection_2__6__5_, connection_2__6__4_, connection_2__6__3_,
         connection_2__6__2_, connection_2__6__1_, connection_2__6__0_,
         connection_2__7__31_, connection_2__7__30_, connection_2__7__29_,
         connection_2__7__28_, connection_2__7__27_, connection_2__7__26_,
         connection_2__7__25_, connection_2__7__24_, connection_2__7__23_,
         connection_2__7__22_, connection_2__7__21_, connection_2__7__20_,
         connection_2__7__19_, connection_2__7__18_, connection_2__7__17_,
         connection_2__7__16_, connection_2__7__15_, connection_2__7__14_,
         connection_2__7__13_, connection_2__7__12_, connection_2__7__11_,
         connection_2__7__10_, connection_2__7__9_, connection_2__7__8_,
         connection_2__7__7_, connection_2__7__6_, connection_2__7__5_,
         connection_2__7__4_, connection_2__7__3_, connection_2__7__2_,
         connection_2__7__1_, connection_2__7__0_, connection_2__8__31_,
         connection_2__8__30_, connection_2__8__29_, connection_2__8__28_,
         connection_2__8__27_, connection_2__8__26_, connection_2__8__25_,
         connection_2__8__24_, connection_2__8__23_, connection_2__8__22_,
         connection_2__8__21_, connection_2__8__20_, connection_2__8__19_,
         connection_2__8__18_, connection_2__8__17_, connection_2__8__16_,
         connection_2__8__15_, connection_2__8__14_, connection_2__8__13_,
         connection_2__8__12_, connection_2__8__11_, connection_2__8__10_,
         connection_2__8__9_, connection_2__8__8_, connection_2__8__7_,
         connection_2__8__6_, connection_2__8__5_, connection_2__8__4_,
         connection_2__8__3_, connection_2__8__2_, connection_2__8__1_,
         connection_2__8__0_, connection_2__9__31_, connection_2__9__30_,
         connection_2__9__29_, connection_2__9__28_, connection_2__9__27_,
         connection_2__9__26_, connection_2__9__25_, connection_2__9__24_,
         connection_2__9__23_, connection_2__9__22_, connection_2__9__21_,
         connection_2__9__20_, connection_2__9__19_, connection_2__9__18_,
         connection_2__9__17_, connection_2__9__16_, connection_2__9__15_,
         connection_2__9__14_, connection_2__9__13_, connection_2__9__12_,
         connection_2__9__11_, connection_2__9__10_, connection_2__9__9_,
         connection_2__9__8_, connection_2__9__7_, connection_2__9__6_,
         connection_2__9__5_, connection_2__9__4_, connection_2__9__3_,
         connection_2__9__2_, connection_2__9__1_, connection_2__9__0_,
         connection_2__10__31_, connection_2__10__30_, connection_2__10__29_,
         connection_2__10__28_, connection_2__10__27_, connection_2__10__26_,
         connection_2__10__25_, connection_2__10__24_, connection_2__10__23_,
         connection_2__10__22_, connection_2__10__21_, connection_2__10__20_,
         connection_2__10__19_, connection_2__10__18_, connection_2__10__17_,
         connection_2__10__16_, connection_2__10__15_, connection_2__10__14_,
         connection_2__10__13_, connection_2__10__12_, connection_2__10__11_,
         connection_2__10__10_, connection_2__10__9_, connection_2__10__8_,
         connection_2__10__7_, connection_2__10__6_, connection_2__10__5_,
         connection_2__10__4_, connection_2__10__3_, connection_2__10__2_,
         connection_2__10__1_, connection_2__10__0_, connection_2__11__31_,
         connection_2__11__30_, connection_2__11__29_, connection_2__11__28_,
         connection_2__11__27_, connection_2__11__26_, connection_2__11__25_,
         connection_2__11__24_, connection_2__11__23_, connection_2__11__22_,
         connection_2__11__21_, connection_2__11__20_, connection_2__11__19_,
         connection_2__11__18_, connection_2__11__17_, connection_2__11__16_,
         connection_2__11__15_, connection_2__11__14_, connection_2__11__13_,
         connection_2__11__12_, connection_2__11__11_, connection_2__11__10_,
         connection_2__11__9_, connection_2__11__8_, connection_2__11__7_,
         connection_2__11__6_, connection_2__11__5_, connection_2__11__4_,
         connection_2__11__3_, connection_2__11__2_, connection_2__11__1_,
         connection_2__11__0_, connection_2__12__31_, connection_2__12__30_,
         connection_2__12__29_, connection_2__12__28_, connection_2__12__27_,
         connection_2__12__26_, connection_2__12__25_, connection_2__12__24_,
         connection_2__12__23_, connection_2__12__22_, connection_2__12__21_,
         connection_2__12__20_, connection_2__12__19_, connection_2__12__18_,
         connection_2__12__17_, connection_2__12__16_, connection_2__12__15_,
         connection_2__12__14_, connection_2__12__13_, connection_2__12__12_,
         connection_2__12__11_, connection_2__12__10_, connection_2__12__9_,
         connection_2__12__8_, connection_2__12__7_, connection_2__12__6_,
         connection_2__12__5_, connection_2__12__4_, connection_2__12__3_,
         connection_2__12__2_, connection_2__12__1_, connection_2__12__0_,
         connection_2__13__31_, connection_2__13__30_, connection_2__13__29_,
         connection_2__13__28_, connection_2__13__27_, connection_2__13__26_,
         connection_2__13__25_, connection_2__13__24_, connection_2__13__23_,
         connection_2__13__22_, connection_2__13__21_, connection_2__13__20_,
         connection_2__13__19_, connection_2__13__18_, connection_2__13__17_,
         connection_2__13__16_, connection_2__13__15_, connection_2__13__14_,
         connection_2__13__13_, connection_2__13__12_, connection_2__13__11_,
         connection_2__13__10_, connection_2__13__9_, connection_2__13__8_,
         connection_2__13__7_, connection_2__13__6_, connection_2__13__5_,
         connection_2__13__4_, connection_2__13__3_, connection_2__13__2_,
         connection_2__13__1_, connection_2__13__0_, connection_2__14__31_,
         connection_2__14__30_, connection_2__14__29_, connection_2__14__28_,
         connection_2__14__27_, connection_2__14__26_, connection_2__14__25_,
         connection_2__14__24_, connection_2__14__23_, connection_2__14__22_,
         connection_2__14__21_, connection_2__14__20_, connection_2__14__19_,
         connection_2__14__18_, connection_2__14__17_, connection_2__14__16_,
         connection_2__14__15_, connection_2__14__14_, connection_2__14__13_,
         connection_2__14__12_, connection_2__14__11_, connection_2__14__10_,
         connection_2__14__9_, connection_2__14__8_, connection_2__14__7_,
         connection_2__14__6_, connection_2__14__5_, connection_2__14__4_,
         connection_2__14__3_, connection_2__14__2_, connection_2__14__1_,
         connection_2__14__0_, connection_2__15__31_, connection_2__15__30_,
         connection_2__15__29_, connection_2__15__28_, connection_2__15__27_,
         connection_2__15__26_, connection_2__15__25_, connection_2__15__24_,
         connection_2__15__23_, connection_2__15__22_, connection_2__15__21_,
         connection_2__15__20_, connection_2__15__19_, connection_2__15__18_,
         connection_2__15__17_, connection_2__15__16_, connection_2__15__15_,
         connection_2__15__14_, connection_2__15__13_, connection_2__15__12_,
         connection_2__15__11_, connection_2__15__10_, connection_2__15__9_,
         connection_2__15__8_, connection_2__15__7_, connection_2__15__6_,
         connection_2__15__5_, connection_2__15__4_, connection_2__15__3_,
         connection_2__15__2_, connection_2__15__1_, connection_2__15__0_,
         connection_2__16__31_, connection_2__16__30_, connection_2__16__29_,
         connection_2__16__28_, connection_2__16__27_, connection_2__16__26_,
         connection_2__16__25_, connection_2__16__24_, connection_2__16__23_,
         connection_2__16__22_, connection_2__16__21_, connection_2__16__20_,
         connection_2__16__19_, connection_2__16__18_, connection_2__16__17_,
         connection_2__16__16_, connection_2__16__15_, connection_2__16__14_,
         connection_2__16__13_, connection_2__16__12_, connection_2__16__11_,
         connection_2__16__10_, connection_2__16__9_, connection_2__16__8_,
         connection_2__16__7_, connection_2__16__6_, connection_2__16__5_,
         connection_2__16__4_, connection_2__16__3_, connection_2__16__2_,
         connection_2__16__1_, connection_2__16__0_, connection_2__17__31_,
         connection_2__17__30_, connection_2__17__29_, connection_2__17__28_,
         connection_2__17__27_, connection_2__17__26_, connection_2__17__25_,
         connection_2__17__24_, connection_2__17__23_, connection_2__17__22_,
         connection_2__17__21_, connection_2__17__20_, connection_2__17__19_,
         connection_2__17__18_, connection_2__17__17_, connection_2__17__16_,
         connection_2__17__15_, connection_2__17__14_, connection_2__17__13_,
         connection_2__17__12_, connection_2__17__11_, connection_2__17__10_,
         connection_2__17__9_, connection_2__17__8_, connection_2__17__7_,
         connection_2__17__6_, connection_2__17__5_, connection_2__17__4_,
         connection_2__17__3_, connection_2__17__2_, connection_2__17__1_,
         connection_2__17__0_, connection_2__18__31_, connection_2__18__30_,
         connection_2__18__29_, connection_2__18__28_, connection_2__18__27_,
         connection_2__18__26_, connection_2__18__25_, connection_2__18__24_,
         connection_2__18__23_, connection_2__18__22_, connection_2__18__21_,
         connection_2__18__20_, connection_2__18__19_, connection_2__18__18_,
         connection_2__18__17_, connection_2__18__16_, connection_2__18__15_,
         connection_2__18__14_, connection_2__18__13_, connection_2__18__12_,
         connection_2__18__11_, connection_2__18__10_, connection_2__18__9_,
         connection_2__18__8_, connection_2__18__7_, connection_2__18__6_,
         connection_2__18__5_, connection_2__18__4_, connection_2__18__3_,
         connection_2__18__2_, connection_2__18__1_, connection_2__18__0_,
         connection_2__19__31_, connection_2__19__30_, connection_2__19__29_,
         connection_2__19__28_, connection_2__19__27_, connection_2__19__26_,
         connection_2__19__25_, connection_2__19__24_, connection_2__19__23_,
         connection_2__19__22_, connection_2__19__21_, connection_2__19__20_,
         connection_2__19__19_, connection_2__19__18_, connection_2__19__17_,
         connection_2__19__16_, connection_2__19__15_, connection_2__19__14_,
         connection_2__19__13_, connection_2__19__12_, connection_2__19__11_,
         connection_2__19__10_, connection_2__19__9_, connection_2__19__8_,
         connection_2__19__7_, connection_2__19__6_, connection_2__19__5_,
         connection_2__19__4_, connection_2__19__3_, connection_2__19__2_,
         connection_2__19__1_, connection_2__19__0_, connection_2__20__31_,
         connection_2__20__30_, connection_2__20__29_, connection_2__20__28_,
         connection_2__20__27_, connection_2__20__26_, connection_2__20__25_,
         connection_2__20__24_, connection_2__20__23_, connection_2__20__22_,
         connection_2__20__21_, connection_2__20__20_, connection_2__20__19_,
         connection_2__20__18_, connection_2__20__17_, connection_2__20__16_,
         connection_2__20__15_, connection_2__20__14_, connection_2__20__13_,
         connection_2__20__12_, connection_2__20__11_, connection_2__20__10_,
         connection_2__20__9_, connection_2__20__8_, connection_2__20__7_,
         connection_2__20__6_, connection_2__20__5_, connection_2__20__4_,
         connection_2__20__3_, connection_2__20__2_, connection_2__20__1_,
         connection_2__20__0_, connection_2__21__31_, connection_2__21__30_,
         connection_2__21__29_, connection_2__21__28_, connection_2__21__27_,
         connection_2__21__26_, connection_2__21__25_, connection_2__21__24_,
         connection_2__21__23_, connection_2__21__22_, connection_2__21__21_,
         connection_2__21__20_, connection_2__21__19_, connection_2__21__18_,
         connection_2__21__17_, connection_2__21__16_, connection_2__21__15_,
         connection_2__21__14_, connection_2__21__13_, connection_2__21__12_,
         connection_2__21__11_, connection_2__21__10_, connection_2__21__9_,
         connection_2__21__8_, connection_2__21__7_, connection_2__21__6_,
         connection_2__21__5_, connection_2__21__4_, connection_2__21__3_,
         connection_2__21__2_, connection_2__21__1_, connection_2__21__0_,
         connection_2__22__31_, connection_2__22__30_, connection_2__22__29_,
         connection_2__22__28_, connection_2__22__27_, connection_2__22__26_,
         connection_2__22__25_, connection_2__22__24_, connection_2__22__23_,
         connection_2__22__22_, connection_2__22__21_, connection_2__22__20_,
         connection_2__22__19_, connection_2__22__18_, connection_2__22__17_,
         connection_2__22__16_, connection_2__22__15_, connection_2__22__14_,
         connection_2__22__13_, connection_2__22__12_, connection_2__22__11_,
         connection_2__22__10_, connection_2__22__9_, connection_2__22__8_,
         connection_2__22__7_, connection_2__22__6_, connection_2__22__5_,
         connection_2__22__4_, connection_2__22__3_, connection_2__22__2_,
         connection_2__22__1_, connection_2__22__0_, connection_2__23__31_,
         connection_2__23__30_, connection_2__23__29_, connection_2__23__28_,
         connection_2__23__27_, connection_2__23__26_, connection_2__23__25_,
         connection_2__23__24_, connection_2__23__23_, connection_2__23__22_,
         connection_2__23__21_, connection_2__23__20_, connection_2__23__19_,
         connection_2__23__18_, connection_2__23__17_, connection_2__23__16_,
         connection_2__23__15_, connection_2__23__14_, connection_2__23__13_,
         connection_2__23__12_, connection_2__23__11_, connection_2__23__10_,
         connection_2__23__9_, connection_2__23__8_, connection_2__23__7_,
         connection_2__23__6_, connection_2__23__5_, connection_2__23__4_,
         connection_2__23__3_, connection_2__23__2_, connection_2__23__1_,
         connection_2__23__0_, connection_2__24__31_, connection_2__24__30_,
         connection_2__24__29_, connection_2__24__28_, connection_2__24__27_,
         connection_2__24__26_, connection_2__24__25_, connection_2__24__24_,
         connection_2__24__23_, connection_2__24__22_, connection_2__24__21_,
         connection_2__24__20_, connection_2__24__19_, connection_2__24__18_,
         connection_2__24__17_, connection_2__24__16_, connection_2__24__15_,
         connection_2__24__14_, connection_2__24__13_, connection_2__24__12_,
         connection_2__24__11_, connection_2__24__10_, connection_2__24__9_,
         connection_2__24__8_, connection_2__24__7_, connection_2__24__6_,
         connection_2__24__5_, connection_2__24__4_, connection_2__24__3_,
         connection_2__24__2_, connection_2__24__1_, connection_2__24__0_,
         connection_2__25__31_, connection_2__25__30_, connection_2__25__29_,
         connection_2__25__28_, connection_2__25__27_, connection_2__25__26_,
         connection_2__25__25_, connection_2__25__24_, connection_2__25__23_,
         connection_2__25__22_, connection_2__25__21_, connection_2__25__20_,
         connection_2__25__19_, connection_2__25__18_, connection_2__25__17_,
         connection_2__25__16_, connection_2__25__15_, connection_2__25__14_,
         connection_2__25__13_, connection_2__25__12_, connection_2__25__11_,
         connection_2__25__10_, connection_2__25__9_, connection_2__25__8_,
         connection_2__25__7_, connection_2__25__6_, connection_2__25__5_,
         connection_2__25__4_, connection_2__25__3_, connection_2__25__2_,
         connection_2__25__1_, connection_2__25__0_, connection_2__26__31_,
         connection_2__26__30_, connection_2__26__29_, connection_2__26__28_,
         connection_2__26__27_, connection_2__26__26_, connection_2__26__25_,
         connection_2__26__24_, connection_2__26__23_, connection_2__26__22_,
         connection_2__26__21_, connection_2__26__20_, connection_2__26__19_,
         connection_2__26__18_, connection_2__26__17_, connection_2__26__16_,
         connection_2__26__15_, connection_2__26__14_, connection_2__26__13_,
         connection_2__26__12_, connection_2__26__11_, connection_2__26__10_,
         connection_2__26__9_, connection_2__26__8_, connection_2__26__7_,
         connection_2__26__6_, connection_2__26__5_, connection_2__26__4_,
         connection_2__26__3_, connection_2__26__2_, connection_2__26__1_,
         connection_2__26__0_, connection_2__27__31_, connection_2__27__30_,
         connection_2__27__29_, connection_2__27__28_, connection_2__27__27_,
         connection_2__27__26_, connection_2__27__25_, connection_2__27__24_,
         connection_2__27__23_, connection_2__27__22_, connection_2__27__21_,
         connection_2__27__20_, connection_2__27__19_, connection_2__27__18_,
         connection_2__27__17_, connection_2__27__16_, connection_2__27__15_,
         connection_2__27__14_, connection_2__27__13_, connection_2__27__12_,
         connection_2__27__11_, connection_2__27__10_, connection_2__27__9_,
         connection_2__27__8_, connection_2__27__7_, connection_2__27__6_,
         connection_2__27__5_, connection_2__27__4_, connection_2__27__3_,
         connection_2__27__2_, connection_2__27__1_, connection_2__27__0_,
         connection_2__28__31_, connection_2__28__30_, connection_2__28__29_,
         connection_2__28__28_, connection_2__28__27_, connection_2__28__26_,
         connection_2__28__25_, connection_2__28__24_, connection_2__28__23_,
         connection_2__28__22_, connection_2__28__21_, connection_2__28__20_,
         connection_2__28__19_, connection_2__28__18_, connection_2__28__17_,
         connection_2__28__16_, connection_2__28__15_, connection_2__28__14_,
         connection_2__28__13_, connection_2__28__12_, connection_2__28__11_,
         connection_2__28__10_, connection_2__28__9_, connection_2__28__8_,
         connection_2__28__7_, connection_2__28__6_, connection_2__28__5_,
         connection_2__28__4_, connection_2__28__3_, connection_2__28__2_,
         connection_2__28__1_, connection_2__28__0_, connection_2__29__31_,
         connection_2__29__30_, connection_2__29__29_, connection_2__29__28_,
         connection_2__29__27_, connection_2__29__26_, connection_2__29__25_,
         connection_2__29__24_, connection_2__29__23_, connection_2__29__22_,
         connection_2__29__21_, connection_2__29__20_, connection_2__29__19_,
         connection_2__29__18_, connection_2__29__17_, connection_2__29__16_,
         connection_2__29__15_, connection_2__29__14_, connection_2__29__13_,
         connection_2__29__12_, connection_2__29__11_, connection_2__29__10_,
         connection_2__29__9_, connection_2__29__8_, connection_2__29__7_,
         connection_2__29__6_, connection_2__29__5_, connection_2__29__4_,
         connection_2__29__3_, connection_2__29__2_, connection_2__29__1_,
         connection_2__29__0_, connection_2__30__31_, connection_2__30__30_,
         connection_2__30__29_, connection_2__30__28_, connection_2__30__27_,
         connection_2__30__26_, connection_2__30__25_, connection_2__30__24_,
         connection_2__30__23_, connection_2__30__22_, connection_2__30__21_,
         connection_2__30__20_, connection_2__30__19_, connection_2__30__18_,
         connection_2__30__17_, connection_2__30__16_, connection_2__30__15_,
         connection_2__30__14_, connection_2__30__13_, connection_2__30__12_,
         connection_2__30__11_, connection_2__30__10_, connection_2__30__9_,
         connection_2__30__8_, connection_2__30__7_, connection_2__30__6_,
         connection_2__30__5_, connection_2__30__4_, connection_2__30__3_,
         connection_2__30__2_, connection_2__30__1_, connection_2__30__0_,
         connection_2__31__31_, connection_2__31__30_, connection_2__31__29_,
         connection_2__31__28_, connection_2__31__27_, connection_2__31__26_,
         connection_2__31__25_, connection_2__31__24_, connection_2__31__23_,
         connection_2__31__22_, connection_2__31__21_, connection_2__31__20_,
         connection_2__31__19_, connection_2__31__18_, connection_2__31__17_,
         connection_2__31__16_, connection_2__31__15_, connection_2__31__14_,
         connection_2__31__13_, connection_2__31__12_, connection_2__31__11_,
         connection_2__31__10_, connection_2__31__9_, connection_2__31__8_,
         connection_2__31__7_, connection_2__31__6_, connection_2__31__5_,
         connection_2__31__4_, connection_2__31__3_, connection_2__31__2_,
         connection_2__31__1_, connection_2__31__0_, connection_3__0__31_,
         connection_3__0__30_, connection_3__0__29_, connection_3__0__28_,
         connection_3__0__27_, connection_3__0__26_, connection_3__0__25_,
         connection_3__0__24_, connection_3__0__23_, connection_3__0__22_,
         connection_3__0__21_, connection_3__0__20_, connection_3__0__19_,
         connection_3__0__18_, connection_3__0__17_, connection_3__0__16_,
         connection_3__0__15_, connection_3__0__14_, connection_3__0__13_,
         connection_3__0__12_, connection_3__0__11_, connection_3__0__10_,
         connection_3__0__9_, connection_3__0__8_, connection_3__0__7_,
         connection_3__0__6_, connection_3__0__5_, connection_3__0__4_,
         connection_3__0__3_, connection_3__0__2_, connection_3__0__1_,
         connection_3__0__0_, connection_3__1__31_, connection_3__1__30_,
         connection_3__1__29_, connection_3__1__28_, connection_3__1__27_,
         connection_3__1__26_, connection_3__1__25_, connection_3__1__24_,
         connection_3__1__23_, connection_3__1__22_, connection_3__1__21_,
         connection_3__1__20_, connection_3__1__19_, connection_3__1__18_,
         connection_3__1__17_, connection_3__1__16_, connection_3__1__15_,
         connection_3__1__14_, connection_3__1__13_, connection_3__1__12_,
         connection_3__1__11_, connection_3__1__10_, connection_3__1__9_,
         connection_3__1__8_, connection_3__1__7_, connection_3__1__6_,
         connection_3__1__5_, connection_3__1__4_, connection_3__1__3_,
         connection_3__1__2_, connection_3__1__1_, connection_3__1__0_,
         connection_3__2__31_, connection_3__2__30_, connection_3__2__29_,
         connection_3__2__28_, connection_3__2__27_, connection_3__2__26_,
         connection_3__2__25_, connection_3__2__24_, connection_3__2__23_,
         connection_3__2__22_, connection_3__2__21_, connection_3__2__20_,
         connection_3__2__19_, connection_3__2__18_, connection_3__2__17_,
         connection_3__2__16_, connection_3__2__15_, connection_3__2__14_,
         connection_3__2__13_, connection_3__2__12_, connection_3__2__11_,
         connection_3__2__10_, connection_3__2__9_, connection_3__2__8_,
         connection_3__2__7_, connection_3__2__6_, connection_3__2__5_,
         connection_3__2__4_, connection_3__2__3_, connection_3__2__2_,
         connection_3__2__1_, connection_3__2__0_, connection_3__3__31_,
         connection_3__3__30_, connection_3__3__29_, connection_3__3__28_,
         connection_3__3__27_, connection_3__3__26_, connection_3__3__25_,
         connection_3__3__24_, connection_3__3__23_, connection_3__3__22_,
         connection_3__3__21_, connection_3__3__20_, connection_3__3__19_,
         connection_3__3__18_, connection_3__3__17_, connection_3__3__16_,
         connection_3__3__15_, connection_3__3__14_, connection_3__3__13_,
         connection_3__3__12_, connection_3__3__11_, connection_3__3__10_,
         connection_3__3__9_, connection_3__3__8_, connection_3__3__7_,
         connection_3__3__6_, connection_3__3__5_, connection_3__3__4_,
         connection_3__3__3_, connection_3__3__2_, connection_3__3__1_,
         connection_3__3__0_, connection_3__4__31_, connection_3__4__30_,
         connection_3__4__29_, connection_3__4__28_, connection_3__4__27_,
         connection_3__4__26_, connection_3__4__25_, connection_3__4__24_,
         connection_3__4__23_, connection_3__4__22_, connection_3__4__21_,
         connection_3__4__20_, connection_3__4__19_, connection_3__4__18_,
         connection_3__4__17_, connection_3__4__16_, connection_3__4__15_,
         connection_3__4__14_, connection_3__4__13_, connection_3__4__12_,
         connection_3__4__11_, connection_3__4__10_, connection_3__4__9_,
         connection_3__4__8_, connection_3__4__7_, connection_3__4__6_,
         connection_3__4__5_, connection_3__4__4_, connection_3__4__3_,
         connection_3__4__2_, connection_3__4__1_, connection_3__4__0_,
         connection_3__5__31_, connection_3__5__30_, connection_3__5__29_,
         connection_3__5__28_, connection_3__5__27_, connection_3__5__26_,
         connection_3__5__25_, connection_3__5__24_, connection_3__5__23_,
         connection_3__5__22_, connection_3__5__21_, connection_3__5__20_,
         connection_3__5__19_, connection_3__5__18_, connection_3__5__17_,
         connection_3__5__16_, connection_3__5__15_, connection_3__5__14_,
         connection_3__5__13_, connection_3__5__12_, connection_3__5__11_,
         connection_3__5__10_, connection_3__5__9_, connection_3__5__8_,
         connection_3__5__7_, connection_3__5__6_, connection_3__5__5_,
         connection_3__5__4_, connection_3__5__3_, connection_3__5__2_,
         connection_3__5__1_, connection_3__5__0_, connection_3__6__31_,
         connection_3__6__30_, connection_3__6__29_, connection_3__6__28_,
         connection_3__6__27_, connection_3__6__26_, connection_3__6__25_,
         connection_3__6__24_, connection_3__6__23_, connection_3__6__22_,
         connection_3__6__21_, connection_3__6__20_, connection_3__6__19_,
         connection_3__6__18_, connection_3__6__17_, connection_3__6__16_,
         connection_3__6__15_, connection_3__6__14_, connection_3__6__13_,
         connection_3__6__12_, connection_3__6__11_, connection_3__6__10_,
         connection_3__6__9_, connection_3__6__8_, connection_3__6__7_,
         connection_3__6__6_, connection_3__6__5_, connection_3__6__4_,
         connection_3__6__3_, connection_3__6__2_, connection_3__6__1_,
         connection_3__6__0_, connection_3__7__31_, connection_3__7__30_,
         connection_3__7__29_, connection_3__7__28_, connection_3__7__27_,
         connection_3__7__26_, connection_3__7__25_, connection_3__7__24_,
         connection_3__7__23_, connection_3__7__22_, connection_3__7__21_,
         connection_3__7__20_, connection_3__7__19_, connection_3__7__18_,
         connection_3__7__17_, connection_3__7__16_, connection_3__7__15_,
         connection_3__7__14_, connection_3__7__13_, connection_3__7__12_,
         connection_3__7__11_, connection_3__7__10_, connection_3__7__9_,
         connection_3__7__8_, connection_3__7__7_, connection_3__7__6_,
         connection_3__7__5_, connection_3__7__4_, connection_3__7__3_,
         connection_3__7__2_, connection_3__7__1_, connection_3__7__0_,
         connection_3__8__31_, connection_3__8__30_, connection_3__8__29_,
         connection_3__8__28_, connection_3__8__27_, connection_3__8__26_,
         connection_3__8__25_, connection_3__8__24_, connection_3__8__23_,
         connection_3__8__22_, connection_3__8__21_, connection_3__8__20_,
         connection_3__8__19_, connection_3__8__18_, connection_3__8__17_,
         connection_3__8__16_, connection_3__8__15_, connection_3__8__14_,
         connection_3__8__13_, connection_3__8__12_, connection_3__8__11_,
         connection_3__8__10_, connection_3__8__9_, connection_3__8__8_,
         connection_3__8__7_, connection_3__8__6_, connection_3__8__5_,
         connection_3__8__4_, connection_3__8__3_, connection_3__8__2_,
         connection_3__8__1_, connection_3__8__0_, connection_3__9__31_,
         connection_3__9__30_, connection_3__9__29_, connection_3__9__28_,
         connection_3__9__27_, connection_3__9__26_, connection_3__9__25_,
         connection_3__9__24_, connection_3__9__23_, connection_3__9__22_,
         connection_3__9__21_, connection_3__9__20_, connection_3__9__19_,
         connection_3__9__18_, connection_3__9__17_, connection_3__9__16_,
         connection_3__9__15_, connection_3__9__14_, connection_3__9__13_,
         connection_3__9__12_, connection_3__9__11_, connection_3__9__10_,
         connection_3__9__9_, connection_3__9__8_, connection_3__9__7_,
         connection_3__9__6_, connection_3__9__5_, connection_3__9__4_,
         connection_3__9__3_, connection_3__9__2_, connection_3__9__1_,
         connection_3__9__0_, connection_3__10__31_, connection_3__10__30_,
         connection_3__10__29_, connection_3__10__28_, connection_3__10__27_,
         connection_3__10__26_, connection_3__10__25_, connection_3__10__24_,
         connection_3__10__23_, connection_3__10__22_, connection_3__10__21_,
         connection_3__10__20_, connection_3__10__19_, connection_3__10__18_,
         connection_3__10__17_, connection_3__10__16_, connection_3__10__15_,
         connection_3__10__14_, connection_3__10__13_, connection_3__10__12_,
         connection_3__10__11_, connection_3__10__10_, connection_3__10__9_,
         connection_3__10__8_, connection_3__10__7_, connection_3__10__6_,
         connection_3__10__5_, connection_3__10__4_, connection_3__10__3_,
         connection_3__10__2_, connection_3__10__1_, connection_3__10__0_,
         connection_3__11__31_, connection_3__11__30_, connection_3__11__29_,
         connection_3__11__28_, connection_3__11__27_, connection_3__11__26_,
         connection_3__11__25_, connection_3__11__24_, connection_3__11__23_,
         connection_3__11__22_, connection_3__11__21_, connection_3__11__20_,
         connection_3__11__19_, connection_3__11__18_, connection_3__11__17_,
         connection_3__11__16_, connection_3__11__15_, connection_3__11__14_,
         connection_3__11__13_, connection_3__11__12_, connection_3__11__11_,
         connection_3__11__10_, connection_3__11__9_, connection_3__11__8_,
         connection_3__11__7_, connection_3__11__6_, connection_3__11__5_,
         connection_3__11__4_, connection_3__11__3_, connection_3__11__2_,
         connection_3__11__1_, connection_3__11__0_, connection_3__12__31_,
         connection_3__12__30_, connection_3__12__29_, connection_3__12__28_,
         connection_3__12__27_, connection_3__12__26_, connection_3__12__25_,
         connection_3__12__24_, connection_3__12__23_, connection_3__12__22_,
         connection_3__12__21_, connection_3__12__20_, connection_3__12__19_,
         connection_3__12__18_, connection_3__12__17_, connection_3__12__16_,
         connection_3__12__15_, connection_3__12__14_, connection_3__12__13_,
         connection_3__12__12_, connection_3__12__11_, connection_3__12__10_,
         connection_3__12__9_, connection_3__12__8_, connection_3__12__7_,
         connection_3__12__6_, connection_3__12__5_, connection_3__12__4_,
         connection_3__12__3_, connection_3__12__2_, connection_3__12__1_,
         connection_3__12__0_, connection_3__13__31_, connection_3__13__30_,
         connection_3__13__29_, connection_3__13__28_, connection_3__13__27_,
         connection_3__13__26_, connection_3__13__25_, connection_3__13__24_,
         connection_3__13__23_, connection_3__13__22_, connection_3__13__21_,
         connection_3__13__20_, connection_3__13__19_, connection_3__13__18_,
         connection_3__13__17_, connection_3__13__16_, connection_3__13__15_,
         connection_3__13__14_, connection_3__13__13_, connection_3__13__12_,
         connection_3__13__11_, connection_3__13__10_, connection_3__13__9_,
         connection_3__13__8_, connection_3__13__7_, connection_3__13__6_,
         connection_3__13__5_, connection_3__13__4_, connection_3__13__3_,
         connection_3__13__2_, connection_3__13__1_, connection_3__13__0_,
         connection_3__14__31_, connection_3__14__30_, connection_3__14__29_,
         connection_3__14__28_, connection_3__14__27_, connection_3__14__26_,
         connection_3__14__25_, connection_3__14__24_, connection_3__14__23_,
         connection_3__14__22_, connection_3__14__21_, connection_3__14__20_,
         connection_3__14__19_, connection_3__14__18_, connection_3__14__17_,
         connection_3__14__16_, connection_3__14__15_, connection_3__14__14_,
         connection_3__14__13_, connection_3__14__12_, connection_3__14__11_,
         connection_3__14__10_, connection_3__14__9_, connection_3__14__8_,
         connection_3__14__7_, connection_3__14__6_, connection_3__14__5_,
         connection_3__14__4_, connection_3__14__3_, connection_3__14__2_,
         connection_3__14__1_, connection_3__14__0_, connection_3__15__31_,
         connection_3__15__30_, connection_3__15__29_, connection_3__15__28_,
         connection_3__15__27_, connection_3__15__26_, connection_3__15__25_,
         connection_3__15__24_, connection_3__15__23_, connection_3__15__22_,
         connection_3__15__21_, connection_3__15__20_, connection_3__15__19_,
         connection_3__15__18_, connection_3__15__17_, connection_3__15__16_,
         connection_3__15__15_, connection_3__15__14_, connection_3__15__13_,
         connection_3__15__12_, connection_3__15__11_, connection_3__15__10_,
         connection_3__15__9_, connection_3__15__8_, connection_3__15__7_,
         connection_3__15__6_, connection_3__15__5_, connection_3__15__4_,
         connection_3__15__3_, connection_3__15__2_, connection_3__15__1_,
         connection_3__15__0_, connection_3__16__31_, connection_3__16__30_,
         connection_3__16__29_, connection_3__16__28_, connection_3__16__27_,
         connection_3__16__26_, connection_3__16__25_, connection_3__16__24_,
         connection_3__16__23_, connection_3__16__22_, connection_3__16__21_,
         connection_3__16__20_, connection_3__16__19_, connection_3__16__18_,
         connection_3__16__17_, connection_3__16__16_, connection_3__16__15_,
         connection_3__16__14_, connection_3__16__13_, connection_3__16__12_,
         connection_3__16__11_, connection_3__16__10_, connection_3__16__9_,
         connection_3__16__8_, connection_3__16__7_, connection_3__16__6_,
         connection_3__16__5_, connection_3__16__4_, connection_3__16__3_,
         connection_3__16__2_, connection_3__16__1_, connection_3__16__0_,
         connection_3__17__31_, connection_3__17__30_, connection_3__17__29_,
         connection_3__17__28_, connection_3__17__27_, connection_3__17__26_,
         connection_3__17__25_, connection_3__17__24_, connection_3__17__23_,
         connection_3__17__22_, connection_3__17__21_, connection_3__17__20_,
         connection_3__17__19_, connection_3__17__18_, connection_3__17__17_,
         connection_3__17__16_, connection_3__17__15_, connection_3__17__14_,
         connection_3__17__13_, connection_3__17__12_, connection_3__17__11_,
         connection_3__17__10_, connection_3__17__9_, connection_3__17__8_,
         connection_3__17__7_, connection_3__17__6_, connection_3__17__5_,
         connection_3__17__4_, connection_3__17__3_, connection_3__17__2_,
         connection_3__17__1_, connection_3__17__0_, connection_3__18__31_,
         connection_3__18__30_, connection_3__18__29_, connection_3__18__28_,
         connection_3__18__27_, connection_3__18__26_, connection_3__18__25_,
         connection_3__18__24_, connection_3__18__23_, connection_3__18__22_,
         connection_3__18__21_, connection_3__18__20_, connection_3__18__19_,
         connection_3__18__18_, connection_3__18__17_, connection_3__18__16_,
         connection_3__18__15_, connection_3__18__14_, connection_3__18__13_,
         connection_3__18__12_, connection_3__18__11_, connection_3__18__10_,
         connection_3__18__9_, connection_3__18__8_, connection_3__18__7_,
         connection_3__18__6_, connection_3__18__5_, connection_3__18__4_,
         connection_3__18__3_, connection_3__18__2_, connection_3__18__1_,
         connection_3__18__0_, connection_3__19__31_, connection_3__19__30_,
         connection_3__19__29_, connection_3__19__28_, connection_3__19__27_,
         connection_3__19__26_, connection_3__19__25_, connection_3__19__24_,
         connection_3__19__23_, connection_3__19__22_, connection_3__19__21_,
         connection_3__19__20_, connection_3__19__19_, connection_3__19__18_,
         connection_3__19__17_, connection_3__19__16_, connection_3__19__15_,
         connection_3__19__14_, connection_3__19__13_, connection_3__19__12_,
         connection_3__19__11_, connection_3__19__10_, connection_3__19__9_,
         connection_3__19__8_, connection_3__19__7_, connection_3__19__6_,
         connection_3__19__5_, connection_3__19__4_, connection_3__19__3_,
         connection_3__19__2_, connection_3__19__1_, connection_3__19__0_,
         connection_3__20__31_, connection_3__20__30_, connection_3__20__29_,
         connection_3__20__28_, connection_3__20__27_, connection_3__20__26_,
         connection_3__20__25_, connection_3__20__24_, connection_3__20__23_,
         connection_3__20__22_, connection_3__20__21_, connection_3__20__20_,
         connection_3__20__19_, connection_3__20__18_, connection_3__20__17_,
         connection_3__20__16_, connection_3__20__15_, connection_3__20__14_,
         connection_3__20__13_, connection_3__20__12_, connection_3__20__11_,
         connection_3__20__10_, connection_3__20__9_, connection_3__20__8_,
         connection_3__20__7_, connection_3__20__6_, connection_3__20__5_,
         connection_3__20__4_, connection_3__20__3_, connection_3__20__2_,
         connection_3__20__1_, connection_3__20__0_, connection_3__21__31_,
         connection_3__21__30_, connection_3__21__29_, connection_3__21__28_,
         connection_3__21__27_, connection_3__21__26_, connection_3__21__25_,
         connection_3__21__24_, connection_3__21__23_, connection_3__21__22_,
         connection_3__21__21_, connection_3__21__20_, connection_3__21__19_,
         connection_3__21__18_, connection_3__21__17_, connection_3__21__16_,
         connection_3__21__15_, connection_3__21__14_, connection_3__21__13_,
         connection_3__21__12_, connection_3__21__11_, connection_3__21__10_,
         connection_3__21__9_, connection_3__21__8_, connection_3__21__7_,
         connection_3__21__6_, connection_3__21__5_, connection_3__21__4_,
         connection_3__21__3_, connection_3__21__2_, connection_3__21__1_,
         connection_3__21__0_, connection_3__22__31_, connection_3__22__30_,
         connection_3__22__29_, connection_3__22__28_, connection_3__22__27_,
         connection_3__22__26_, connection_3__22__25_, connection_3__22__24_,
         connection_3__22__23_, connection_3__22__22_, connection_3__22__21_,
         connection_3__22__20_, connection_3__22__19_, connection_3__22__18_,
         connection_3__22__17_, connection_3__22__16_, connection_3__22__15_,
         connection_3__22__14_, connection_3__22__13_, connection_3__22__12_,
         connection_3__22__11_, connection_3__22__10_, connection_3__22__9_,
         connection_3__22__8_, connection_3__22__7_, connection_3__22__6_,
         connection_3__22__5_, connection_3__22__4_, connection_3__22__3_,
         connection_3__22__2_, connection_3__22__1_, connection_3__22__0_,
         connection_3__23__31_, connection_3__23__30_, connection_3__23__29_,
         connection_3__23__28_, connection_3__23__27_, connection_3__23__26_,
         connection_3__23__25_, connection_3__23__24_, connection_3__23__23_,
         connection_3__23__22_, connection_3__23__21_, connection_3__23__20_,
         connection_3__23__19_, connection_3__23__18_, connection_3__23__17_,
         connection_3__23__16_, connection_3__23__15_, connection_3__23__14_,
         connection_3__23__13_, connection_3__23__12_, connection_3__23__11_,
         connection_3__23__10_, connection_3__23__9_, connection_3__23__8_,
         connection_3__23__7_, connection_3__23__6_, connection_3__23__5_,
         connection_3__23__4_, connection_3__23__3_, connection_3__23__2_,
         connection_3__23__1_, connection_3__23__0_, connection_3__24__31_,
         connection_3__24__30_, connection_3__24__29_, connection_3__24__28_,
         connection_3__24__27_, connection_3__24__26_, connection_3__24__25_,
         connection_3__24__24_, connection_3__24__23_, connection_3__24__22_,
         connection_3__24__21_, connection_3__24__20_, connection_3__24__19_,
         connection_3__24__18_, connection_3__24__17_, connection_3__24__16_,
         connection_3__24__15_, connection_3__24__14_, connection_3__24__13_,
         connection_3__24__12_, connection_3__24__11_, connection_3__24__10_,
         connection_3__24__9_, connection_3__24__8_, connection_3__24__7_,
         connection_3__24__6_, connection_3__24__5_, connection_3__24__4_,
         connection_3__24__3_, connection_3__24__2_, connection_3__24__1_,
         connection_3__24__0_, connection_3__25__31_, connection_3__25__30_,
         connection_3__25__29_, connection_3__25__28_, connection_3__25__27_,
         connection_3__25__26_, connection_3__25__25_, connection_3__25__24_,
         connection_3__25__23_, connection_3__25__22_, connection_3__25__21_,
         connection_3__25__20_, connection_3__25__19_, connection_3__25__18_,
         connection_3__25__17_, connection_3__25__16_, connection_3__25__15_,
         connection_3__25__14_, connection_3__25__13_, connection_3__25__12_,
         connection_3__25__11_, connection_3__25__10_, connection_3__25__9_,
         connection_3__25__8_, connection_3__25__7_, connection_3__25__6_,
         connection_3__25__5_, connection_3__25__4_, connection_3__25__3_,
         connection_3__25__2_, connection_3__25__1_, connection_3__25__0_,
         connection_3__26__31_, connection_3__26__30_, connection_3__26__29_,
         connection_3__26__28_, connection_3__26__27_, connection_3__26__26_,
         connection_3__26__25_, connection_3__26__24_, connection_3__26__23_,
         connection_3__26__22_, connection_3__26__21_, connection_3__26__20_,
         connection_3__26__19_, connection_3__26__18_, connection_3__26__17_,
         connection_3__26__16_, connection_3__26__15_, connection_3__26__14_,
         connection_3__26__13_, connection_3__26__12_, connection_3__26__11_,
         connection_3__26__10_, connection_3__26__9_, connection_3__26__8_,
         connection_3__26__7_, connection_3__26__6_, connection_3__26__5_,
         connection_3__26__4_, connection_3__26__3_, connection_3__26__2_,
         connection_3__26__1_, connection_3__26__0_, connection_3__27__31_,
         connection_3__27__30_, connection_3__27__29_, connection_3__27__28_,
         connection_3__27__27_, connection_3__27__26_, connection_3__27__25_,
         connection_3__27__24_, connection_3__27__23_, connection_3__27__22_,
         connection_3__27__21_, connection_3__27__20_, connection_3__27__19_,
         connection_3__27__18_, connection_3__27__17_, connection_3__27__16_,
         connection_3__27__15_, connection_3__27__14_, connection_3__27__13_,
         connection_3__27__12_, connection_3__27__11_, connection_3__27__10_,
         connection_3__27__9_, connection_3__27__8_, connection_3__27__7_,
         connection_3__27__6_, connection_3__27__5_, connection_3__27__4_,
         connection_3__27__3_, connection_3__27__2_, connection_3__27__1_,
         connection_3__27__0_, connection_3__28__31_, connection_3__28__30_,
         connection_3__28__29_, connection_3__28__28_, connection_3__28__27_,
         connection_3__28__26_, connection_3__28__25_, connection_3__28__24_,
         connection_3__28__23_, connection_3__28__22_, connection_3__28__21_,
         connection_3__28__20_, connection_3__28__19_, connection_3__28__18_,
         connection_3__28__17_, connection_3__28__16_, connection_3__28__15_,
         connection_3__28__14_, connection_3__28__13_, connection_3__28__12_,
         connection_3__28__11_, connection_3__28__10_, connection_3__28__9_,
         connection_3__28__8_, connection_3__28__7_, connection_3__28__6_,
         connection_3__28__5_, connection_3__28__4_, connection_3__28__3_,
         connection_3__28__2_, connection_3__28__1_, connection_3__28__0_,
         connection_3__29__31_, connection_3__29__30_, connection_3__29__29_,
         connection_3__29__28_, connection_3__29__27_, connection_3__29__26_,
         connection_3__29__25_, connection_3__29__24_, connection_3__29__23_,
         connection_3__29__22_, connection_3__29__21_, connection_3__29__20_,
         connection_3__29__19_, connection_3__29__18_, connection_3__29__17_,
         connection_3__29__16_, connection_3__29__15_, connection_3__29__14_,
         connection_3__29__13_, connection_3__29__12_, connection_3__29__11_,
         connection_3__29__10_, connection_3__29__9_, connection_3__29__8_,
         connection_3__29__7_, connection_3__29__6_, connection_3__29__5_,
         connection_3__29__4_, connection_3__29__3_, connection_3__29__2_,
         connection_3__29__1_, connection_3__29__0_, connection_3__30__31_,
         connection_3__30__30_, connection_3__30__29_, connection_3__30__28_,
         connection_3__30__27_, connection_3__30__26_, connection_3__30__25_,
         connection_3__30__24_, connection_3__30__23_, connection_3__30__22_,
         connection_3__30__21_, connection_3__30__20_, connection_3__30__19_,
         connection_3__30__18_, connection_3__30__17_, connection_3__30__16_,
         connection_3__30__15_, connection_3__30__14_, connection_3__30__13_,
         connection_3__30__12_, connection_3__30__11_, connection_3__30__10_,
         connection_3__30__9_, connection_3__30__8_, connection_3__30__7_,
         connection_3__30__6_, connection_3__30__5_, connection_3__30__4_,
         connection_3__30__3_, connection_3__30__2_, connection_3__30__1_,
         connection_3__30__0_, connection_3__31__31_, connection_3__31__30_,
         connection_3__31__29_, connection_3__31__28_, connection_3__31__27_,
         connection_3__31__26_, connection_3__31__25_, connection_3__31__24_,
         connection_3__31__23_, connection_3__31__22_, connection_3__31__21_,
         connection_3__31__20_, connection_3__31__19_, connection_3__31__18_,
         connection_3__31__17_, connection_3__31__16_, connection_3__31__15_,
         connection_3__31__14_, connection_3__31__13_, connection_3__31__12_,
         connection_3__31__11_, connection_3__31__10_, connection_3__31__9_,
         connection_3__31__8_, connection_3__31__7_, connection_3__31__6_,
         connection_3__31__5_, connection_3__31__4_, connection_3__31__3_,
         connection_3__31__2_, connection_3__31__1_, connection_3__31__0_,
         connection_4__0__31_, connection_4__0__30_, connection_4__0__29_,
         connection_4__0__28_, connection_4__0__27_, connection_4__0__26_,
         connection_4__0__25_, connection_4__0__24_, connection_4__0__23_,
         connection_4__0__22_, connection_4__0__21_, connection_4__0__20_,
         connection_4__0__19_, connection_4__0__18_, connection_4__0__17_,
         connection_4__0__16_, connection_4__0__15_, connection_4__0__14_,
         connection_4__0__13_, connection_4__0__12_, connection_4__0__11_,
         connection_4__0__10_, connection_4__0__9_, connection_4__0__8_,
         connection_4__0__7_, connection_4__0__6_, connection_4__0__5_,
         connection_4__0__4_, connection_4__0__3_, connection_4__0__2_,
         connection_4__0__1_, connection_4__0__0_, connection_4__1__31_,
         connection_4__1__30_, connection_4__1__29_, connection_4__1__28_,
         connection_4__1__27_, connection_4__1__26_, connection_4__1__25_,
         connection_4__1__24_, connection_4__1__23_, connection_4__1__22_,
         connection_4__1__21_, connection_4__1__20_, connection_4__1__19_,
         connection_4__1__18_, connection_4__1__17_, connection_4__1__16_,
         connection_4__1__15_, connection_4__1__14_, connection_4__1__13_,
         connection_4__1__12_, connection_4__1__11_, connection_4__1__10_,
         connection_4__1__9_, connection_4__1__8_, connection_4__1__7_,
         connection_4__1__6_, connection_4__1__5_, connection_4__1__4_,
         connection_4__1__3_, connection_4__1__2_, connection_4__1__1_,
         connection_4__1__0_, connection_4__2__31_, connection_4__2__30_,
         connection_4__2__29_, connection_4__2__28_, connection_4__2__27_,
         connection_4__2__26_, connection_4__2__25_, connection_4__2__24_,
         connection_4__2__23_, connection_4__2__22_, connection_4__2__21_,
         connection_4__2__20_, connection_4__2__19_, connection_4__2__18_,
         connection_4__2__17_, connection_4__2__16_, connection_4__2__15_,
         connection_4__2__14_, connection_4__2__13_, connection_4__2__12_,
         connection_4__2__11_, connection_4__2__10_, connection_4__2__9_,
         connection_4__2__8_, connection_4__2__7_, connection_4__2__6_,
         connection_4__2__5_, connection_4__2__4_, connection_4__2__3_,
         connection_4__2__2_, connection_4__2__1_, connection_4__2__0_,
         connection_4__3__31_, connection_4__3__30_, connection_4__3__29_,
         connection_4__3__28_, connection_4__3__27_, connection_4__3__26_,
         connection_4__3__25_, connection_4__3__24_, connection_4__3__23_,
         connection_4__3__22_, connection_4__3__21_, connection_4__3__20_,
         connection_4__3__19_, connection_4__3__18_, connection_4__3__17_,
         connection_4__3__16_, connection_4__3__15_, connection_4__3__14_,
         connection_4__3__13_, connection_4__3__12_, connection_4__3__11_,
         connection_4__3__10_, connection_4__3__9_, connection_4__3__8_,
         connection_4__3__7_, connection_4__3__6_, connection_4__3__5_,
         connection_4__3__4_, connection_4__3__3_, connection_4__3__2_,
         connection_4__3__1_, connection_4__3__0_, connection_4__4__31_,
         connection_4__4__30_, connection_4__4__29_, connection_4__4__28_,
         connection_4__4__27_, connection_4__4__26_, connection_4__4__25_,
         connection_4__4__24_, connection_4__4__23_, connection_4__4__22_,
         connection_4__4__21_, connection_4__4__20_, connection_4__4__19_,
         connection_4__4__18_, connection_4__4__17_, connection_4__4__16_,
         connection_4__4__15_, connection_4__4__14_, connection_4__4__13_,
         connection_4__4__12_, connection_4__4__11_, connection_4__4__10_,
         connection_4__4__9_, connection_4__4__8_, connection_4__4__7_,
         connection_4__4__6_, connection_4__4__5_, connection_4__4__4_,
         connection_4__4__3_, connection_4__4__2_, connection_4__4__1_,
         connection_4__4__0_, connection_4__5__31_, connection_4__5__30_,
         connection_4__5__29_, connection_4__5__28_, connection_4__5__27_,
         connection_4__5__26_, connection_4__5__25_, connection_4__5__24_,
         connection_4__5__23_, connection_4__5__22_, connection_4__5__21_,
         connection_4__5__20_, connection_4__5__19_, connection_4__5__18_,
         connection_4__5__17_, connection_4__5__16_, connection_4__5__15_,
         connection_4__5__14_, connection_4__5__13_, connection_4__5__12_,
         connection_4__5__11_, connection_4__5__10_, connection_4__5__9_,
         connection_4__5__8_, connection_4__5__7_, connection_4__5__6_,
         connection_4__5__5_, connection_4__5__4_, connection_4__5__3_,
         connection_4__5__2_, connection_4__5__1_, connection_4__5__0_,
         connection_4__6__31_, connection_4__6__30_, connection_4__6__29_,
         connection_4__6__28_, connection_4__6__27_, connection_4__6__26_,
         connection_4__6__25_, connection_4__6__24_, connection_4__6__23_,
         connection_4__6__22_, connection_4__6__21_, connection_4__6__20_,
         connection_4__6__19_, connection_4__6__18_, connection_4__6__17_,
         connection_4__6__16_, connection_4__6__15_, connection_4__6__14_,
         connection_4__6__13_, connection_4__6__12_, connection_4__6__11_,
         connection_4__6__10_, connection_4__6__9_, connection_4__6__8_,
         connection_4__6__7_, connection_4__6__6_, connection_4__6__5_,
         connection_4__6__4_, connection_4__6__3_, connection_4__6__2_,
         connection_4__6__1_, connection_4__6__0_, connection_4__7__31_,
         connection_4__7__30_, connection_4__7__29_, connection_4__7__28_,
         connection_4__7__27_, connection_4__7__26_, connection_4__7__25_,
         connection_4__7__24_, connection_4__7__23_, connection_4__7__22_,
         connection_4__7__21_, connection_4__7__20_, connection_4__7__19_,
         connection_4__7__18_, connection_4__7__17_, connection_4__7__16_,
         connection_4__7__15_, connection_4__7__14_, connection_4__7__13_,
         connection_4__7__12_, connection_4__7__11_, connection_4__7__10_,
         connection_4__7__9_, connection_4__7__8_, connection_4__7__7_,
         connection_4__7__6_, connection_4__7__5_, connection_4__7__4_,
         connection_4__7__3_, connection_4__7__2_, connection_4__7__1_,
         connection_4__7__0_, connection_4__8__31_, connection_4__8__30_,
         connection_4__8__29_, connection_4__8__28_, connection_4__8__27_,
         connection_4__8__26_, connection_4__8__25_, connection_4__8__24_,
         connection_4__8__23_, connection_4__8__22_, connection_4__8__21_,
         connection_4__8__20_, connection_4__8__19_, connection_4__8__18_,
         connection_4__8__17_, connection_4__8__16_, connection_4__8__15_,
         connection_4__8__14_, connection_4__8__13_, connection_4__8__12_,
         connection_4__8__11_, connection_4__8__10_, connection_4__8__9_,
         connection_4__8__8_, connection_4__8__7_, connection_4__8__6_,
         connection_4__8__5_, connection_4__8__4_, connection_4__8__3_,
         connection_4__8__2_, connection_4__8__1_, connection_4__8__0_,
         connection_4__9__31_, connection_4__9__30_, connection_4__9__29_,
         connection_4__9__28_, connection_4__9__27_, connection_4__9__26_,
         connection_4__9__25_, connection_4__9__24_, connection_4__9__23_,
         connection_4__9__22_, connection_4__9__21_, connection_4__9__20_,
         connection_4__9__19_, connection_4__9__18_, connection_4__9__17_,
         connection_4__9__16_, connection_4__9__15_, connection_4__9__14_,
         connection_4__9__13_, connection_4__9__12_, connection_4__9__11_,
         connection_4__9__10_, connection_4__9__9_, connection_4__9__8_,
         connection_4__9__7_, connection_4__9__6_, connection_4__9__5_,
         connection_4__9__4_, connection_4__9__3_, connection_4__9__2_,
         connection_4__9__1_, connection_4__9__0_, connection_4__10__31_,
         connection_4__10__30_, connection_4__10__29_, connection_4__10__28_,
         connection_4__10__27_, connection_4__10__26_, connection_4__10__25_,
         connection_4__10__24_, connection_4__10__23_, connection_4__10__22_,
         connection_4__10__21_, connection_4__10__20_, connection_4__10__19_,
         connection_4__10__18_, connection_4__10__17_, connection_4__10__16_,
         connection_4__10__15_, connection_4__10__14_, connection_4__10__13_,
         connection_4__10__12_, connection_4__10__11_, connection_4__10__10_,
         connection_4__10__9_, connection_4__10__8_, connection_4__10__7_,
         connection_4__10__6_, connection_4__10__5_, connection_4__10__4_,
         connection_4__10__3_, connection_4__10__2_, connection_4__10__1_,
         connection_4__10__0_, connection_4__11__31_, connection_4__11__30_,
         connection_4__11__29_, connection_4__11__28_, connection_4__11__27_,
         connection_4__11__26_, connection_4__11__25_, connection_4__11__24_,
         connection_4__11__23_, connection_4__11__22_, connection_4__11__21_,
         connection_4__11__20_, connection_4__11__19_, connection_4__11__18_,
         connection_4__11__17_, connection_4__11__16_, connection_4__11__15_,
         connection_4__11__14_, connection_4__11__13_, connection_4__11__12_,
         connection_4__11__11_, connection_4__11__10_, connection_4__11__9_,
         connection_4__11__8_, connection_4__11__7_, connection_4__11__6_,
         connection_4__11__5_, connection_4__11__4_, connection_4__11__3_,
         connection_4__11__2_, connection_4__11__1_, connection_4__11__0_,
         connection_4__12__31_, connection_4__12__30_, connection_4__12__29_,
         connection_4__12__28_, connection_4__12__27_, connection_4__12__26_,
         connection_4__12__25_, connection_4__12__24_, connection_4__12__23_,
         connection_4__12__22_, connection_4__12__21_, connection_4__12__20_,
         connection_4__12__19_, connection_4__12__18_, connection_4__12__17_,
         connection_4__12__16_, connection_4__12__15_, connection_4__12__14_,
         connection_4__12__13_, connection_4__12__12_, connection_4__12__11_,
         connection_4__12__10_, connection_4__12__9_, connection_4__12__8_,
         connection_4__12__7_, connection_4__12__6_, connection_4__12__5_,
         connection_4__12__4_, connection_4__12__3_, connection_4__12__2_,
         connection_4__12__1_, connection_4__12__0_, connection_4__13__31_,
         connection_4__13__30_, connection_4__13__29_, connection_4__13__28_,
         connection_4__13__27_, connection_4__13__26_, connection_4__13__25_,
         connection_4__13__24_, connection_4__13__23_, connection_4__13__22_,
         connection_4__13__21_, connection_4__13__20_, connection_4__13__19_,
         connection_4__13__18_, connection_4__13__17_, connection_4__13__16_,
         connection_4__13__15_, connection_4__13__14_, connection_4__13__13_,
         connection_4__13__12_, connection_4__13__11_, connection_4__13__10_,
         connection_4__13__9_, connection_4__13__8_, connection_4__13__7_,
         connection_4__13__6_, connection_4__13__5_, connection_4__13__4_,
         connection_4__13__3_, connection_4__13__2_, connection_4__13__1_,
         connection_4__13__0_, connection_4__14__31_, connection_4__14__30_,
         connection_4__14__29_, connection_4__14__28_, connection_4__14__27_,
         connection_4__14__26_, connection_4__14__25_, connection_4__14__24_,
         connection_4__14__23_, connection_4__14__22_, connection_4__14__21_,
         connection_4__14__20_, connection_4__14__19_, connection_4__14__18_,
         connection_4__14__17_, connection_4__14__16_, connection_4__14__15_,
         connection_4__14__14_, connection_4__14__13_, connection_4__14__12_,
         connection_4__14__11_, connection_4__14__10_, connection_4__14__9_,
         connection_4__14__8_, connection_4__14__7_, connection_4__14__6_,
         connection_4__14__5_, connection_4__14__4_, connection_4__14__3_,
         connection_4__14__2_, connection_4__14__1_, connection_4__14__0_,
         connection_4__15__31_, connection_4__15__30_, connection_4__15__29_,
         connection_4__15__28_, connection_4__15__27_, connection_4__15__26_,
         connection_4__15__25_, connection_4__15__24_, connection_4__15__23_,
         connection_4__15__22_, connection_4__15__21_, connection_4__15__20_,
         connection_4__15__19_, connection_4__15__18_, connection_4__15__17_,
         connection_4__15__16_, connection_4__15__15_, connection_4__15__14_,
         connection_4__15__13_, connection_4__15__12_, connection_4__15__11_,
         connection_4__15__10_, connection_4__15__9_, connection_4__15__8_,
         connection_4__15__7_, connection_4__15__6_, connection_4__15__5_,
         connection_4__15__4_, connection_4__15__3_, connection_4__15__2_,
         connection_4__15__1_, connection_4__15__0_, connection_4__16__31_,
         connection_4__16__30_, connection_4__16__29_, connection_4__16__28_,
         connection_4__16__27_, connection_4__16__26_, connection_4__16__25_,
         connection_4__16__24_, connection_4__16__23_, connection_4__16__22_,
         connection_4__16__21_, connection_4__16__20_, connection_4__16__19_,
         connection_4__16__18_, connection_4__16__17_, connection_4__16__16_,
         connection_4__16__15_, connection_4__16__14_, connection_4__16__13_,
         connection_4__16__12_, connection_4__16__11_, connection_4__16__10_,
         connection_4__16__9_, connection_4__16__8_, connection_4__16__7_,
         connection_4__16__6_, connection_4__16__5_, connection_4__16__4_,
         connection_4__16__3_, connection_4__16__2_, connection_4__16__1_,
         connection_4__16__0_, connection_4__17__31_, connection_4__17__30_,
         connection_4__17__29_, connection_4__17__28_, connection_4__17__27_,
         connection_4__17__26_, connection_4__17__25_, connection_4__17__24_,
         connection_4__17__23_, connection_4__17__22_, connection_4__17__21_,
         connection_4__17__20_, connection_4__17__19_, connection_4__17__18_,
         connection_4__17__17_, connection_4__17__16_, connection_4__17__15_,
         connection_4__17__14_, connection_4__17__13_, connection_4__17__12_,
         connection_4__17__11_, connection_4__17__10_, connection_4__17__9_,
         connection_4__17__8_, connection_4__17__7_, connection_4__17__6_,
         connection_4__17__5_, connection_4__17__4_, connection_4__17__3_,
         connection_4__17__2_, connection_4__17__1_, connection_4__17__0_,
         connection_4__18__31_, connection_4__18__30_, connection_4__18__29_,
         connection_4__18__28_, connection_4__18__27_, connection_4__18__26_,
         connection_4__18__25_, connection_4__18__24_, connection_4__18__23_,
         connection_4__18__22_, connection_4__18__21_, connection_4__18__20_,
         connection_4__18__19_, connection_4__18__18_, connection_4__18__17_,
         connection_4__18__16_, connection_4__18__15_, connection_4__18__14_,
         connection_4__18__13_, connection_4__18__12_, connection_4__18__11_,
         connection_4__18__10_, connection_4__18__9_, connection_4__18__8_,
         connection_4__18__7_, connection_4__18__6_, connection_4__18__5_,
         connection_4__18__4_, connection_4__18__3_, connection_4__18__2_,
         connection_4__18__1_, connection_4__18__0_, connection_4__19__31_,
         connection_4__19__30_, connection_4__19__29_, connection_4__19__28_,
         connection_4__19__27_, connection_4__19__26_, connection_4__19__25_,
         connection_4__19__24_, connection_4__19__23_, connection_4__19__22_,
         connection_4__19__21_, connection_4__19__20_, connection_4__19__19_,
         connection_4__19__18_, connection_4__19__17_, connection_4__19__16_,
         connection_4__19__15_, connection_4__19__14_, connection_4__19__13_,
         connection_4__19__12_, connection_4__19__11_, connection_4__19__10_,
         connection_4__19__9_, connection_4__19__8_, connection_4__19__7_,
         connection_4__19__6_, connection_4__19__5_, connection_4__19__4_,
         connection_4__19__3_, connection_4__19__2_, connection_4__19__1_,
         connection_4__19__0_, connection_4__20__31_, connection_4__20__30_,
         connection_4__20__29_, connection_4__20__28_, connection_4__20__27_,
         connection_4__20__26_, connection_4__20__25_, connection_4__20__24_,
         connection_4__20__23_, connection_4__20__22_, connection_4__20__21_,
         connection_4__20__20_, connection_4__20__19_, connection_4__20__18_,
         connection_4__20__17_, connection_4__20__16_, connection_4__20__15_,
         connection_4__20__14_, connection_4__20__13_, connection_4__20__12_,
         connection_4__20__11_, connection_4__20__10_, connection_4__20__9_,
         connection_4__20__8_, connection_4__20__7_, connection_4__20__6_,
         connection_4__20__5_, connection_4__20__4_, connection_4__20__3_,
         connection_4__20__2_, connection_4__20__1_, connection_4__20__0_,
         connection_4__21__31_, connection_4__21__30_, connection_4__21__29_,
         connection_4__21__28_, connection_4__21__27_, connection_4__21__26_,
         connection_4__21__25_, connection_4__21__24_, connection_4__21__23_,
         connection_4__21__22_, connection_4__21__21_, connection_4__21__20_,
         connection_4__21__19_, connection_4__21__18_, connection_4__21__17_,
         connection_4__21__16_, connection_4__21__15_, connection_4__21__14_,
         connection_4__21__13_, connection_4__21__12_, connection_4__21__11_,
         connection_4__21__10_, connection_4__21__9_, connection_4__21__8_,
         connection_4__21__7_, connection_4__21__6_, connection_4__21__5_,
         connection_4__21__4_, connection_4__21__3_, connection_4__21__2_,
         connection_4__21__1_, connection_4__21__0_, connection_4__22__31_,
         connection_4__22__30_, connection_4__22__29_, connection_4__22__28_,
         connection_4__22__27_, connection_4__22__26_, connection_4__22__25_,
         connection_4__22__24_, connection_4__22__23_, connection_4__22__22_,
         connection_4__22__21_, connection_4__22__20_, connection_4__22__19_,
         connection_4__22__18_, connection_4__22__17_, connection_4__22__16_,
         connection_4__22__15_, connection_4__22__14_, connection_4__22__13_,
         connection_4__22__12_, connection_4__22__11_, connection_4__22__10_,
         connection_4__22__9_, connection_4__22__8_, connection_4__22__7_,
         connection_4__22__6_, connection_4__22__5_, connection_4__22__4_,
         connection_4__22__3_, connection_4__22__2_, connection_4__22__1_,
         connection_4__22__0_, connection_4__23__31_, connection_4__23__30_,
         connection_4__23__29_, connection_4__23__28_, connection_4__23__27_,
         connection_4__23__26_, connection_4__23__25_, connection_4__23__24_,
         connection_4__23__23_, connection_4__23__22_, connection_4__23__21_,
         connection_4__23__20_, connection_4__23__19_, connection_4__23__18_,
         connection_4__23__17_, connection_4__23__16_, connection_4__23__15_,
         connection_4__23__14_, connection_4__23__13_, connection_4__23__12_,
         connection_4__23__11_, connection_4__23__10_, connection_4__23__9_,
         connection_4__23__8_, connection_4__23__7_, connection_4__23__6_,
         connection_4__23__5_, connection_4__23__4_, connection_4__23__3_,
         connection_4__23__2_, connection_4__23__1_, connection_4__23__0_,
         connection_4__24__31_, connection_4__24__30_, connection_4__24__29_,
         connection_4__24__28_, connection_4__24__27_, connection_4__24__26_,
         connection_4__24__25_, connection_4__24__24_, connection_4__24__23_,
         connection_4__24__22_, connection_4__24__21_, connection_4__24__20_,
         connection_4__24__19_, connection_4__24__18_, connection_4__24__17_,
         connection_4__24__16_, connection_4__24__15_, connection_4__24__14_,
         connection_4__24__13_, connection_4__24__12_, connection_4__24__11_,
         connection_4__24__10_, connection_4__24__9_, connection_4__24__8_,
         connection_4__24__7_, connection_4__24__6_, connection_4__24__5_,
         connection_4__24__4_, connection_4__24__3_, connection_4__24__2_,
         connection_4__24__1_, connection_4__24__0_, connection_4__25__31_,
         connection_4__25__30_, connection_4__25__29_, connection_4__25__28_,
         connection_4__25__27_, connection_4__25__26_, connection_4__25__25_,
         connection_4__25__24_, connection_4__25__23_, connection_4__25__22_,
         connection_4__25__21_, connection_4__25__20_, connection_4__25__19_,
         connection_4__25__18_, connection_4__25__17_, connection_4__25__16_,
         connection_4__25__15_, connection_4__25__14_, connection_4__25__13_,
         connection_4__25__12_, connection_4__25__11_, connection_4__25__10_,
         connection_4__25__9_, connection_4__25__8_, connection_4__25__7_,
         connection_4__25__6_, connection_4__25__5_, connection_4__25__4_,
         connection_4__25__3_, connection_4__25__2_, connection_4__25__1_,
         connection_4__25__0_, connection_4__26__31_, connection_4__26__30_,
         connection_4__26__29_, connection_4__26__28_, connection_4__26__27_,
         connection_4__26__26_, connection_4__26__25_, connection_4__26__24_,
         connection_4__26__23_, connection_4__26__22_, connection_4__26__21_,
         connection_4__26__20_, connection_4__26__19_, connection_4__26__18_,
         connection_4__26__17_, connection_4__26__16_, connection_4__26__15_,
         connection_4__26__14_, connection_4__26__13_, connection_4__26__12_,
         connection_4__26__11_, connection_4__26__10_, connection_4__26__9_,
         connection_4__26__8_, connection_4__26__7_, connection_4__26__6_,
         connection_4__26__5_, connection_4__26__4_, connection_4__26__3_,
         connection_4__26__2_, connection_4__26__1_, connection_4__26__0_,
         connection_4__27__31_, connection_4__27__30_, connection_4__27__29_,
         connection_4__27__28_, connection_4__27__27_, connection_4__27__26_,
         connection_4__27__25_, connection_4__27__24_, connection_4__27__23_,
         connection_4__27__22_, connection_4__27__21_, connection_4__27__20_,
         connection_4__27__19_, connection_4__27__18_, connection_4__27__17_,
         connection_4__27__16_, connection_4__27__15_, connection_4__27__14_,
         connection_4__27__13_, connection_4__27__12_, connection_4__27__11_,
         connection_4__27__10_, connection_4__27__9_, connection_4__27__8_,
         connection_4__27__7_, connection_4__27__6_, connection_4__27__5_,
         connection_4__27__4_, connection_4__27__3_, connection_4__27__2_,
         connection_4__27__1_, connection_4__27__0_, connection_4__28__31_,
         connection_4__28__30_, connection_4__28__29_, connection_4__28__28_,
         connection_4__28__27_, connection_4__28__26_, connection_4__28__25_,
         connection_4__28__24_, connection_4__28__23_, connection_4__28__22_,
         connection_4__28__21_, connection_4__28__20_, connection_4__28__19_,
         connection_4__28__18_, connection_4__28__17_, connection_4__28__16_,
         connection_4__28__15_, connection_4__28__14_, connection_4__28__13_,
         connection_4__28__12_, connection_4__28__11_, connection_4__28__10_,
         connection_4__28__9_, connection_4__28__8_, connection_4__28__7_,
         connection_4__28__6_, connection_4__28__5_, connection_4__28__4_,
         connection_4__28__3_, connection_4__28__2_, connection_4__28__1_,
         connection_4__28__0_, connection_4__29__31_, connection_4__29__30_,
         connection_4__29__29_, connection_4__29__28_, connection_4__29__27_,
         connection_4__29__26_, connection_4__29__25_, connection_4__29__24_,
         connection_4__29__23_, connection_4__29__22_, connection_4__29__21_,
         connection_4__29__20_, connection_4__29__19_, connection_4__29__18_,
         connection_4__29__17_, connection_4__29__16_, connection_4__29__15_,
         connection_4__29__14_, connection_4__29__13_, connection_4__29__12_,
         connection_4__29__11_, connection_4__29__10_, connection_4__29__9_,
         connection_4__29__8_, connection_4__29__7_, connection_4__29__6_,
         connection_4__29__5_, connection_4__29__4_, connection_4__29__3_,
         connection_4__29__2_, connection_4__29__1_, connection_4__29__0_,
         connection_4__30__31_, connection_4__30__30_, connection_4__30__29_,
         connection_4__30__28_, connection_4__30__27_, connection_4__30__26_,
         connection_4__30__25_, connection_4__30__24_, connection_4__30__23_,
         connection_4__30__22_, connection_4__30__21_, connection_4__30__20_,
         connection_4__30__19_, connection_4__30__18_, connection_4__30__17_,
         connection_4__30__16_, connection_4__30__15_, connection_4__30__14_,
         connection_4__30__13_, connection_4__30__12_, connection_4__30__11_,
         connection_4__30__10_, connection_4__30__9_, connection_4__30__8_,
         connection_4__30__7_, connection_4__30__6_, connection_4__30__5_,
         connection_4__30__4_, connection_4__30__3_, connection_4__30__2_,
         connection_4__30__1_, connection_4__30__0_, connection_4__31__31_,
         connection_4__31__30_, connection_4__31__29_, connection_4__31__28_,
         connection_4__31__27_, connection_4__31__26_, connection_4__31__25_,
         connection_4__31__24_, connection_4__31__23_, connection_4__31__22_,
         connection_4__31__21_, connection_4__31__20_, connection_4__31__19_,
         connection_4__31__18_, connection_4__31__17_, connection_4__31__16_,
         connection_4__31__15_, connection_4__31__14_, connection_4__31__13_,
         connection_4__31__12_, connection_4__31__11_, connection_4__31__10_,
         connection_4__31__9_, connection_4__31__8_, connection_4__31__7_,
         connection_4__31__6_, connection_4__31__5_, connection_4__31__4_,
         connection_4__31__3_, connection_4__31__2_, connection_4__31__1_,
         connection_4__31__0_, connection_5__0__31_, connection_5__0__30_,
         connection_5__0__29_, connection_5__0__28_, connection_5__0__27_,
         connection_5__0__26_, connection_5__0__25_, connection_5__0__24_,
         connection_5__0__23_, connection_5__0__22_, connection_5__0__21_,
         connection_5__0__20_, connection_5__0__19_, connection_5__0__18_,
         connection_5__0__17_, connection_5__0__16_, connection_5__0__15_,
         connection_5__0__14_, connection_5__0__13_, connection_5__0__12_,
         connection_5__0__11_, connection_5__0__10_, connection_5__0__9_,
         connection_5__0__8_, connection_5__0__7_, connection_5__0__6_,
         connection_5__0__5_, connection_5__0__4_, connection_5__0__3_,
         connection_5__0__2_, connection_5__0__1_, connection_5__0__0_,
         connection_5__1__31_, connection_5__1__30_, connection_5__1__29_,
         connection_5__1__28_, connection_5__1__27_, connection_5__1__26_,
         connection_5__1__25_, connection_5__1__24_, connection_5__1__23_,
         connection_5__1__22_, connection_5__1__21_, connection_5__1__20_,
         connection_5__1__19_, connection_5__1__18_, connection_5__1__17_,
         connection_5__1__16_, connection_5__1__15_, connection_5__1__14_,
         connection_5__1__13_, connection_5__1__12_, connection_5__1__11_,
         connection_5__1__10_, connection_5__1__9_, connection_5__1__8_,
         connection_5__1__7_, connection_5__1__6_, connection_5__1__5_,
         connection_5__1__4_, connection_5__1__3_, connection_5__1__2_,
         connection_5__1__1_, connection_5__1__0_, connection_5__2__31_,
         connection_5__2__30_, connection_5__2__29_, connection_5__2__28_,
         connection_5__2__27_, connection_5__2__26_, connection_5__2__25_,
         connection_5__2__24_, connection_5__2__23_, connection_5__2__22_,
         connection_5__2__21_, connection_5__2__20_, connection_5__2__19_,
         connection_5__2__18_, connection_5__2__17_, connection_5__2__16_,
         connection_5__2__15_, connection_5__2__14_, connection_5__2__13_,
         connection_5__2__12_, connection_5__2__11_, connection_5__2__10_,
         connection_5__2__9_, connection_5__2__8_, connection_5__2__7_,
         connection_5__2__6_, connection_5__2__5_, connection_5__2__4_,
         connection_5__2__3_, connection_5__2__2_, connection_5__2__1_,
         connection_5__2__0_, connection_5__3__31_, connection_5__3__30_,
         connection_5__3__29_, connection_5__3__28_, connection_5__3__27_,
         connection_5__3__26_, connection_5__3__25_, connection_5__3__24_,
         connection_5__3__23_, connection_5__3__22_, connection_5__3__21_,
         connection_5__3__20_, connection_5__3__19_, connection_5__3__18_,
         connection_5__3__17_, connection_5__3__16_, connection_5__3__15_,
         connection_5__3__14_, connection_5__3__13_, connection_5__3__12_,
         connection_5__3__11_, connection_5__3__10_, connection_5__3__9_,
         connection_5__3__8_, connection_5__3__7_, connection_5__3__6_,
         connection_5__3__5_, connection_5__3__4_, connection_5__3__3_,
         connection_5__3__2_, connection_5__3__1_, connection_5__3__0_,
         connection_5__4__31_, connection_5__4__30_, connection_5__4__29_,
         connection_5__4__28_, connection_5__4__27_, connection_5__4__26_,
         connection_5__4__25_, connection_5__4__24_, connection_5__4__23_,
         connection_5__4__22_, connection_5__4__21_, connection_5__4__20_,
         connection_5__4__19_, connection_5__4__18_, connection_5__4__17_,
         connection_5__4__16_, connection_5__4__15_, connection_5__4__14_,
         connection_5__4__13_, connection_5__4__12_, connection_5__4__11_,
         connection_5__4__10_, connection_5__4__9_, connection_5__4__8_,
         connection_5__4__7_, connection_5__4__6_, connection_5__4__5_,
         connection_5__4__4_, connection_5__4__3_, connection_5__4__2_,
         connection_5__4__1_, connection_5__4__0_, connection_5__5__31_,
         connection_5__5__30_, connection_5__5__29_, connection_5__5__28_,
         connection_5__5__27_, connection_5__5__26_, connection_5__5__25_,
         connection_5__5__24_, connection_5__5__23_, connection_5__5__22_,
         connection_5__5__21_, connection_5__5__20_, connection_5__5__19_,
         connection_5__5__18_, connection_5__5__17_, connection_5__5__16_,
         connection_5__5__15_, connection_5__5__14_, connection_5__5__13_,
         connection_5__5__12_, connection_5__5__11_, connection_5__5__10_,
         connection_5__5__9_, connection_5__5__8_, connection_5__5__7_,
         connection_5__5__6_, connection_5__5__5_, connection_5__5__4_,
         connection_5__5__3_, connection_5__5__2_, connection_5__5__1_,
         connection_5__5__0_, connection_5__6__31_, connection_5__6__30_,
         connection_5__6__29_, connection_5__6__28_, connection_5__6__27_,
         connection_5__6__26_, connection_5__6__25_, connection_5__6__24_,
         connection_5__6__23_, connection_5__6__22_, connection_5__6__21_,
         connection_5__6__20_, connection_5__6__19_, connection_5__6__18_,
         connection_5__6__17_, connection_5__6__16_, connection_5__6__15_,
         connection_5__6__14_, connection_5__6__13_, connection_5__6__12_,
         connection_5__6__11_, connection_5__6__10_, connection_5__6__9_,
         connection_5__6__8_, connection_5__6__7_, connection_5__6__6_,
         connection_5__6__5_, connection_5__6__4_, connection_5__6__3_,
         connection_5__6__2_, connection_5__6__1_, connection_5__6__0_,
         connection_5__7__31_, connection_5__7__30_, connection_5__7__29_,
         connection_5__7__28_, connection_5__7__27_, connection_5__7__26_,
         connection_5__7__25_, connection_5__7__24_, connection_5__7__23_,
         connection_5__7__22_, connection_5__7__21_, connection_5__7__20_,
         connection_5__7__19_, connection_5__7__18_, connection_5__7__17_,
         connection_5__7__16_, connection_5__7__15_, connection_5__7__14_,
         connection_5__7__13_, connection_5__7__12_, connection_5__7__11_,
         connection_5__7__10_, connection_5__7__9_, connection_5__7__8_,
         connection_5__7__7_, connection_5__7__6_, connection_5__7__5_,
         connection_5__7__4_, connection_5__7__3_, connection_5__7__2_,
         connection_5__7__1_, connection_5__7__0_, connection_5__8__31_,
         connection_5__8__30_, connection_5__8__29_, connection_5__8__28_,
         connection_5__8__27_, connection_5__8__26_, connection_5__8__25_,
         connection_5__8__24_, connection_5__8__23_, connection_5__8__22_,
         connection_5__8__21_, connection_5__8__20_, connection_5__8__19_,
         connection_5__8__18_, connection_5__8__17_, connection_5__8__16_,
         connection_5__8__15_, connection_5__8__14_, connection_5__8__13_,
         connection_5__8__12_, connection_5__8__11_, connection_5__8__10_,
         connection_5__8__9_, connection_5__8__8_, connection_5__8__7_,
         connection_5__8__6_, connection_5__8__5_, connection_5__8__4_,
         connection_5__8__3_, connection_5__8__2_, connection_5__8__1_,
         connection_5__8__0_, connection_5__9__31_, connection_5__9__30_,
         connection_5__9__29_, connection_5__9__28_, connection_5__9__27_,
         connection_5__9__26_, connection_5__9__25_, connection_5__9__24_,
         connection_5__9__23_, connection_5__9__22_, connection_5__9__21_,
         connection_5__9__20_, connection_5__9__19_, connection_5__9__18_,
         connection_5__9__17_, connection_5__9__16_, connection_5__9__15_,
         connection_5__9__14_, connection_5__9__13_, connection_5__9__12_,
         connection_5__9__11_, connection_5__9__10_, connection_5__9__9_,
         connection_5__9__8_, connection_5__9__7_, connection_5__9__6_,
         connection_5__9__5_, connection_5__9__4_, connection_5__9__3_,
         connection_5__9__2_, connection_5__9__1_, connection_5__9__0_,
         connection_5__10__31_, connection_5__10__30_, connection_5__10__29_,
         connection_5__10__28_, connection_5__10__27_, connection_5__10__26_,
         connection_5__10__25_, connection_5__10__24_, connection_5__10__23_,
         connection_5__10__22_, connection_5__10__21_, connection_5__10__20_,
         connection_5__10__19_, connection_5__10__18_, connection_5__10__17_,
         connection_5__10__16_, connection_5__10__15_, connection_5__10__14_,
         connection_5__10__13_, connection_5__10__12_, connection_5__10__11_,
         connection_5__10__10_, connection_5__10__9_, connection_5__10__8_,
         connection_5__10__7_, connection_5__10__6_, connection_5__10__5_,
         connection_5__10__4_, connection_5__10__3_, connection_5__10__2_,
         connection_5__10__1_, connection_5__10__0_, connection_5__11__31_,
         connection_5__11__30_, connection_5__11__29_, connection_5__11__28_,
         connection_5__11__27_, connection_5__11__26_, connection_5__11__25_,
         connection_5__11__24_, connection_5__11__23_, connection_5__11__22_,
         connection_5__11__21_, connection_5__11__20_, connection_5__11__19_,
         connection_5__11__18_, connection_5__11__17_, connection_5__11__16_,
         connection_5__11__15_, connection_5__11__14_, connection_5__11__13_,
         connection_5__11__12_, connection_5__11__11_, connection_5__11__10_,
         connection_5__11__9_, connection_5__11__8_, connection_5__11__7_,
         connection_5__11__6_, connection_5__11__5_, connection_5__11__4_,
         connection_5__11__3_, connection_5__11__2_, connection_5__11__1_,
         connection_5__11__0_, connection_5__12__31_, connection_5__12__30_,
         connection_5__12__29_, connection_5__12__28_, connection_5__12__27_,
         connection_5__12__26_, connection_5__12__25_, connection_5__12__24_,
         connection_5__12__23_, connection_5__12__22_, connection_5__12__21_,
         connection_5__12__20_, connection_5__12__19_, connection_5__12__18_,
         connection_5__12__17_, connection_5__12__16_, connection_5__12__15_,
         connection_5__12__14_, connection_5__12__13_, connection_5__12__12_,
         connection_5__12__11_, connection_5__12__10_, connection_5__12__9_,
         connection_5__12__8_, connection_5__12__7_, connection_5__12__6_,
         connection_5__12__5_, connection_5__12__4_, connection_5__12__3_,
         connection_5__12__2_, connection_5__12__1_, connection_5__12__0_,
         connection_5__13__31_, connection_5__13__30_, connection_5__13__29_,
         connection_5__13__28_, connection_5__13__27_, connection_5__13__26_,
         connection_5__13__25_, connection_5__13__24_, connection_5__13__23_,
         connection_5__13__22_, connection_5__13__21_, connection_5__13__20_,
         connection_5__13__19_, connection_5__13__18_, connection_5__13__17_,
         connection_5__13__16_, connection_5__13__15_, connection_5__13__14_,
         connection_5__13__13_, connection_5__13__12_, connection_5__13__11_,
         connection_5__13__10_, connection_5__13__9_, connection_5__13__8_,
         connection_5__13__7_, connection_5__13__6_, connection_5__13__5_,
         connection_5__13__4_, connection_5__13__3_, connection_5__13__2_,
         connection_5__13__1_, connection_5__13__0_, connection_5__14__31_,
         connection_5__14__30_, connection_5__14__29_, connection_5__14__28_,
         connection_5__14__27_, connection_5__14__26_, connection_5__14__25_,
         connection_5__14__24_, connection_5__14__23_, connection_5__14__22_,
         connection_5__14__21_, connection_5__14__20_, connection_5__14__19_,
         connection_5__14__18_, connection_5__14__17_, connection_5__14__16_,
         connection_5__14__15_, connection_5__14__14_, connection_5__14__13_,
         connection_5__14__12_, connection_5__14__11_, connection_5__14__10_,
         connection_5__14__9_, connection_5__14__8_, connection_5__14__7_,
         connection_5__14__6_, connection_5__14__5_, connection_5__14__4_,
         connection_5__14__3_, connection_5__14__2_, connection_5__14__1_,
         connection_5__14__0_, connection_5__15__31_, connection_5__15__30_,
         connection_5__15__29_, connection_5__15__28_, connection_5__15__27_,
         connection_5__15__26_, connection_5__15__25_, connection_5__15__24_,
         connection_5__15__23_, connection_5__15__22_, connection_5__15__21_,
         connection_5__15__20_, connection_5__15__19_, connection_5__15__18_,
         connection_5__15__17_, connection_5__15__16_, connection_5__15__15_,
         connection_5__15__14_, connection_5__15__13_, connection_5__15__12_,
         connection_5__15__11_, connection_5__15__10_, connection_5__15__9_,
         connection_5__15__8_, connection_5__15__7_, connection_5__15__6_,
         connection_5__15__5_, connection_5__15__4_, connection_5__15__3_,
         connection_5__15__2_, connection_5__15__1_, connection_5__15__0_,
         connection_5__16__31_, connection_5__16__30_, connection_5__16__29_,
         connection_5__16__28_, connection_5__16__27_, connection_5__16__26_,
         connection_5__16__25_, connection_5__16__24_, connection_5__16__23_,
         connection_5__16__22_, connection_5__16__21_, connection_5__16__20_,
         connection_5__16__19_, connection_5__16__18_, connection_5__16__17_,
         connection_5__16__16_, connection_5__16__15_, connection_5__16__14_,
         connection_5__16__13_, connection_5__16__12_, connection_5__16__11_,
         connection_5__16__10_, connection_5__16__9_, connection_5__16__8_,
         connection_5__16__7_, connection_5__16__6_, connection_5__16__5_,
         connection_5__16__4_, connection_5__16__3_, connection_5__16__2_,
         connection_5__16__1_, connection_5__16__0_, connection_5__17__31_,
         connection_5__17__30_, connection_5__17__29_, connection_5__17__28_,
         connection_5__17__27_, connection_5__17__26_, connection_5__17__25_,
         connection_5__17__24_, connection_5__17__23_, connection_5__17__22_,
         connection_5__17__21_, connection_5__17__20_, connection_5__17__19_,
         connection_5__17__18_, connection_5__17__17_, connection_5__17__16_,
         connection_5__17__15_, connection_5__17__14_, connection_5__17__13_,
         connection_5__17__12_, connection_5__17__11_, connection_5__17__10_,
         connection_5__17__9_, connection_5__17__8_, connection_5__17__7_,
         connection_5__17__6_, connection_5__17__5_, connection_5__17__4_,
         connection_5__17__3_, connection_5__17__2_, connection_5__17__1_,
         connection_5__17__0_, connection_5__18__31_, connection_5__18__30_,
         connection_5__18__29_, connection_5__18__28_, connection_5__18__27_,
         connection_5__18__26_, connection_5__18__25_, connection_5__18__24_,
         connection_5__18__23_, connection_5__18__22_, connection_5__18__21_,
         connection_5__18__20_, connection_5__18__19_, connection_5__18__18_,
         connection_5__18__17_, connection_5__18__16_, connection_5__18__15_,
         connection_5__18__14_, connection_5__18__13_, connection_5__18__12_,
         connection_5__18__11_, connection_5__18__10_, connection_5__18__9_,
         connection_5__18__8_, connection_5__18__7_, connection_5__18__6_,
         connection_5__18__5_, connection_5__18__4_, connection_5__18__3_,
         connection_5__18__2_, connection_5__18__1_, connection_5__18__0_,
         connection_5__19__31_, connection_5__19__30_, connection_5__19__29_,
         connection_5__19__28_, connection_5__19__27_, connection_5__19__26_,
         connection_5__19__25_, connection_5__19__24_, connection_5__19__23_,
         connection_5__19__22_, connection_5__19__21_, connection_5__19__20_,
         connection_5__19__19_, connection_5__19__18_, connection_5__19__17_,
         connection_5__19__16_, connection_5__19__15_, connection_5__19__14_,
         connection_5__19__13_, connection_5__19__12_, connection_5__19__11_,
         connection_5__19__10_, connection_5__19__9_, connection_5__19__8_,
         connection_5__19__7_, connection_5__19__6_, connection_5__19__5_,
         connection_5__19__4_, connection_5__19__3_, connection_5__19__2_,
         connection_5__19__1_, connection_5__19__0_, connection_5__20__31_,
         connection_5__20__30_, connection_5__20__29_, connection_5__20__28_,
         connection_5__20__27_, connection_5__20__26_, connection_5__20__25_,
         connection_5__20__24_, connection_5__20__23_, connection_5__20__22_,
         connection_5__20__21_, connection_5__20__20_, connection_5__20__19_,
         connection_5__20__18_, connection_5__20__17_, connection_5__20__16_,
         connection_5__20__15_, connection_5__20__14_, connection_5__20__13_,
         connection_5__20__12_, connection_5__20__11_, connection_5__20__10_,
         connection_5__20__9_, connection_5__20__8_, connection_5__20__7_,
         connection_5__20__6_, connection_5__20__5_, connection_5__20__4_,
         connection_5__20__3_, connection_5__20__2_, connection_5__20__1_,
         connection_5__20__0_, connection_5__21__31_, connection_5__21__30_,
         connection_5__21__29_, connection_5__21__28_, connection_5__21__27_,
         connection_5__21__26_, connection_5__21__25_, connection_5__21__24_,
         connection_5__21__23_, connection_5__21__22_, connection_5__21__21_,
         connection_5__21__20_, connection_5__21__19_, connection_5__21__18_,
         connection_5__21__17_, connection_5__21__16_, connection_5__21__15_,
         connection_5__21__14_, connection_5__21__13_, connection_5__21__12_,
         connection_5__21__11_, connection_5__21__10_, connection_5__21__9_,
         connection_5__21__8_, connection_5__21__7_, connection_5__21__6_,
         connection_5__21__5_, connection_5__21__4_, connection_5__21__3_,
         connection_5__21__2_, connection_5__21__1_, connection_5__21__0_,
         connection_5__22__31_, connection_5__22__30_, connection_5__22__29_,
         connection_5__22__28_, connection_5__22__27_, connection_5__22__26_,
         connection_5__22__25_, connection_5__22__24_, connection_5__22__23_,
         connection_5__22__22_, connection_5__22__21_, connection_5__22__20_,
         connection_5__22__19_, connection_5__22__18_, connection_5__22__17_,
         connection_5__22__16_, connection_5__22__15_, connection_5__22__14_,
         connection_5__22__13_, connection_5__22__12_, connection_5__22__11_,
         connection_5__22__10_, connection_5__22__9_, connection_5__22__8_,
         connection_5__22__7_, connection_5__22__6_, connection_5__22__5_,
         connection_5__22__4_, connection_5__22__3_, connection_5__22__2_,
         connection_5__22__1_, connection_5__22__0_, connection_5__23__31_,
         connection_5__23__30_, connection_5__23__29_, connection_5__23__28_,
         connection_5__23__27_, connection_5__23__26_, connection_5__23__25_,
         connection_5__23__24_, connection_5__23__23_, connection_5__23__22_,
         connection_5__23__21_, connection_5__23__20_, connection_5__23__19_,
         connection_5__23__18_, connection_5__23__17_, connection_5__23__16_,
         connection_5__23__15_, connection_5__23__14_, connection_5__23__13_,
         connection_5__23__12_, connection_5__23__11_, connection_5__23__10_,
         connection_5__23__9_, connection_5__23__8_, connection_5__23__7_,
         connection_5__23__6_, connection_5__23__5_, connection_5__23__4_,
         connection_5__23__3_, connection_5__23__2_, connection_5__23__1_,
         connection_5__23__0_, connection_5__24__31_, connection_5__24__30_,
         connection_5__24__29_, connection_5__24__28_, connection_5__24__27_,
         connection_5__24__26_, connection_5__24__25_, connection_5__24__24_,
         connection_5__24__23_, connection_5__24__22_, connection_5__24__21_,
         connection_5__24__20_, connection_5__24__19_, connection_5__24__18_,
         connection_5__24__17_, connection_5__24__16_, connection_5__24__15_,
         connection_5__24__14_, connection_5__24__13_, connection_5__24__12_,
         connection_5__24__11_, connection_5__24__10_, connection_5__24__9_,
         connection_5__24__8_, connection_5__24__7_, connection_5__24__6_,
         connection_5__24__5_, connection_5__24__4_, connection_5__24__3_,
         connection_5__24__2_, connection_5__24__1_, connection_5__24__0_,
         connection_5__25__31_, connection_5__25__30_, connection_5__25__29_,
         connection_5__25__28_, connection_5__25__27_, connection_5__25__26_,
         connection_5__25__25_, connection_5__25__24_, connection_5__25__23_,
         connection_5__25__22_, connection_5__25__21_, connection_5__25__20_,
         connection_5__25__19_, connection_5__25__18_, connection_5__25__17_,
         connection_5__25__16_, connection_5__25__15_, connection_5__25__14_,
         connection_5__25__13_, connection_5__25__12_, connection_5__25__11_,
         connection_5__25__10_, connection_5__25__9_, connection_5__25__8_,
         connection_5__25__7_, connection_5__25__6_, connection_5__25__5_,
         connection_5__25__4_, connection_5__25__3_, connection_5__25__2_,
         connection_5__25__1_, connection_5__25__0_, connection_5__26__31_,
         connection_5__26__30_, connection_5__26__29_, connection_5__26__28_,
         connection_5__26__27_, connection_5__26__26_, connection_5__26__25_,
         connection_5__26__24_, connection_5__26__23_, connection_5__26__22_,
         connection_5__26__21_, connection_5__26__20_, connection_5__26__19_,
         connection_5__26__18_, connection_5__26__17_, connection_5__26__16_,
         connection_5__26__15_, connection_5__26__14_, connection_5__26__13_,
         connection_5__26__12_, connection_5__26__11_, connection_5__26__10_,
         connection_5__26__9_, connection_5__26__8_, connection_5__26__7_,
         connection_5__26__6_, connection_5__26__5_, connection_5__26__4_,
         connection_5__26__3_, connection_5__26__2_, connection_5__26__1_,
         connection_5__26__0_, connection_5__27__31_, connection_5__27__30_,
         connection_5__27__29_, connection_5__27__28_, connection_5__27__27_,
         connection_5__27__26_, connection_5__27__25_, connection_5__27__24_,
         connection_5__27__23_, connection_5__27__22_, connection_5__27__21_,
         connection_5__27__20_, connection_5__27__19_, connection_5__27__18_,
         connection_5__27__17_, connection_5__27__16_, connection_5__27__15_,
         connection_5__27__14_, connection_5__27__13_, connection_5__27__12_,
         connection_5__27__11_, connection_5__27__10_, connection_5__27__9_,
         connection_5__27__8_, connection_5__27__7_, connection_5__27__6_,
         connection_5__27__5_, connection_5__27__4_, connection_5__27__3_,
         connection_5__27__2_, connection_5__27__1_, connection_5__27__0_,
         connection_5__28__31_, connection_5__28__30_, connection_5__28__29_,
         connection_5__28__28_, connection_5__28__27_, connection_5__28__26_,
         connection_5__28__25_, connection_5__28__24_, connection_5__28__23_,
         connection_5__28__22_, connection_5__28__21_, connection_5__28__20_,
         connection_5__28__19_, connection_5__28__18_, connection_5__28__17_,
         connection_5__28__16_, connection_5__28__15_, connection_5__28__14_,
         connection_5__28__13_, connection_5__28__12_, connection_5__28__11_,
         connection_5__28__10_, connection_5__28__9_, connection_5__28__8_,
         connection_5__28__7_, connection_5__28__6_, connection_5__28__5_,
         connection_5__28__4_, connection_5__28__3_, connection_5__28__2_,
         connection_5__28__1_, connection_5__28__0_, connection_5__29__31_,
         connection_5__29__30_, connection_5__29__29_, connection_5__29__28_,
         connection_5__29__27_, connection_5__29__26_, connection_5__29__25_,
         connection_5__29__24_, connection_5__29__23_, connection_5__29__22_,
         connection_5__29__21_, connection_5__29__20_, connection_5__29__19_,
         connection_5__29__18_, connection_5__29__17_, connection_5__29__16_,
         connection_5__29__15_, connection_5__29__14_, connection_5__29__13_,
         connection_5__29__12_, connection_5__29__11_, connection_5__29__10_,
         connection_5__29__9_, connection_5__29__8_, connection_5__29__7_,
         connection_5__29__6_, connection_5__29__5_, connection_5__29__4_,
         connection_5__29__3_, connection_5__29__2_, connection_5__29__1_,
         connection_5__29__0_, connection_5__30__31_, connection_5__30__30_,
         connection_5__30__29_, connection_5__30__28_, connection_5__30__27_,
         connection_5__30__26_, connection_5__30__25_, connection_5__30__24_,
         connection_5__30__23_, connection_5__30__22_, connection_5__30__21_,
         connection_5__30__20_, connection_5__30__19_, connection_5__30__18_,
         connection_5__30__17_, connection_5__30__16_, connection_5__30__15_,
         connection_5__30__14_, connection_5__30__13_, connection_5__30__12_,
         connection_5__30__11_, connection_5__30__10_, connection_5__30__9_,
         connection_5__30__8_, connection_5__30__7_, connection_5__30__6_,
         connection_5__30__5_, connection_5__30__4_, connection_5__30__3_,
         connection_5__30__2_, connection_5__30__1_, connection_5__30__0_,
         connection_5__31__31_, connection_5__31__30_, connection_5__31__29_,
         connection_5__31__28_, connection_5__31__27_, connection_5__31__26_,
         connection_5__31__25_, connection_5__31__24_, connection_5__31__23_,
         connection_5__31__22_, connection_5__31__21_, connection_5__31__20_,
         connection_5__31__19_, connection_5__31__18_, connection_5__31__17_,
         connection_5__31__16_, connection_5__31__15_, connection_5__31__14_,
         connection_5__31__13_, connection_5__31__12_, connection_5__31__11_,
         connection_5__31__10_, connection_5__31__9_, connection_5__31__8_,
         connection_5__31__7_, connection_5__31__6_, connection_5__31__5_,
         connection_5__31__4_, connection_5__31__3_, connection_5__31__2_,
         connection_5__31__1_, connection_5__31__0_, connection_6__0__31_,
         connection_6__0__30_, connection_6__0__29_, connection_6__0__28_,
         connection_6__0__27_, connection_6__0__26_, connection_6__0__25_,
         connection_6__0__24_, connection_6__0__23_, connection_6__0__22_,
         connection_6__0__21_, connection_6__0__20_, connection_6__0__19_,
         connection_6__0__18_, connection_6__0__17_, connection_6__0__16_,
         connection_6__0__15_, connection_6__0__14_, connection_6__0__13_,
         connection_6__0__12_, connection_6__0__11_, connection_6__0__10_,
         connection_6__0__9_, connection_6__0__8_, connection_6__0__7_,
         connection_6__0__6_, connection_6__0__5_, connection_6__0__4_,
         connection_6__0__3_, connection_6__0__2_, connection_6__0__1_,
         connection_6__0__0_, connection_6__1__31_, connection_6__1__30_,
         connection_6__1__29_, connection_6__1__28_, connection_6__1__27_,
         connection_6__1__26_, connection_6__1__25_, connection_6__1__24_,
         connection_6__1__23_, connection_6__1__22_, connection_6__1__21_,
         connection_6__1__20_, connection_6__1__19_, connection_6__1__18_,
         connection_6__1__17_, connection_6__1__16_, connection_6__1__15_,
         connection_6__1__14_, connection_6__1__13_, connection_6__1__12_,
         connection_6__1__11_, connection_6__1__10_, connection_6__1__9_,
         connection_6__1__8_, connection_6__1__7_, connection_6__1__6_,
         connection_6__1__5_, connection_6__1__4_, connection_6__1__3_,
         connection_6__1__2_, connection_6__1__1_, connection_6__1__0_,
         connection_6__2__31_, connection_6__2__30_, connection_6__2__29_,
         connection_6__2__28_, connection_6__2__27_, connection_6__2__26_,
         connection_6__2__25_, connection_6__2__24_, connection_6__2__23_,
         connection_6__2__22_, connection_6__2__21_, connection_6__2__20_,
         connection_6__2__19_, connection_6__2__18_, connection_6__2__17_,
         connection_6__2__16_, connection_6__2__15_, connection_6__2__14_,
         connection_6__2__13_, connection_6__2__12_, connection_6__2__11_,
         connection_6__2__10_, connection_6__2__9_, connection_6__2__8_,
         connection_6__2__7_, connection_6__2__6_, connection_6__2__5_,
         connection_6__2__4_, connection_6__2__3_, connection_6__2__2_,
         connection_6__2__1_, connection_6__2__0_, connection_6__3__31_,
         connection_6__3__30_, connection_6__3__29_, connection_6__3__28_,
         connection_6__3__27_, connection_6__3__26_, connection_6__3__25_,
         connection_6__3__24_, connection_6__3__23_, connection_6__3__22_,
         connection_6__3__21_, connection_6__3__20_, connection_6__3__19_,
         connection_6__3__18_, connection_6__3__17_, connection_6__3__16_,
         connection_6__3__15_, connection_6__3__14_, connection_6__3__13_,
         connection_6__3__12_, connection_6__3__11_, connection_6__3__10_,
         connection_6__3__9_, connection_6__3__8_, connection_6__3__7_,
         connection_6__3__6_, connection_6__3__5_, connection_6__3__4_,
         connection_6__3__3_, connection_6__3__2_, connection_6__3__1_,
         connection_6__3__0_, connection_6__4__31_, connection_6__4__30_,
         connection_6__4__29_, connection_6__4__28_, connection_6__4__27_,
         connection_6__4__26_, connection_6__4__25_, connection_6__4__24_,
         connection_6__4__23_, connection_6__4__22_, connection_6__4__21_,
         connection_6__4__20_, connection_6__4__19_, connection_6__4__18_,
         connection_6__4__17_, connection_6__4__16_, connection_6__4__15_,
         connection_6__4__14_, connection_6__4__13_, connection_6__4__12_,
         connection_6__4__11_, connection_6__4__10_, connection_6__4__9_,
         connection_6__4__8_, connection_6__4__7_, connection_6__4__6_,
         connection_6__4__5_, connection_6__4__4_, connection_6__4__3_,
         connection_6__4__2_, connection_6__4__1_, connection_6__4__0_,
         connection_6__5__31_, connection_6__5__30_, connection_6__5__29_,
         connection_6__5__28_, connection_6__5__27_, connection_6__5__26_,
         connection_6__5__25_, connection_6__5__24_, connection_6__5__23_,
         connection_6__5__22_, connection_6__5__21_, connection_6__5__20_,
         connection_6__5__19_, connection_6__5__18_, connection_6__5__17_,
         connection_6__5__16_, connection_6__5__15_, connection_6__5__14_,
         connection_6__5__13_, connection_6__5__12_, connection_6__5__11_,
         connection_6__5__10_, connection_6__5__9_, connection_6__5__8_,
         connection_6__5__7_, connection_6__5__6_, connection_6__5__5_,
         connection_6__5__4_, connection_6__5__3_, connection_6__5__2_,
         connection_6__5__1_, connection_6__5__0_, connection_6__6__31_,
         connection_6__6__30_, connection_6__6__29_, connection_6__6__28_,
         connection_6__6__27_, connection_6__6__26_, connection_6__6__25_,
         connection_6__6__24_, connection_6__6__23_, connection_6__6__22_,
         connection_6__6__21_, connection_6__6__20_, connection_6__6__19_,
         connection_6__6__18_, connection_6__6__17_, connection_6__6__16_,
         connection_6__6__15_, connection_6__6__14_, connection_6__6__13_,
         connection_6__6__12_, connection_6__6__11_, connection_6__6__10_,
         connection_6__6__9_, connection_6__6__8_, connection_6__6__7_,
         connection_6__6__6_, connection_6__6__5_, connection_6__6__4_,
         connection_6__6__3_, connection_6__6__2_, connection_6__6__1_,
         connection_6__6__0_, connection_6__7__31_, connection_6__7__30_,
         connection_6__7__29_, connection_6__7__28_, connection_6__7__27_,
         connection_6__7__26_, connection_6__7__25_, connection_6__7__24_,
         connection_6__7__23_, connection_6__7__22_, connection_6__7__21_,
         connection_6__7__20_, connection_6__7__19_, connection_6__7__18_,
         connection_6__7__17_, connection_6__7__16_, connection_6__7__15_,
         connection_6__7__14_, connection_6__7__13_, connection_6__7__12_,
         connection_6__7__11_, connection_6__7__10_, connection_6__7__9_,
         connection_6__7__8_, connection_6__7__7_, connection_6__7__6_,
         connection_6__7__5_, connection_6__7__4_, connection_6__7__3_,
         connection_6__7__2_, connection_6__7__1_, connection_6__7__0_,
         connection_6__8__31_, connection_6__8__30_, connection_6__8__29_,
         connection_6__8__28_, connection_6__8__27_, connection_6__8__26_,
         connection_6__8__25_, connection_6__8__24_, connection_6__8__23_,
         connection_6__8__22_, connection_6__8__21_, connection_6__8__20_,
         connection_6__8__19_, connection_6__8__18_, connection_6__8__17_,
         connection_6__8__16_, connection_6__8__15_, connection_6__8__14_,
         connection_6__8__13_, connection_6__8__12_, connection_6__8__11_,
         connection_6__8__10_, connection_6__8__9_, connection_6__8__8_,
         connection_6__8__7_, connection_6__8__6_, connection_6__8__5_,
         connection_6__8__4_, connection_6__8__3_, connection_6__8__2_,
         connection_6__8__1_, connection_6__8__0_, connection_6__9__31_,
         connection_6__9__30_, connection_6__9__29_, connection_6__9__28_,
         connection_6__9__27_, connection_6__9__26_, connection_6__9__25_,
         connection_6__9__24_, connection_6__9__23_, connection_6__9__22_,
         connection_6__9__21_, connection_6__9__20_, connection_6__9__19_,
         connection_6__9__18_, connection_6__9__17_, connection_6__9__16_,
         connection_6__9__15_, connection_6__9__14_, connection_6__9__13_,
         connection_6__9__12_, connection_6__9__11_, connection_6__9__10_,
         connection_6__9__9_, connection_6__9__8_, connection_6__9__7_,
         connection_6__9__6_, connection_6__9__5_, connection_6__9__4_,
         connection_6__9__3_, connection_6__9__2_, connection_6__9__1_,
         connection_6__9__0_, connection_6__10__31_, connection_6__10__30_,
         connection_6__10__29_, connection_6__10__28_, connection_6__10__27_,
         connection_6__10__26_, connection_6__10__25_, connection_6__10__24_,
         connection_6__10__23_, connection_6__10__22_, connection_6__10__21_,
         connection_6__10__20_, connection_6__10__19_, connection_6__10__18_,
         connection_6__10__17_, connection_6__10__16_, connection_6__10__15_,
         connection_6__10__14_, connection_6__10__13_, connection_6__10__12_,
         connection_6__10__11_, connection_6__10__10_, connection_6__10__9_,
         connection_6__10__8_, connection_6__10__7_, connection_6__10__6_,
         connection_6__10__5_, connection_6__10__4_, connection_6__10__3_,
         connection_6__10__2_, connection_6__10__1_, connection_6__10__0_,
         connection_6__11__31_, connection_6__11__30_, connection_6__11__29_,
         connection_6__11__28_, connection_6__11__27_, connection_6__11__26_,
         connection_6__11__25_, connection_6__11__24_, connection_6__11__23_,
         connection_6__11__22_, connection_6__11__21_, connection_6__11__20_,
         connection_6__11__19_, connection_6__11__18_, connection_6__11__17_,
         connection_6__11__16_, connection_6__11__15_, connection_6__11__14_,
         connection_6__11__13_, connection_6__11__12_, connection_6__11__11_,
         connection_6__11__10_, connection_6__11__9_, connection_6__11__8_,
         connection_6__11__7_, connection_6__11__6_, connection_6__11__5_,
         connection_6__11__4_, connection_6__11__3_, connection_6__11__2_,
         connection_6__11__1_, connection_6__11__0_, connection_6__12__31_,
         connection_6__12__30_, connection_6__12__29_, connection_6__12__28_,
         connection_6__12__27_, connection_6__12__26_, connection_6__12__25_,
         connection_6__12__24_, connection_6__12__23_, connection_6__12__22_,
         connection_6__12__21_, connection_6__12__20_, connection_6__12__19_,
         connection_6__12__18_, connection_6__12__17_, connection_6__12__16_,
         connection_6__12__15_, connection_6__12__14_, connection_6__12__13_,
         connection_6__12__12_, connection_6__12__11_, connection_6__12__10_,
         connection_6__12__9_, connection_6__12__8_, connection_6__12__7_,
         connection_6__12__6_, connection_6__12__5_, connection_6__12__4_,
         connection_6__12__3_, connection_6__12__2_, connection_6__12__1_,
         connection_6__12__0_, connection_6__13__31_, connection_6__13__30_,
         connection_6__13__29_, connection_6__13__28_, connection_6__13__27_,
         connection_6__13__26_, connection_6__13__25_, connection_6__13__24_,
         connection_6__13__23_, connection_6__13__22_, connection_6__13__21_,
         connection_6__13__20_, connection_6__13__19_, connection_6__13__18_,
         connection_6__13__17_, connection_6__13__16_, connection_6__13__15_,
         connection_6__13__14_, connection_6__13__13_, connection_6__13__12_,
         connection_6__13__11_, connection_6__13__10_, connection_6__13__9_,
         connection_6__13__8_, connection_6__13__7_, connection_6__13__6_,
         connection_6__13__5_, connection_6__13__4_, connection_6__13__3_,
         connection_6__13__2_, connection_6__13__1_, connection_6__13__0_,
         connection_6__14__31_, connection_6__14__30_, connection_6__14__29_,
         connection_6__14__28_, connection_6__14__27_, connection_6__14__26_,
         connection_6__14__25_, connection_6__14__24_, connection_6__14__23_,
         connection_6__14__22_, connection_6__14__21_, connection_6__14__20_,
         connection_6__14__19_, connection_6__14__18_, connection_6__14__17_,
         connection_6__14__16_, connection_6__14__15_, connection_6__14__14_,
         connection_6__14__13_, connection_6__14__12_, connection_6__14__11_,
         connection_6__14__10_, connection_6__14__9_, connection_6__14__8_,
         connection_6__14__7_, connection_6__14__6_, connection_6__14__5_,
         connection_6__14__4_, connection_6__14__3_, connection_6__14__2_,
         connection_6__14__1_, connection_6__14__0_, connection_6__15__31_,
         connection_6__15__30_, connection_6__15__29_, connection_6__15__28_,
         connection_6__15__27_, connection_6__15__26_, connection_6__15__25_,
         connection_6__15__24_, connection_6__15__23_, connection_6__15__22_,
         connection_6__15__21_, connection_6__15__20_, connection_6__15__19_,
         connection_6__15__18_, connection_6__15__17_, connection_6__15__16_,
         connection_6__15__15_, connection_6__15__14_, connection_6__15__13_,
         connection_6__15__12_, connection_6__15__11_, connection_6__15__10_,
         connection_6__15__9_, connection_6__15__8_, connection_6__15__7_,
         connection_6__15__6_, connection_6__15__5_, connection_6__15__4_,
         connection_6__15__3_, connection_6__15__2_, connection_6__15__1_,
         connection_6__15__0_, connection_6__16__31_, connection_6__16__30_,
         connection_6__16__29_, connection_6__16__28_, connection_6__16__27_,
         connection_6__16__26_, connection_6__16__25_, connection_6__16__24_,
         connection_6__16__23_, connection_6__16__22_, connection_6__16__21_,
         connection_6__16__20_, connection_6__16__19_, connection_6__16__18_,
         connection_6__16__17_, connection_6__16__16_, connection_6__16__15_,
         connection_6__16__14_, connection_6__16__13_, connection_6__16__12_,
         connection_6__16__11_, connection_6__16__10_, connection_6__16__9_,
         connection_6__16__8_, connection_6__16__7_, connection_6__16__6_,
         connection_6__16__5_, connection_6__16__4_, connection_6__16__3_,
         connection_6__16__2_, connection_6__16__1_, connection_6__16__0_,
         connection_6__17__31_, connection_6__17__30_, connection_6__17__29_,
         connection_6__17__28_, connection_6__17__27_, connection_6__17__26_,
         connection_6__17__25_, connection_6__17__24_, connection_6__17__23_,
         connection_6__17__22_, connection_6__17__21_, connection_6__17__20_,
         connection_6__17__19_, connection_6__17__18_, connection_6__17__17_,
         connection_6__17__16_, connection_6__17__15_, connection_6__17__14_,
         connection_6__17__13_, connection_6__17__12_, connection_6__17__11_,
         connection_6__17__10_, connection_6__17__9_, connection_6__17__8_,
         connection_6__17__7_, connection_6__17__6_, connection_6__17__5_,
         connection_6__17__4_, connection_6__17__3_, connection_6__17__2_,
         connection_6__17__1_, connection_6__17__0_, connection_6__18__31_,
         connection_6__18__30_, connection_6__18__29_, connection_6__18__28_,
         connection_6__18__27_, connection_6__18__26_, connection_6__18__25_,
         connection_6__18__24_, connection_6__18__23_, connection_6__18__22_,
         connection_6__18__21_, connection_6__18__20_, connection_6__18__19_,
         connection_6__18__18_, connection_6__18__17_, connection_6__18__16_,
         connection_6__18__15_, connection_6__18__14_, connection_6__18__13_,
         connection_6__18__12_, connection_6__18__11_, connection_6__18__10_,
         connection_6__18__9_, connection_6__18__8_, connection_6__18__7_,
         connection_6__18__6_, connection_6__18__5_, connection_6__18__4_,
         connection_6__18__3_, connection_6__18__2_, connection_6__18__1_,
         connection_6__18__0_, connection_6__19__31_, connection_6__19__30_,
         connection_6__19__29_, connection_6__19__28_, connection_6__19__27_,
         connection_6__19__26_, connection_6__19__25_, connection_6__19__24_,
         connection_6__19__23_, connection_6__19__22_, connection_6__19__21_,
         connection_6__19__20_, connection_6__19__19_, connection_6__19__18_,
         connection_6__19__17_, connection_6__19__16_, connection_6__19__15_,
         connection_6__19__14_, connection_6__19__13_, connection_6__19__12_,
         connection_6__19__11_, connection_6__19__10_, connection_6__19__9_,
         connection_6__19__8_, connection_6__19__7_, connection_6__19__6_,
         connection_6__19__5_, connection_6__19__4_, connection_6__19__3_,
         connection_6__19__2_, connection_6__19__1_, connection_6__19__0_,
         connection_6__20__31_, connection_6__20__30_, connection_6__20__29_,
         connection_6__20__28_, connection_6__20__27_, connection_6__20__26_,
         connection_6__20__25_, connection_6__20__24_, connection_6__20__23_,
         connection_6__20__22_, connection_6__20__21_, connection_6__20__20_,
         connection_6__20__19_, connection_6__20__18_, connection_6__20__17_,
         connection_6__20__16_, connection_6__20__15_, connection_6__20__14_,
         connection_6__20__13_, connection_6__20__12_, connection_6__20__11_,
         connection_6__20__10_, connection_6__20__9_, connection_6__20__8_,
         connection_6__20__7_, connection_6__20__6_, connection_6__20__5_,
         connection_6__20__4_, connection_6__20__3_, connection_6__20__2_,
         connection_6__20__1_, connection_6__20__0_, connection_6__21__31_,
         connection_6__21__30_, connection_6__21__29_, connection_6__21__28_,
         connection_6__21__27_, connection_6__21__26_, connection_6__21__25_,
         connection_6__21__24_, connection_6__21__23_, connection_6__21__22_,
         connection_6__21__21_, connection_6__21__20_, connection_6__21__19_,
         connection_6__21__18_, connection_6__21__17_, connection_6__21__16_,
         connection_6__21__15_, connection_6__21__14_, connection_6__21__13_,
         connection_6__21__12_, connection_6__21__11_, connection_6__21__10_,
         connection_6__21__9_, connection_6__21__8_, connection_6__21__7_,
         connection_6__21__6_, connection_6__21__5_, connection_6__21__4_,
         connection_6__21__3_, connection_6__21__2_, connection_6__21__1_,
         connection_6__21__0_, connection_6__22__31_, connection_6__22__30_,
         connection_6__22__29_, connection_6__22__28_, connection_6__22__27_,
         connection_6__22__26_, connection_6__22__25_, connection_6__22__24_,
         connection_6__22__23_, connection_6__22__22_, connection_6__22__21_,
         connection_6__22__20_, connection_6__22__19_, connection_6__22__18_,
         connection_6__22__17_, connection_6__22__16_, connection_6__22__15_,
         connection_6__22__14_, connection_6__22__13_, connection_6__22__12_,
         connection_6__22__11_, connection_6__22__10_, connection_6__22__9_,
         connection_6__22__8_, connection_6__22__7_, connection_6__22__6_,
         connection_6__22__5_, connection_6__22__4_, connection_6__22__3_,
         connection_6__22__2_, connection_6__22__1_, connection_6__22__0_,
         connection_6__23__31_, connection_6__23__30_, connection_6__23__29_,
         connection_6__23__28_, connection_6__23__27_, connection_6__23__26_,
         connection_6__23__25_, connection_6__23__24_, connection_6__23__23_,
         connection_6__23__22_, connection_6__23__21_, connection_6__23__20_,
         connection_6__23__19_, connection_6__23__18_, connection_6__23__17_,
         connection_6__23__16_, connection_6__23__15_, connection_6__23__14_,
         connection_6__23__13_, connection_6__23__12_, connection_6__23__11_,
         connection_6__23__10_, connection_6__23__9_, connection_6__23__8_,
         connection_6__23__7_, connection_6__23__6_, connection_6__23__5_,
         connection_6__23__4_, connection_6__23__3_, connection_6__23__2_,
         connection_6__23__1_, connection_6__23__0_, connection_6__24__31_,
         connection_6__24__30_, connection_6__24__29_, connection_6__24__28_,
         connection_6__24__27_, connection_6__24__26_, connection_6__24__25_,
         connection_6__24__24_, connection_6__24__23_, connection_6__24__22_,
         connection_6__24__21_, connection_6__24__20_, connection_6__24__19_,
         connection_6__24__18_, connection_6__24__17_, connection_6__24__16_,
         connection_6__24__15_, connection_6__24__14_, connection_6__24__13_,
         connection_6__24__12_, connection_6__24__11_, connection_6__24__10_,
         connection_6__24__9_, connection_6__24__8_, connection_6__24__7_,
         connection_6__24__6_, connection_6__24__5_, connection_6__24__4_,
         connection_6__24__3_, connection_6__24__2_, connection_6__24__1_,
         connection_6__24__0_, connection_6__25__31_, connection_6__25__30_,
         connection_6__25__29_, connection_6__25__28_, connection_6__25__27_,
         connection_6__25__26_, connection_6__25__25_, connection_6__25__24_,
         connection_6__25__23_, connection_6__25__22_, connection_6__25__21_,
         connection_6__25__20_, connection_6__25__19_, connection_6__25__18_,
         connection_6__25__17_, connection_6__25__16_, connection_6__25__15_,
         connection_6__25__14_, connection_6__25__13_, connection_6__25__12_,
         connection_6__25__11_, connection_6__25__10_, connection_6__25__9_,
         connection_6__25__8_, connection_6__25__7_, connection_6__25__6_,
         connection_6__25__5_, connection_6__25__4_, connection_6__25__3_,
         connection_6__25__2_, connection_6__25__1_, connection_6__25__0_,
         connection_6__26__31_, connection_6__26__30_, connection_6__26__29_,
         connection_6__26__28_, connection_6__26__27_, connection_6__26__26_,
         connection_6__26__25_, connection_6__26__24_, connection_6__26__23_,
         connection_6__26__22_, connection_6__26__21_, connection_6__26__20_,
         connection_6__26__19_, connection_6__26__18_, connection_6__26__17_,
         connection_6__26__16_, connection_6__26__15_, connection_6__26__14_,
         connection_6__26__13_, connection_6__26__12_, connection_6__26__11_,
         connection_6__26__10_, connection_6__26__9_, connection_6__26__8_,
         connection_6__26__7_, connection_6__26__6_, connection_6__26__5_,
         connection_6__26__4_, connection_6__26__3_, connection_6__26__2_,
         connection_6__26__1_, connection_6__26__0_, connection_6__27__31_,
         connection_6__27__30_, connection_6__27__29_, connection_6__27__28_,
         connection_6__27__27_, connection_6__27__26_, connection_6__27__25_,
         connection_6__27__24_, connection_6__27__23_, connection_6__27__22_,
         connection_6__27__21_, connection_6__27__20_, connection_6__27__19_,
         connection_6__27__18_, connection_6__27__17_, connection_6__27__16_,
         connection_6__27__15_, connection_6__27__14_, connection_6__27__13_,
         connection_6__27__12_, connection_6__27__11_, connection_6__27__10_,
         connection_6__27__9_, connection_6__27__8_, connection_6__27__7_,
         connection_6__27__6_, connection_6__27__5_, connection_6__27__4_,
         connection_6__27__3_, connection_6__27__2_, connection_6__27__1_,
         connection_6__27__0_, connection_6__28__31_, connection_6__28__30_,
         connection_6__28__29_, connection_6__28__28_, connection_6__28__27_,
         connection_6__28__26_, connection_6__28__25_, connection_6__28__24_,
         connection_6__28__23_, connection_6__28__22_, connection_6__28__21_,
         connection_6__28__20_, connection_6__28__19_, connection_6__28__18_,
         connection_6__28__17_, connection_6__28__16_, connection_6__28__15_,
         connection_6__28__14_, connection_6__28__13_, connection_6__28__12_,
         connection_6__28__11_, connection_6__28__10_, connection_6__28__9_,
         connection_6__28__8_, connection_6__28__7_, connection_6__28__6_,
         connection_6__28__5_, connection_6__28__4_, connection_6__28__3_,
         connection_6__28__2_, connection_6__28__1_, connection_6__28__0_,
         connection_6__29__31_, connection_6__29__30_, connection_6__29__29_,
         connection_6__29__28_, connection_6__29__27_, connection_6__29__26_,
         connection_6__29__25_, connection_6__29__24_, connection_6__29__23_,
         connection_6__29__22_, connection_6__29__21_, connection_6__29__20_,
         connection_6__29__19_, connection_6__29__18_, connection_6__29__17_,
         connection_6__29__16_, connection_6__29__15_, connection_6__29__14_,
         connection_6__29__13_, connection_6__29__12_, connection_6__29__11_,
         connection_6__29__10_, connection_6__29__9_, connection_6__29__8_,
         connection_6__29__7_, connection_6__29__6_, connection_6__29__5_,
         connection_6__29__4_, connection_6__29__3_, connection_6__29__2_,
         connection_6__29__1_, connection_6__29__0_, connection_6__30__31_,
         connection_6__30__30_, connection_6__30__29_, connection_6__30__28_,
         connection_6__30__27_, connection_6__30__26_, connection_6__30__25_,
         connection_6__30__24_, connection_6__30__23_, connection_6__30__22_,
         connection_6__30__21_, connection_6__30__20_, connection_6__30__19_,
         connection_6__30__18_, connection_6__30__17_, connection_6__30__16_,
         connection_6__30__15_, connection_6__30__14_, connection_6__30__13_,
         connection_6__30__12_, connection_6__30__11_, connection_6__30__10_,
         connection_6__30__9_, connection_6__30__8_, connection_6__30__7_,
         connection_6__30__6_, connection_6__30__5_, connection_6__30__4_,
         connection_6__30__3_, connection_6__30__2_, connection_6__30__1_,
         connection_6__30__0_, connection_6__31__31_, connection_6__31__30_,
         connection_6__31__29_, connection_6__31__28_, connection_6__31__27_,
         connection_6__31__26_, connection_6__31__25_, connection_6__31__24_,
         connection_6__31__23_, connection_6__31__22_, connection_6__31__21_,
         connection_6__31__20_, connection_6__31__19_, connection_6__31__18_,
         connection_6__31__17_, connection_6__31__16_, connection_6__31__15_,
         connection_6__31__14_, connection_6__31__13_, connection_6__31__12_,
         connection_6__31__11_, connection_6__31__10_, connection_6__31__9_,
         connection_6__31__8_, connection_6__31__7_, connection_6__31__6_,
         connection_6__31__5_, connection_6__31__4_, connection_6__31__3_,
         connection_6__31__2_, connection_6__31__1_, connection_6__31__0_,
         connection_7__0__31_, connection_7__0__30_, connection_7__0__29_,
         connection_7__0__28_, connection_7__0__27_, connection_7__0__26_,
         connection_7__0__25_, connection_7__0__24_, connection_7__0__23_,
         connection_7__0__22_, connection_7__0__21_, connection_7__0__20_,
         connection_7__0__19_, connection_7__0__18_, connection_7__0__17_,
         connection_7__0__16_, connection_7__0__15_, connection_7__0__14_,
         connection_7__0__13_, connection_7__0__12_, connection_7__0__11_,
         connection_7__0__10_, connection_7__0__9_, connection_7__0__8_,
         connection_7__0__7_, connection_7__0__6_, connection_7__0__5_,
         connection_7__0__4_, connection_7__0__3_, connection_7__0__2_,
         connection_7__0__1_, connection_7__0__0_, connection_7__1__31_,
         connection_7__1__30_, connection_7__1__29_, connection_7__1__28_,
         connection_7__1__27_, connection_7__1__26_, connection_7__1__25_,
         connection_7__1__24_, connection_7__1__23_, connection_7__1__22_,
         connection_7__1__21_, connection_7__1__20_, connection_7__1__19_,
         connection_7__1__18_, connection_7__1__17_, connection_7__1__16_,
         connection_7__1__15_, connection_7__1__14_, connection_7__1__13_,
         connection_7__1__12_, connection_7__1__11_, connection_7__1__10_,
         connection_7__1__9_, connection_7__1__8_, connection_7__1__7_,
         connection_7__1__6_, connection_7__1__5_, connection_7__1__4_,
         connection_7__1__3_, connection_7__1__2_, connection_7__1__1_,
         connection_7__1__0_, connection_7__2__31_, connection_7__2__30_,
         connection_7__2__29_, connection_7__2__28_, connection_7__2__27_,
         connection_7__2__26_, connection_7__2__25_, connection_7__2__24_,
         connection_7__2__23_, connection_7__2__22_, connection_7__2__21_,
         connection_7__2__20_, connection_7__2__19_, connection_7__2__18_,
         connection_7__2__17_, connection_7__2__16_, connection_7__2__15_,
         connection_7__2__14_, connection_7__2__13_, connection_7__2__12_,
         connection_7__2__11_, connection_7__2__10_, connection_7__2__9_,
         connection_7__2__8_, connection_7__2__7_, connection_7__2__6_,
         connection_7__2__5_, connection_7__2__4_, connection_7__2__3_,
         connection_7__2__2_, connection_7__2__1_, connection_7__2__0_,
         connection_7__3__31_, connection_7__3__30_, connection_7__3__29_,
         connection_7__3__28_, connection_7__3__27_, connection_7__3__26_,
         connection_7__3__25_, connection_7__3__24_, connection_7__3__23_,
         connection_7__3__22_, connection_7__3__21_, connection_7__3__20_,
         connection_7__3__19_, connection_7__3__18_, connection_7__3__17_,
         connection_7__3__16_, connection_7__3__15_, connection_7__3__14_,
         connection_7__3__13_, connection_7__3__12_, connection_7__3__11_,
         connection_7__3__10_, connection_7__3__9_, connection_7__3__8_,
         connection_7__3__7_, connection_7__3__6_, connection_7__3__5_,
         connection_7__3__4_, connection_7__3__3_, connection_7__3__2_,
         connection_7__3__1_, connection_7__3__0_, connection_7__4__31_,
         connection_7__4__30_, connection_7__4__29_, connection_7__4__28_,
         connection_7__4__27_, connection_7__4__26_, connection_7__4__25_,
         connection_7__4__24_, connection_7__4__23_, connection_7__4__22_,
         connection_7__4__21_, connection_7__4__20_, connection_7__4__19_,
         connection_7__4__18_, connection_7__4__17_, connection_7__4__16_,
         connection_7__4__15_, connection_7__4__14_, connection_7__4__13_,
         connection_7__4__12_, connection_7__4__11_, connection_7__4__10_,
         connection_7__4__9_, connection_7__4__8_, connection_7__4__7_,
         connection_7__4__6_, connection_7__4__5_, connection_7__4__4_,
         connection_7__4__3_, connection_7__4__2_, connection_7__4__1_,
         connection_7__4__0_, connection_7__5__31_, connection_7__5__30_,
         connection_7__5__29_, connection_7__5__28_, connection_7__5__27_,
         connection_7__5__26_, connection_7__5__25_, connection_7__5__24_,
         connection_7__5__23_, connection_7__5__22_, connection_7__5__21_,
         connection_7__5__20_, connection_7__5__19_, connection_7__5__18_,
         connection_7__5__17_, connection_7__5__16_, connection_7__5__15_,
         connection_7__5__14_, connection_7__5__13_, connection_7__5__12_,
         connection_7__5__11_, connection_7__5__10_, connection_7__5__9_,
         connection_7__5__8_, connection_7__5__7_, connection_7__5__6_,
         connection_7__5__5_, connection_7__5__4_, connection_7__5__3_,
         connection_7__5__2_, connection_7__5__1_, connection_7__5__0_,
         connection_7__6__31_, connection_7__6__30_, connection_7__6__29_,
         connection_7__6__28_, connection_7__6__27_, connection_7__6__26_,
         connection_7__6__25_, connection_7__6__24_, connection_7__6__23_,
         connection_7__6__22_, connection_7__6__21_, connection_7__6__20_,
         connection_7__6__19_, connection_7__6__18_, connection_7__6__17_,
         connection_7__6__16_, connection_7__6__15_, connection_7__6__14_,
         connection_7__6__13_, connection_7__6__12_, connection_7__6__11_,
         connection_7__6__10_, connection_7__6__9_, connection_7__6__8_,
         connection_7__6__7_, connection_7__6__6_, connection_7__6__5_,
         connection_7__6__4_, connection_7__6__3_, connection_7__6__2_,
         connection_7__6__1_, connection_7__6__0_, connection_7__7__31_,
         connection_7__7__30_, connection_7__7__29_, connection_7__7__28_,
         connection_7__7__27_, connection_7__7__26_, connection_7__7__25_,
         connection_7__7__24_, connection_7__7__23_, connection_7__7__22_,
         connection_7__7__21_, connection_7__7__20_, connection_7__7__19_,
         connection_7__7__18_, connection_7__7__17_, connection_7__7__16_,
         connection_7__7__15_, connection_7__7__14_, connection_7__7__13_,
         connection_7__7__12_, connection_7__7__11_, connection_7__7__10_,
         connection_7__7__9_, connection_7__7__8_, connection_7__7__7_,
         connection_7__7__6_, connection_7__7__5_, connection_7__7__4_,
         connection_7__7__3_, connection_7__7__2_, connection_7__7__1_,
         connection_7__7__0_, connection_7__8__31_, connection_7__8__30_,
         connection_7__8__29_, connection_7__8__28_, connection_7__8__27_,
         connection_7__8__26_, connection_7__8__25_, connection_7__8__24_,
         connection_7__8__23_, connection_7__8__22_, connection_7__8__21_,
         connection_7__8__20_, connection_7__8__19_, connection_7__8__18_,
         connection_7__8__17_, connection_7__8__16_, connection_7__8__15_,
         connection_7__8__14_, connection_7__8__13_, connection_7__8__12_,
         connection_7__8__11_, connection_7__8__10_, connection_7__8__9_,
         connection_7__8__8_, connection_7__8__7_, connection_7__8__6_,
         connection_7__8__5_, connection_7__8__4_, connection_7__8__3_,
         connection_7__8__2_, connection_7__8__1_, connection_7__8__0_,
         connection_7__9__31_, connection_7__9__30_, connection_7__9__29_,
         connection_7__9__28_, connection_7__9__27_, connection_7__9__26_,
         connection_7__9__25_, connection_7__9__24_, connection_7__9__23_,
         connection_7__9__22_, connection_7__9__21_, connection_7__9__20_,
         connection_7__9__19_, connection_7__9__18_, connection_7__9__17_,
         connection_7__9__16_, connection_7__9__15_, connection_7__9__14_,
         connection_7__9__13_, connection_7__9__12_, connection_7__9__11_,
         connection_7__9__10_, connection_7__9__9_, connection_7__9__8_,
         connection_7__9__7_, connection_7__9__6_, connection_7__9__5_,
         connection_7__9__4_, connection_7__9__3_, connection_7__9__2_,
         connection_7__9__1_, connection_7__9__0_, connection_7__10__31_,
         connection_7__10__30_, connection_7__10__29_, connection_7__10__28_,
         connection_7__10__27_, connection_7__10__26_, connection_7__10__25_,
         connection_7__10__24_, connection_7__10__23_, connection_7__10__22_,
         connection_7__10__21_, connection_7__10__20_, connection_7__10__19_,
         connection_7__10__18_, connection_7__10__17_, connection_7__10__16_,
         connection_7__10__15_, connection_7__10__14_, connection_7__10__13_,
         connection_7__10__12_, connection_7__10__11_, connection_7__10__10_,
         connection_7__10__9_, connection_7__10__8_, connection_7__10__7_,
         connection_7__10__6_, connection_7__10__5_, connection_7__10__4_,
         connection_7__10__3_, connection_7__10__2_, connection_7__10__1_,
         connection_7__10__0_, connection_7__11__31_, connection_7__11__30_,
         connection_7__11__29_, connection_7__11__28_, connection_7__11__27_,
         connection_7__11__26_, connection_7__11__25_, connection_7__11__24_,
         connection_7__11__23_, connection_7__11__22_, connection_7__11__21_,
         connection_7__11__20_, connection_7__11__19_, connection_7__11__18_,
         connection_7__11__17_, connection_7__11__16_, connection_7__11__15_,
         connection_7__11__14_, connection_7__11__13_, connection_7__11__12_,
         connection_7__11__11_, connection_7__11__10_, connection_7__11__9_,
         connection_7__11__8_, connection_7__11__7_, connection_7__11__6_,
         connection_7__11__5_, connection_7__11__4_, connection_7__11__3_,
         connection_7__11__2_, connection_7__11__1_, connection_7__11__0_,
         connection_7__12__31_, connection_7__12__30_, connection_7__12__29_,
         connection_7__12__28_, connection_7__12__27_, connection_7__12__26_,
         connection_7__12__25_, connection_7__12__24_, connection_7__12__23_,
         connection_7__12__22_, connection_7__12__21_, connection_7__12__20_,
         connection_7__12__19_, connection_7__12__18_, connection_7__12__17_,
         connection_7__12__16_, connection_7__12__15_, connection_7__12__14_,
         connection_7__12__13_, connection_7__12__12_, connection_7__12__11_,
         connection_7__12__10_, connection_7__12__9_, connection_7__12__8_,
         connection_7__12__7_, connection_7__12__6_, connection_7__12__5_,
         connection_7__12__4_, connection_7__12__3_, connection_7__12__2_,
         connection_7__12__1_, connection_7__12__0_, connection_7__13__31_,
         connection_7__13__30_, connection_7__13__29_, connection_7__13__28_,
         connection_7__13__27_, connection_7__13__26_, connection_7__13__25_,
         connection_7__13__24_, connection_7__13__23_, connection_7__13__22_,
         connection_7__13__21_, connection_7__13__20_, connection_7__13__19_,
         connection_7__13__18_, connection_7__13__17_, connection_7__13__16_,
         connection_7__13__15_, connection_7__13__14_, connection_7__13__13_,
         connection_7__13__12_, connection_7__13__11_, connection_7__13__10_,
         connection_7__13__9_, connection_7__13__8_, connection_7__13__7_,
         connection_7__13__6_, connection_7__13__5_, connection_7__13__4_,
         connection_7__13__3_, connection_7__13__2_, connection_7__13__1_,
         connection_7__13__0_, connection_7__14__31_, connection_7__14__30_,
         connection_7__14__29_, connection_7__14__28_, connection_7__14__27_,
         connection_7__14__26_, connection_7__14__25_, connection_7__14__24_,
         connection_7__14__23_, connection_7__14__22_, connection_7__14__21_,
         connection_7__14__20_, connection_7__14__19_, connection_7__14__18_,
         connection_7__14__17_, connection_7__14__16_, connection_7__14__15_,
         connection_7__14__14_, connection_7__14__13_, connection_7__14__12_,
         connection_7__14__11_, connection_7__14__10_, connection_7__14__9_,
         connection_7__14__8_, connection_7__14__7_, connection_7__14__6_,
         connection_7__14__5_, connection_7__14__4_, connection_7__14__3_,
         connection_7__14__2_, connection_7__14__1_, connection_7__14__0_,
         connection_7__15__31_, connection_7__15__30_, connection_7__15__29_,
         connection_7__15__28_, connection_7__15__27_, connection_7__15__26_,
         connection_7__15__25_, connection_7__15__24_, connection_7__15__23_,
         connection_7__15__22_, connection_7__15__21_, connection_7__15__20_,
         connection_7__15__19_, connection_7__15__18_, connection_7__15__17_,
         connection_7__15__16_, connection_7__15__15_, connection_7__15__14_,
         connection_7__15__13_, connection_7__15__12_, connection_7__15__11_,
         connection_7__15__10_, connection_7__15__9_, connection_7__15__8_,
         connection_7__15__7_, connection_7__15__6_, connection_7__15__5_,
         connection_7__15__4_, connection_7__15__3_, connection_7__15__2_,
         connection_7__15__1_, connection_7__15__0_, connection_7__16__31_,
         connection_7__16__30_, connection_7__16__29_, connection_7__16__28_,
         connection_7__16__27_, connection_7__16__26_, connection_7__16__25_,
         connection_7__16__24_, connection_7__16__23_, connection_7__16__22_,
         connection_7__16__21_, connection_7__16__20_, connection_7__16__19_,
         connection_7__16__18_, connection_7__16__17_, connection_7__16__16_,
         connection_7__16__15_, connection_7__16__14_, connection_7__16__13_,
         connection_7__16__12_, connection_7__16__11_, connection_7__16__10_,
         connection_7__16__9_, connection_7__16__8_, connection_7__16__7_,
         connection_7__16__6_, connection_7__16__5_, connection_7__16__4_,
         connection_7__16__3_, connection_7__16__2_, connection_7__16__1_,
         connection_7__16__0_, connection_7__17__31_, connection_7__17__30_,
         connection_7__17__29_, connection_7__17__28_, connection_7__17__27_,
         connection_7__17__26_, connection_7__17__25_, connection_7__17__24_,
         connection_7__17__23_, connection_7__17__22_, connection_7__17__21_,
         connection_7__17__20_, connection_7__17__19_, connection_7__17__18_,
         connection_7__17__17_, connection_7__17__16_, connection_7__17__15_,
         connection_7__17__14_, connection_7__17__13_, connection_7__17__12_,
         connection_7__17__11_, connection_7__17__10_, connection_7__17__9_,
         connection_7__17__8_, connection_7__17__7_, connection_7__17__6_,
         connection_7__17__5_, connection_7__17__4_, connection_7__17__3_,
         connection_7__17__2_, connection_7__17__1_, connection_7__17__0_,
         connection_7__18__31_, connection_7__18__30_, connection_7__18__29_,
         connection_7__18__28_, connection_7__18__27_, connection_7__18__26_,
         connection_7__18__25_, connection_7__18__24_, connection_7__18__23_,
         connection_7__18__22_, connection_7__18__21_, connection_7__18__20_,
         connection_7__18__19_, connection_7__18__18_, connection_7__18__17_,
         connection_7__18__16_, connection_7__18__15_, connection_7__18__14_,
         connection_7__18__13_, connection_7__18__12_, connection_7__18__11_,
         connection_7__18__10_, connection_7__18__9_, connection_7__18__8_,
         connection_7__18__7_, connection_7__18__6_, connection_7__18__5_,
         connection_7__18__4_, connection_7__18__3_, connection_7__18__2_,
         connection_7__18__1_, connection_7__18__0_, connection_7__19__31_,
         connection_7__19__30_, connection_7__19__29_, connection_7__19__28_,
         connection_7__19__27_, connection_7__19__26_, connection_7__19__25_,
         connection_7__19__24_, connection_7__19__23_, connection_7__19__22_,
         connection_7__19__21_, connection_7__19__20_, connection_7__19__19_,
         connection_7__19__18_, connection_7__19__17_, connection_7__19__16_,
         connection_7__19__15_, connection_7__19__14_, connection_7__19__13_,
         connection_7__19__12_, connection_7__19__11_, connection_7__19__10_,
         connection_7__19__9_, connection_7__19__8_, connection_7__19__7_,
         connection_7__19__6_, connection_7__19__5_, connection_7__19__4_,
         connection_7__19__3_, connection_7__19__2_, connection_7__19__1_,
         connection_7__19__0_, connection_7__20__31_, connection_7__20__30_,
         connection_7__20__29_, connection_7__20__28_, connection_7__20__27_,
         connection_7__20__26_, connection_7__20__25_, connection_7__20__24_,
         connection_7__20__23_, connection_7__20__22_, connection_7__20__21_,
         connection_7__20__20_, connection_7__20__19_, connection_7__20__18_,
         connection_7__20__17_, connection_7__20__16_, connection_7__20__15_,
         connection_7__20__14_, connection_7__20__13_, connection_7__20__12_,
         connection_7__20__11_, connection_7__20__10_, connection_7__20__9_,
         connection_7__20__8_, connection_7__20__7_, connection_7__20__6_,
         connection_7__20__5_, connection_7__20__4_, connection_7__20__3_,
         connection_7__20__2_, connection_7__20__1_, connection_7__20__0_,
         connection_7__21__31_, connection_7__21__30_, connection_7__21__29_,
         connection_7__21__28_, connection_7__21__27_, connection_7__21__26_,
         connection_7__21__25_, connection_7__21__24_, connection_7__21__23_,
         connection_7__21__22_, connection_7__21__21_, connection_7__21__20_,
         connection_7__21__19_, connection_7__21__18_, connection_7__21__17_,
         connection_7__21__16_, connection_7__21__15_, connection_7__21__14_,
         connection_7__21__13_, connection_7__21__12_, connection_7__21__11_,
         connection_7__21__10_, connection_7__21__9_, connection_7__21__8_,
         connection_7__21__7_, connection_7__21__6_, connection_7__21__5_,
         connection_7__21__4_, connection_7__21__3_, connection_7__21__2_,
         connection_7__21__1_, connection_7__21__0_, connection_7__22__31_,
         connection_7__22__30_, connection_7__22__29_, connection_7__22__28_,
         connection_7__22__27_, connection_7__22__26_, connection_7__22__25_,
         connection_7__22__24_, connection_7__22__23_, connection_7__22__22_,
         connection_7__22__21_, connection_7__22__20_, connection_7__22__19_,
         connection_7__22__18_, connection_7__22__17_, connection_7__22__16_,
         connection_7__22__15_, connection_7__22__14_, connection_7__22__13_,
         connection_7__22__12_, connection_7__22__11_, connection_7__22__10_,
         connection_7__22__9_, connection_7__22__8_, connection_7__22__7_,
         connection_7__22__6_, connection_7__22__5_, connection_7__22__4_,
         connection_7__22__3_, connection_7__22__2_, connection_7__22__1_,
         connection_7__22__0_, connection_7__23__31_, connection_7__23__30_,
         connection_7__23__29_, connection_7__23__28_, connection_7__23__27_,
         connection_7__23__26_, connection_7__23__25_, connection_7__23__24_,
         connection_7__23__23_, connection_7__23__22_, connection_7__23__21_,
         connection_7__23__20_, connection_7__23__19_, connection_7__23__18_,
         connection_7__23__17_, connection_7__23__16_, connection_7__23__15_,
         connection_7__23__14_, connection_7__23__13_, connection_7__23__12_,
         connection_7__23__11_, connection_7__23__10_, connection_7__23__9_,
         connection_7__23__8_, connection_7__23__7_, connection_7__23__6_,
         connection_7__23__5_, connection_7__23__4_, connection_7__23__3_,
         connection_7__23__2_, connection_7__23__1_, connection_7__23__0_,
         connection_7__24__31_, connection_7__24__30_, connection_7__24__29_,
         connection_7__24__28_, connection_7__24__27_, connection_7__24__26_,
         connection_7__24__25_, connection_7__24__24_, connection_7__24__23_,
         connection_7__24__22_, connection_7__24__21_, connection_7__24__20_,
         connection_7__24__19_, connection_7__24__18_, connection_7__24__17_,
         connection_7__24__16_, connection_7__24__15_, connection_7__24__14_,
         connection_7__24__13_, connection_7__24__12_, connection_7__24__11_,
         connection_7__24__10_, connection_7__24__9_, connection_7__24__8_,
         connection_7__24__7_, connection_7__24__6_, connection_7__24__5_,
         connection_7__24__4_, connection_7__24__3_, connection_7__24__2_,
         connection_7__24__1_, connection_7__24__0_, connection_7__25__31_,
         connection_7__25__30_, connection_7__25__29_, connection_7__25__28_,
         connection_7__25__27_, connection_7__25__26_, connection_7__25__25_,
         connection_7__25__24_, connection_7__25__23_, connection_7__25__22_,
         connection_7__25__21_, connection_7__25__20_, connection_7__25__19_,
         connection_7__25__18_, connection_7__25__17_, connection_7__25__16_,
         connection_7__25__15_, connection_7__25__14_, connection_7__25__13_,
         connection_7__25__12_, connection_7__25__11_, connection_7__25__10_,
         connection_7__25__9_, connection_7__25__8_, connection_7__25__7_,
         connection_7__25__6_, connection_7__25__5_, connection_7__25__4_,
         connection_7__25__3_, connection_7__25__2_, connection_7__25__1_,
         connection_7__25__0_, connection_7__26__31_, connection_7__26__30_,
         connection_7__26__29_, connection_7__26__28_, connection_7__26__27_,
         connection_7__26__26_, connection_7__26__25_, connection_7__26__24_,
         connection_7__26__23_, connection_7__26__22_, connection_7__26__21_,
         connection_7__26__20_, connection_7__26__19_, connection_7__26__18_,
         connection_7__26__17_, connection_7__26__16_, connection_7__26__15_,
         connection_7__26__14_, connection_7__26__13_, connection_7__26__12_,
         connection_7__26__11_, connection_7__26__10_, connection_7__26__9_,
         connection_7__26__8_, connection_7__26__7_, connection_7__26__6_,
         connection_7__26__5_, connection_7__26__4_, connection_7__26__3_,
         connection_7__26__2_, connection_7__26__1_, connection_7__26__0_,
         connection_7__27__31_, connection_7__27__30_, connection_7__27__29_,
         connection_7__27__28_, connection_7__27__27_, connection_7__27__26_,
         connection_7__27__25_, connection_7__27__24_, connection_7__27__23_,
         connection_7__27__22_, connection_7__27__21_, connection_7__27__20_,
         connection_7__27__19_, connection_7__27__18_, connection_7__27__17_,
         connection_7__27__16_, connection_7__27__15_, connection_7__27__14_,
         connection_7__27__13_, connection_7__27__12_, connection_7__27__11_,
         connection_7__27__10_, connection_7__27__9_, connection_7__27__8_,
         connection_7__27__7_, connection_7__27__6_, connection_7__27__5_,
         connection_7__27__4_, connection_7__27__3_, connection_7__27__2_,
         connection_7__27__1_, connection_7__27__0_, connection_7__28__31_,
         connection_7__28__30_, connection_7__28__29_, connection_7__28__28_,
         connection_7__28__27_, connection_7__28__26_, connection_7__28__25_,
         connection_7__28__24_, connection_7__28__23_, connection_7__28__22_,
         connection_7__28__21_, connection_7__28__20_, connection_7__28__19_,
         connection_7__28__18_, connection_7__28__17_, connection_7__28__16_,
         connection_7__28__15_, connection_7__28__14_, connection_7__28__13_,
         connection_7__28__12_, connection_7__28__11_, connection_7__28__10_,
         connection_7__28__9_, connection_7__28__8_, connection_7__28__7_,
         connection_7__28__6_, connection_7__28__5_, connection_7__28__4_,
         connection_7__28__3_, connection_7__28__2_, connection_7__28__1_,
         connection_7__28__0_, connection_7__29__31_, connection_7__29__30_,
         connection_7__29__29_, connection_7__29__28_, connection_7__29__27_,
         connection_7__29__26_, connection_7__29__25_, connection_7__29__24_,
         connection_7__29__23_, connection_7__29__22_, connection_7__29__21_,
         connection_7__29__20_, connection_7__29__19_, connection_7__29__18_,
         connection_7__29__17_, connection_7__29__16_, connection_7__29__15_,
         connection_7__29__14_, connection_7__29__13_, connection_7__29__12_,
         connection_7__29__11_, connection_7__29__10_, connection_7__29__9_,
         connection_7__29__8_, connection_7__29__7_, connection_7__29__6_,
         connection_7__29__5_, connection_7__29__4_, connection_7__29__3_,
         connection_7__29__2_, connection_7__29__1_, connection_7__29__0_,
         connection_7__30__31_, connection_7__30__30_, connection_7__30__29_,
         connection_7__30__28_, connection_7__30__27_, connection_7__30__26_,
         connection_7__30__25_, connection_7__30__24_, connection_7__30__23_,
         connection_7__30__22_, connection_7__30__21_, connection_7__30__20_,
         connection_7__30__19_, connection_7__30__18_, connection_7__30__17_,
         connection_7__30__16_, connection_7__30__15_, connection_7__30__14_,
         connection_7__30__13_, connection_7__30__12_, connection_7__30__11_,
         connection_7__30__10_, connection_7__30__9_, connection_7__30__8_,
         connection_7__30__7_, connection_7__30__6_, connection_7__30__5_,
         connection_7__30__4_, connection_7__30__3_, connection_7__30__2_,
         connection_7__30__1_, connection_7__30__0_, connection_7__31__31_,
         connection_7__31__30_, connection_7__31__29_, connection_7__31__28_,
         connection_7__31__27_, connection_7__31__26_, connection_7__31__25_,
         connection_7__31__24_, connection_7__31__23_, connection_7__31__22_,
         connection_7__31__21_, connection_7__31__20_, connection_7__31__19_,
         connection_7__31__18_, connection_7__31__17_, connection_7__31__16_,
         connection_7__31__15_, connection_7__31__14_, connection_7__31__13_,
         connection_7__31__12_, connection_7__31__11_, connection_7__31__10_,
         connection_7__31__9_, connection_7__31__8_, connection_7__31__7_,
         connection_7__31__6_, connection_7__31__5_, connection_7__31__4_,
         connection_7__31__3_, connection_7__31__2_, connection_7__31__1_,
         connection_7__31__0_, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n1538, n1541, n1544, n1547,
         n1550, n1553, n1556, n1559, n1562, n1565, n1568, n1571, n1574, n1577,
         n1580, n1583;
  wire   [255:0] cmd_pipeline_stage_0__pipeline_i_cmd_reg;
  wire   [223:0] cmd_pipeline_stage_1__pipeline_i_cmd_reg;
  wire   [191:0] cmd_pipeline_stage_2__pipeline_i_cmd_reg;
  wire   [159:0] cmd_pipeline_stage_3__pipeline_i_cmd_reg;
  wire   [127:0] cmd_pipeline_stage_4__pipeline_i_cmd_reg;
  wire   [95:0] cmd_pipeline_stage_5__pipeline_i_cmd_reg;
  wire   [63:0] cmd_pipeline_stage_6__pipeline_i_cmd_reg;
  wire   [31:0] cmd_pipeline_stage_7__pipeline_i_cmd_reg;

  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_0 first_stage_switch_0__first_stage ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[1:0]), .i_data_bus(
        i_data_bus[63:0]), .o_valid({connection_valid_0__1_, 
        connection_valid_0__0_}), .o_data_bus({connection_0__1__31_, 
        connection_0__1__30_, connection_0__1__29_, connection_0__1__28_, 
        connection_0__1__27_, connection_0__1__26_, connection_0__1__25_, 
        connection_0__1__24_, connection_0__1__23_, connection_0__1__22_, 
        connection_0__1__21_, connection_0__1__20_, connection_0__1__19_, 
        connection_0__1__18_, connection_0__1__17_, connection_0__1__16_, 
        connection_0__1__15_, connection_0__1__14_, connection_0__1__13_, 
        connection_0__1__12_, connection_0__1__11_, connection_0__1__10_, 
        connection_0__1__9_, connection_0__1__8_, connection_0__1__7_, 
        connection_0__1__6_, connection_0__1__5_, connection_0__1__4_, 
        connection_0__1__3_, connection_0__1__2_, connection_0__1__1_, 
        connection_0__1__0_, connection_0__0__31_, connection_0__0__30_, 
        connection_0__0__29_, connection_0__0__28_, connection_0__0__27_, 
        connection_0__0__26_, connection_0__0__25_, connection_0__0__24_, 
        connection_0__0__23_, connection_0__0__22_, connection_0__0__21_, 
        connection_0__0__20_, connection_0__0__19_, connection_0__0__18_, 
        connection_0__0__17_, connection_0__0__16_, connection_0__0__15_, 
        connection_0__0__14_, connection_0__0__13_, connection_0__0__12_, 
        connection_0__0__11_, connection_0__0__10_, connection_0__0__9_, 
        connection_0__0__8_, connection_0__0__7_, connection_0__0__6_, 
        connection_0__0__5_, connection_0__0__4_, connection_0__0__3_, 
        connection_0__0__2_, connection_0__0__1_, connection_0__0__0_}), 
        .i_en(i_en), .i_cmd(i_cmd[1:0]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_143 first_stage_switch_1__first_stage ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[3:2]), .i_data_bus(
        i_data_bus[127:64]), .o_valid({connection_valid_0__3_, 
        connection_valid_0__2_}), .o_data_bus({connection_0__3__31_, 
        connection_0__3__30_, connection_0__3__29_, connection_0__3__28_, 
        connection_0__3__27_, connection_0__3__26_, connection_0__3__25_, 
        connection_0__3__24_, connection_0__3__23_, connection_0__3__22_, 
        connection_0__3__21_, connection_0__3__20_, connection_0__3__19_, 
        connection_0__3__18_, connection_0__3__17_, connection_0__3__16_, 
        connection_0__3__15_, connection_0__3__14_, connection_0__3__13_, 
        connection_0__3__12_, connection_0__3__11_, connection_0__3__10_, 
        connection_0__3__9_, connection_0__3__8_, connection_0__3__7_, 
        connection_0__3__6_, connection_0__3__5_, connection_0__3__4_, 
        connection_0__3__3_, connection_0__3__2_, connection_0__3__1_, 
        connection_0__3__0_, connection_0__2__31_, connection_0__2__30_, 
        connection_0__2__29_, connection_0__2__28_, connection_0__2__27_, 
        connection_0__2__26_, connection_0__2__25_, connection_0__2__24_, 
        connection_0__2__23_, connection_0__2__22_, connection_0__2__21_, 
        connection_0__2__20_, connection_0__2__19_, connection_0__2__18_, 
        connection_0__2__17_, connection_0__2__16_, connection_0__2__15_, 
        connection_0__2__14_, connection_0__2__13_, connection_0__2__12_, 
        connection_0__2__11_, connection_0__2__10_, connection_0__2__9_, 
        connection_0__2__8_, connection_0__2__7_, connection_0__2__6_, 
        connection_0__2__5_, connection_0__2__4_, connection_0__2__3_, 
        connection_0__2__2_, connection_0__2__1_, connection_0__2__0_}), 
        .i_en(i_en), .i_cmd(i_cmd[3:2]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_142 first_stage_switch_2__first_stage ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[5:4]), .i_data_bus(
        i_data_bus[191:128]), .o_valid({connection_valid_0__5_, 
        connection_valid_0__4_}), .o_data_bus({connection_0__5__31_, 
        connection_0__5__30_, connection_0__5__29_, connection_0__5__28_, 
        connection_0__5__27_, connection_0__5__26_, connection_0__5__25_, 
        connection_0__5__24_, connection_0__5__23_, connection_0__5__22_, 
        connection_0__5__21_, connection_0__5__20_, connection_0__5__19_, 
        connection_0__5__18_, connection_0__5__17_, connection_0__5__16_, 
        connection_0__5__15_, connection_0__5__14_, connection_0__5__13_, 
        connection_0__5__12_, connection_0__5__11_, connection_0__5__10_, 
        connection_0__5__9_, connection_0__5__8_, connection_0__5__7_, 
        connection_0__5__6_, connection_0__5__5_, connection_0__5__4_, 
        connection_0__5__3_, connection_0__5__2_, connection_0__5__1_, 
        connection_0__5__0_, connection_0__4__31_, connection_0__4__30_, 
        connection_0__4__29_, connection_0__4__28_, connection_0__4__27_, 
        connection_0__4__26_, connection_0__4__25_, connection_0__4__24_, 
        connection_0__4__23_, connection_0__4__22_, connection_0__4__21_, 
        connection_0__4__20_, connection_0__4__19_, connection_0__4__18_, 
        connection_0__4__17_, connection_0__4__16_, connection_0__4__15_, 
        connection_0__4__14_, connection_0__4__13_, connection_0__4__12_, 
        connection_0__4__11_, connection_0__4__10_, connection_0__4__9_, 
        connection_0__4__8_, connection_0__4__7_, connection_0__4__6_, 
        connection_0__4__5_, connection_0__4__4_, connection_0__4__3_, 
        connection_0__4__2_, connection_0__4__1_, connection_0__4__0_}), 
        .i_en(i_en), .i_cmd(i_cmd[5:4]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_141 first_stage_switch_3__first_stage ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[7:6]), .i_data_bus(
        i_data_bus[255:192]), .o_valid({connection_valid_0__7_, 
        connection_valid_0__6_}), .o_data_bus({connection_0__7__31_, 
        connection_0__7__30_, connection_0__7__29_, connection_0__7__28_, 
        connection_0__7__27_, connection_0__7__26_, connection_0__7__25_, 
        connection_0__7__24_, connection_0__7__23_, connection_0__7__22_, 
        connection_0__7__21_, connection_0__7__20_, connection_0__7__19_, 
        connection_0__7__18_, connection_0__7__17_, connection_0__7__16_, 
        connection_0__7__15_, connection_0__7__14_, connection_0__7__13_, 
        connection_0__7__12_, connection_0__7__11_, connection_0__7__10_, 
        connection_0__7__9_, connection_0__7__8_, connection_0__7__7_, 
        connection_0__7__6_, connection_0__7__5_, connection_0__7__4_, 
        connection_0__7__3_, connection_0__7__2_, connection_0__7__1_, 
        connection_0__7__0_, connection_0__6__31_, connection_0__6__30_, 
        connection_0__6__29_, connection_0__6__28_, connection_0__6__27_, 
        connection_0__6__26_, connection_0__6__25_, connection_0__6__24_, 
        connection_0__6__23_, connection_0__6__22_, connection_0__6__21_, 
        connection_0__6__20_, connection_0__6__19_, connection_0__6__18_, 
        connection_0__6__17_, connection_0__6__16_, connection_0__6__15_, 
        connection_0__6__14_, connection_0__6__13_, connection_0__6__12_, 
        connection_0__6__11_, connection_0__6__10_, connection_0__6__9_, 
        connection_0__6__8_, connection_0__6__7_, connection_0__6__6_, 
        connection_0__6__5_, connection_0__6__4_, connection_0__6__3_, 
        connection_0__6__2_, connection_0__6__1_, connection_0__6__0_}), 
        .i_en(i_en), .i_cmd(i_cmd[7:6]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_140 first_stage_switch_4__first_stage ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[9:8]), .i_data_bus(
        i_data_bus[319:256]), .o_valid({connection_valid_0__9_, 
        connection_valid_0__8_}), .o_data_bus({connection_0__9__31_, 
        connection_0__9__30_, connection_0__9__29_, connection_0__9__28_, 
        connection_0__9__27_, connection_0__9__26_, connection_0__9__25_, 
        connection_0__9__24_, connection_0__9__23_, connection_0__9__22_, 
        connection_0__9__21_, connection_0__9__20_, connection_0__9__19_, 
        connection_0__9__18_, connection_0__9__17_, connection_0__9__16_, 
        connection_0__9__15_, connection_0__9__14_, connection_0__9__13_, 
        connection_0__9__12_, connection_0__9__11_, connection_0__9__10_, 
        connection_0__9__9_, connection_0__9__8_, connection_0__9__7_, 
        connection_0__9__6_, connection_0__9__5_, connection_0__9__4_, 
        connection_0__9__3_, connection_0__9__2_, connection_0__9__1_, 
        connection_0__9__0_, connection_0__8__31_, connection_0__8__30_, 
        connection_0__8__29_, connection_0__8__28_, connection_0__8__27_, 
        connection_0__8__26_, connection_0__8__25_, connection_0__8__24_, 
        connection_0__8__23_, connection_0__8__22_, connection_0__8__21_, 
        connection_0__8__20_, connection_0__8__19_, connection_0__8__18_, 
        connection_0__8__17_, connection_0__8__16_, connection_0__8__15_, 
        connection_0__8__14_, connection_0__8__13_, connection_0__8__12_, 
        connection_0__8__11_, connection_0__8__10_, connection_0__8__9_, 
        connection_0__8__8_, connection_0__8__7_, connection_0__8__6_, 
        connection_0__8__5_, connection_0__8__4_, connection_0__8__3_, 
        connection_0__8__2_, connection_0__8__1_, connection_0__8__0_}), 
        .i_en(i_en), .i_cmd(i_cmd[9:8]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_139 first_stage_switch_5__first_stage ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[11:10]), .i_data_bus(
        i_data_bus[383:320]), .o_valid({connection_valid_0__11_, 
        connection_valid_0__10_}), .o_data_bus({connection_0__11__31_, 
        connection_0__11__30_, connection_0__11__29_, connection_0__11__28_, 
        connection_0__11__27_, connection_0__11__26_, connection_0__11__25_, 
        connection_0__11__24_, connection_0__11__23_, connection_0__11__22_, 
        connection_0__11__21_, connection_0__11__20_, connection_0__11__19_, 
        connection_0__11__18_, connection_0__11__17_, connection_0__11__16_, 
        connection_0__11__15_, connection_0__11__14_, connection_0__11__13_, 
        connection_0__11__12_, connection_0__11__11_, connection_0__11__10_, 
        connection_0__11__9_, connection_0__11__8_, connection_0__11__7_, 
        connection_0__11__6_, connection_0__11__5_, connection_0__11__4_, 
        connection_0__11__3_, connection_0__11__2_, connection_0__11__1_, 
        connection_0__11__0_, connection_0__10__31_, connection_0__10__30_, 
        connection_0__10__29_, connection_0__10__28_, connection_0__10__27_, 
        connection_0__10__26_, connection_0__10__25_, connection_0__10__24_, 
        connection_0__10__23_, connection_0__10__22_, connection_0__10__21_, 
        connection_0__10__20_, connection_0__10__19_, connection_0__10__18_, 
        connection_0__10__17_, connection_0__10__16_, connection_0__10__15_, 
        connection_0__10__14_, connection_0__10__13_, connection_0__10__12_, 
        connection_0__10__11_, connection_0__10__10_, connection_0__10__9_, 
        connection_0__10__8_, connection_0__10__7_, connection_0__10__6_, 
        connection_0__10__5_, connection_0__10__4_, connection_0__10__3_, 
        connection_0__10__2_, connection_0__10__1_, connection_0__10__0_}), 
        .i_en(i_en), .i_cmd(i_cmd[11:10]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_138 first_stage_switch_6__first_stage ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[13:12]), .i_data_bus(
        i_data_bus[447:384]), .o_valid({connection_valid_0__13_, 
        connection_valid_0__12_}), .o_data_bus({connection_0__13__31_, 
        connection_0__13__30_, connection_0__13__29_, connection_0__13__28_, 
        connection_0__13__27_, connection_0__13__26_, connection_0__13__25_, 
        connection_0__13__24_, connection_0__13__23_, connection_0__13__22_, 
        connection_0__13__21_, connection_0__13__20_, connection_0__13__19_, 
        connection_0__13__18_, connection_0__13__17_, connection_0__13__16_, 
        connection_0__13__15_, connection_0__13__14_, connection_0__13__13_, 
        connection_0__13__12_, connection_0__13__11_, connection_0__13__10_, 
        connection_0__13__9_, connection_0__13__8_, connection_0__13__7_, 
        connection_0__13__6_, connection_0__13__5_, connection_0__13__4_, 
        connection_0__13__3_, connection_0__13__2_, connection_0__13__1_, 
        connection_0__13__0_, connection_0__12__31_, connection_0__12__30_, 
        connection_0__12__29_, connection_0__12__28_, connection_0__12__27_, 
        connection_0__12__26_, connection_0__12__25_, connection_0__12__24_, 
        connection_0__12__23_, connection_0__12__22_, connection_0__12__21_, 
        connection_0__12__20_, connection_0__12__19_, connection_0__12__18_, 
        connection_0__12__17_, connection_0__12__16_, connection_0__12__15_, 
        connection_0__12__14_, connection_0__12__13_, connection_0__12__12_, 
        connection_0__12__11_, connection_0__12__10_, connection_0__12__9_, 
        connection_0__12__8_, connection_0__12__7_, connection_0__12__6_, 
        connection_0__12__5_, connection_0__12__4_, connection_0__12__3_, 
        connection_0__12__2_, connection_0__12__1_, connection_0__12__0_}), 
        .i_en(i_en), .i_cmd(i_cmd[13:12]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_137 first_stage_switch_7__first_stage ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[15:14]), .i_data_bus(
        i_data_bus[511:448]), .o_valid({connection_valid_0__15_, 
        connection_valid_0__14_}), .o_data_bus({connection_0__15__31_, 
        connection_0__15__30_, connection_0__15__29_, connection_0__15__28_, 
        connection_0__15__27_, connection_0__15__26_, connection_0__15__25_, 
        connection_0__15__24_, connection_0__15__23_, connection_0__15__22_, 
        connection_0__15__21_, connection_0__15__20_, connection_0__15__19_, 
        connection_0__15__18_, connection_0__15__17_, connection_0__15__16_, 
        connection_0__15__15_, connection_0__15__14_, connection_0__15__13_, 
        connection_0__15__12_, connection_0__15__11_, connection_0__15__10_, 
        connection_0__15__9_, connection_0__15__8_, connection_0__15__7_, 
        connection_0__15__6_, connection_0__15__5_, connection_0__15__4_, 
        connection_0__15__3_, connection_0__15__2_, connection_0__15__1_, 
        connection_0__15__0_, connection_0__14__31_, connection_0__14__30_, 
        connection_0__14__29_, connection_0__14__28_, connection_0__14__27_, 
        connection_0__14__26_, connection_0__14__25_, connection_0__14__24_, 
        connection_0__14__23_, connection_0__14__22_, connection_0__14__21_, 
        connection_0__14__20_, connection_0__14__19_, connection_0__14__18_, 
        connection_0__14__17_, connection_0__14__16_, connection_0__14__15_, 
        connection_0__14__14_, connection_0__14__13_, connection_0__14__12_, 
        connection_0__14__11_, connection_0__14__10_, connection_0__14__9_, 
        connection_0__14__8_, connection_0__14__7_, connection_0__14__6_, 
        connection_0__14__5_, connection_0__14__4_, connection_0__14__3_, 
        connection_0__14__2_, connection_0__14__1_, connection_0__14__0_}), 
        .i_en(i_en), .i_cmd(i_cmd[15:14]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_136 first_stage_switch_8__first_stage ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[17:16]), .i_data_bus(
        i_data_bus[575:512]), .o_valid({connection_valid_0__17_, 
        connection_valid_0__16_}), .o_data_bus({connection_0__17__31_, 
        connection_0__17__30_, connection_0__17__29_, connection_0__17__28_, 
        connection_0__17__27_, connection_0__17__26_, connection_0__17__25_, 
        connection_0__17__24_, connection_0__17__23_, connection_0__17__22_, 
        connection_0__17__21_, connection_0__17__20_, connection_0__17__19_, 
        connection_0__17__18_, connection_0__17__17_, connection_0__17__16_, 
        connection_0__17__15_, connection_0__17__14_, connection_0__17__13_, 
        connection_0__17__12_, connection_0__17__11_, connection_0__17__10_, 
        connection_0__17__9_, connection_0__17__8_, connection_0__17__7_, 
        connection_0__17__6_, connection_0__17__5_, connection_0__17__4_, 
        connection_0__17__3_, connection_0__17__2_, connection_0__17__1_, 
        connection_0__17__0_, connection_0__16__31_, connection_0__16__30_, 
        connection_0__16__29_, connection_0__16__28_, connection_0__16__27_, 
        connection_0__16__26_, connection_0__16__25_, connection_0__16__24_, 
        connection_0__16__23_, connection_0__16__22_, connection_0__16__21_, 
        connection_0__16__20_, connection_0__16__19_, connection_0__16__18_, 
        connection_0__16__17_, connection_0__16__16_, connection_0__16__15_, 
        connection_0__16__14_, connection_0__16__13_, connection_0__16__12_, 
        connection_0__16__11_, connection_0__16__10_, connection_0__16__9_, 
        connection_0__16__8_, connection_0__16__7_, connection_0__16__6_, 
        connection_0__16__5_, connection_0__16__4_, connection_0__16__3_, 
        connection_0__16__2_, connection_0__16__1_, connection_0__16__0_}), 
        .i_en(i_en), .i_cmd(i_cmd[17:16]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_135 first_stage_switch_9__first_stage ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[19:18]), .i_data_bus(
        i_data_bus[639:576]), .o_valid({connection_valid_0__19_, 
        connection_valid_0__18_}), .o_data_bus({connection_0__19__31_, 
        connection_0__19__30_, connection_0__19__29_, connection_0__19__28_, 
        connection_0__19__27_, connection_0__19__26_, connection_0__19__25_, 
        connection_0__19__24_, connection_0__19__23_, connection_0__19__22_, 
        connection_0__19__21_, connection_0__19__20_, connection_0__19__19_, 
        connection_0__19__18_, connection_0__19__17_, connection_0__19__16_, 
        connection_0__19__15_, connection_0__19__14_, connection_0__19__13_, 
        connection_0__19__12_, connection_0__19__11_, connection_0__19__10_, 
        connection_0__19__9_, connection_0__19__8_, connection_0__19__7_, 
        connection_0__19__6_, connection_0__19__5_, connection_0__19__4_, 
        connection_0__19__3_, connection_0__19__2_, connection_0__19__1_, 
        connection_0__19__0_, connection_0__18__31_, connection_0__18__30_, 
        connection_0__18__29_, connection_0__18__28_, connection_0__18__27_, 
        connection_0__18__26_, connection_0__18__25_, connection_0__18__24_, 
        connection_0__18__23_, connection_0__18__22_, connection_0__18__21_, 
        connection_0__18__20_, connection_0__18__19_, connection_0__18__18_, 
        connection_0__18__17_, connection_0__18__16_, connection_0__18__15_, 
        connection_0__18__14_, connection_0__18__13_, connection_0__18__12_, 
        connection_0__18__11_, connection_0__18__10_, connection_0__18__9_, 
        connection_0__18__8_, connection_0__18__7_, connection_0__18__6_, 
        connection_0__18__5_, connection_0__18__4_, connection_0__18__3_, 
        connection_0__18__2_, connection_0__18__1_, connection_0__18__0_}), 
        .i_en(i_en), .i_cmd(i_cmd[19:18]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_134 first_stage_switch_10__first_stage ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[21:20]), .i_data_bus(
        i_data_bus[703:640]), .o_valid({connection_valid_0__21_, 
        connection_valid_0__20_}), .o_data_bus({connection_0__21__31_, 
        connection_0__21__30_, connection_0__21__29_, connection_0__21__28_, 
        connection_0__21__27_, connection_0__21__26_, connection_0__21__25_, 
        connection_0__21__24_, connection_0__21__23_, connection_0__21__22_, 
        connection_0__21__21_, connection_0__21__20_, connection_0__21__19_, 
        connection_0__21__18_, connection_0__21__17_, connection_0__21__16_, 
        connection_0__21__15_, connection_0__21__14_, connection_0__21__13_, 
        connection_0__21__12_, connection_0__21__11_, connection_0__21__10_, 
        connection_0__21__9_, connection_0__21__8_, connection_0__21__7_, 
        connection_0__21__6_, connection_0__21__5_, connection_0__21__4_, 
        connection_0__21__3_, connection_0__21__2_, connection_0__21__1_, 
        connection_0__21__0_, connection_0__20__31_, connection_0__20__30_, 
        connection_0__20__29_, connection_0__20__28_, connection_0__20__27_, 
        connection_0__20__26_, connection_0__20__25_, connection_0__20__24_, 
        connection_0__20__23_, connection_0__20__22_, connection_0__20__21_, 
        connection_0__20__20_, connection_0__20__19_, connection_0__20__18_, 
        connection_0__20__17_, connection_0__20__16_, connection_0__20__15_, 
        connection_0__20__14_, connection_0__20__13_, connection_0__20__12_, 
        connection_0__20__11_, connection_0__20__10_, connection_0__20__9_, 
        connection_0__20__8_, connection_0__20__7_, connection_0__20__6_, 
        connection_0__20__5_, connection_0__20__4_, connection_0__20__3_, 
        connection_0__20__2_, connection_0__20__1_, connection_0__20__0_}), 
        .i_en(i_en), .i_cmd(i_cmd[21:20]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_133 first_stage_switch_11__first_stage ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[23:22]), .i_data_bus(
        i_data_bus[767:704]), .o_valid({connection_valid_0__23_, 
        connection_valid_0__22_}), .o_data_bus({connection_0__23__31_, 
        connection_0__23__30_, connection_0__23__29_, connection_0__23__28_, 
        connection_0__23__27_, connection_0__23__26_, connection_0__23__25_, 
        connection_0__23__24_, connection_0__23__23_, connection_0__23__22_, 
        connection_0__23__21_, connection_0__23__20_, connection_0__23__19_, 
        connection_0__23__18_, connection_0__23__17_, connection_0__23__16_, 
        connection_0__23__15_, connection_0__23__14_, connection_0__23__13_, 
        connection_0__23__12_, connection_0__23__11_, connection_0__23__10_, 
        connection_0__23__9_, connection_0__23__8_, connection_0__23__7_, 
        connection_0__23__6_, connection_0__23__5_, connection_0__23__4_, 
        connection_0__23__3_, connection_0__23__2_, connection_0__23__1_, 
        connection_0__23__0_, connection_0__22__31_, connection_0__22__30_, 
        connection_0__22__29_, connection_0__22__28_, connection_0__22__27_, 
        connection_0__22__26_, connection_0__22__25_, connection_0__22__24_, 
        connection_0__22__23_, connection_0__22__22_, connection_0__22__21_, 
        connection_0__22__20_, connection_0__22__19_, connection_0__22__18_, 
        connection_0__22__17_, connection_0__22__16_, connection_0__22__15_, 
        connection_0__22__14_, connection_0__22__13_, connection_0__22__12_, 
        connection_0__22__11_, connection_0__22__10_, connection_0__22__9_, 
        connection_0__22__8_, connection_0__22__7_, connection_0__22__6_, 
        connection_0__22__5_, connection_0__22__4_, connection_0__22__3_, 
        connection_0__22__2_, connection_0__22__1_, connection_0__22__0_}), 
        .i_en(i_en), .i_cmd(i_cmd[23:22]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_132 first_stage_switch_12__first_stage ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[25:24]), .i_data_bus(
        i_data_bus[831:768]), .o_valid({connection_valid_0__25_, 
        connection_valid_0__24_}), .o_data_bus({connection_0__25__31_, 
        connection_0__25__30_, connection_0__25__29_, connection_0__25__28_, 
        connection_0__25__27_, connection_0__25__26_, connection_0__25__25_, 
        connection_0__25__24_, connection_0__25__23_, connection_0__25__22_, 
        connection_0__25__21_, connection_0__25__20_, connection_0__25__19_, 
        connection_0__25__18_, connection_0__25__17_, connection_0__25__16_, 
        connection_0__25__15_, connection_0__25__14_, connection_0__25__13_, 
        connection_0__25__12_, connection_0__25__11_, connection_0__25__10_, 
        connection_0__25__9_, connection_0__25__8_, connection_0__25__7_, 
        connection_0__25__6_, connection_0__25__5_, connection_0__25__4_, 
        connection_0__25__3_, connection_0__25__2_, connection_0__25__1_, 
        connection_0__25__0_, connection_0__24__31_, connection_0__24__30_, 
        connection_0__24__29_, connection_0__24__28_, connection_0__24__27_, 
        connection_0__24__26_, connection_0__24__25_, connection_0__24__24_, 
        connection_0__24__23_, connection_0__24__22_, connection_0__24__21_, 
        connection_0__24__20_, connection_0__24__19_, connection_0__24__18_, 
        connection_0__24__17_, connection_0__24__16_, connection_0__24__15_, 
        connection_0__24__14_, connection_0__24__13_, connection_0__24__12_, 
        connection_0__24__11_, connection_0__24__10_, connection_0__24__9_, 
        connection_0__24__8_, connection_0__24__7_, connection_0__24__6_, 
        connection_0__24__5_, connection_0__24__4_, connection_0__24__3_, 
        connection_0__24__2_, connection_0__24__1_, connection_0__24__0_}), 
        .i_en(i_en), .i_cmd(i_cmd[25:24]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_131 first_stage_switch_13__first_stage ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[27:26]), .i_data_bus(
        i_data_bus[895:832]), .o_valid({connection_valid_0__27_, 
        connection_valid_0__26_}), .o_data_bus({connection_0__27__31_, 
        connection_0__27__30_, connection_0__27__29_, connection_0__27__28_, 
        connection_0__27__27_, connection_0__27__26_, connection_0__27__25_, 
        connection_0__27__24_, connection_0__27__23_, connection_0__27__22_, 
        connection_0__27__21_, connection_0__27__20_, connection_0__27__19_, 
        connection_0__27__18_, connection_0__27__17_, connection_0__27__16_, 
        connection_0__27__15_, connection_0__27__14_, connection_0__27__13_, 
        connection_0__27__12_, connection_0__27__11_, connection_0__27__10_, 
        connection_0__27__9_, connection_0__27__8_, connection_0__27__7_, 
        connection_0__27__6_, connection_0__27__5_, connection_0__27__4_, 
        connection_0__27__3_, connection_0__27__2_, connection_0__27__1_, 
        connection_0__27__0_, connection_0__26__31_, connection_0__26__30_, 
        connection_0__26__29_, connection_0__26__28_, connection_0__26__27_, 
        connection_0__26__26_, connection_0__26__25_, connection_0__26__24_, 
        connection_0__26__23_, connection_0__26__22_, connection_0__26__21_, 
        connection_0__26__20_, connection_0__26__19_, connection_0__26__18_, 
        connection_0__26__17_, connection_0__26__16_, connection_0__26__15_, 
        connection_0__26__14_, connection_0__26__13_, connection_0__26__12_, 
        connection_0__26__11_, connection_0__26__10_, connection_0__26__9_, 
        connection_0__26__8_, connection_0__26__7_, connection_0__26__6_, 
        connection_0__26__5_, connection_0__26__4_, connection_0__26__3_, 
        connection_0__26__2_, connection_0__26__1_, connection_0__26__0_}), 
        .i_en(i_en), .i_cmd(i_cmd[27:26]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_130 first_stage_switch_14__first_stage ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[29:28]), .i_data_bus(
        i_data_bus[959:896]), .o_valid({connection_valid_0__29_, 
        connection_valid_0__28_}), .o_data_bus({connection_0__29__31_, 
        connection_0__29__30_, connection_0__29__29_, connection_0__29__28_, 
        connection_0__29__27_, connection_0__29__26_, connection_0__29__25_, 
        connection_0__29__24_, connection_0__29__23_, connection_0__29__22_, 
        connection_0__29__21_, connection_0__29__20_, connection_0__29__19_, 
        connection_0__29__18_, connection_0__29__17_, connection_0__29__16_, 
        connection_0__29__15_, connection_0__29__14_, connection_0__29__13_, 
        connection_0__29__12_, connection_0__29__11_, connection_0__29__10_, 
        connection_0__29__9_, connection_0__29__8_, connection_0__29__7_, 
        connection_0__29__6_, connection_0__29__5_, connection_0__29__4_, 
        connection_0__29__3_, connection_0__29__2_, connection_0__29__1_, 
        connection_0__29__0_, connection_0__28__31_, connection_0__28__30_, 
        connection_0__28__29_, connection_0__28__28_, connection_0__28__27_, 
        connection_0__28__26_, connection_0__28__25_, connection_0__28__24_, 
        connection_0__28__23_, connection_0__28__22_, connection_0__28__21_, 
        connection_0__28__20_, connection_0__28__19_, connection_0__28__18_, 
        connection_0__28__17_, connection_0__28__16_, connection_0__28__15_, 
        connection_0__28__14_, connection_0__28__13_, connection_0__28__12_, 
        connection_0__28__11_, connection_0__28__10_, connection_0__28__9_, 
        connection_0__28__8_, connection_0__28__7_, connection_0__28__6_, 
        connection_0__28__5_, connection_0__28__4_, connection_0__28__3_, 
        connection_0__28__2_, connection_0__28__1_, connection_0__28__0_}), 
        .i_en(i_en), .i_cmd(i_cmd[29:28]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_129 first_stage_switch_15__first_stage ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[31:30]), .i_data_bus(
        i_data_bus[1023:960]), .o_valid({connection_valid_0__31_, 
        connection_valid_0__30_}), .o_data_bus({connection_0__31__31_, 
        connection_0__31__30_, connection_0__31__29_, connection_0__31__28_, 
        connection_0__31__27_, connection_0__31__26_, connection_0__31__25_, 
        connection_0__31__24_, connection_0__31__23_, connection_0__31__22_, 
        connection_0__31__21_, connection_0__31__20_, connection_0__31__19_, 
        connection_0__31__18_, connection_0__31__17_, connection_0__31__16_, 
        connection_0__31__15_, connection_0__31__14_, connection_0__31__13_, 
        connection_0__31__12_, connection_0__31__11_, connection_0__31__10_, 
        connection_0__31__9_, connection_0__31__8_, connection_0__31__7_, 
        connection_0__31__6_, connection_0__31__5_, connection_0__31__4_, 
        connection_0__31__3_, connection_0__31__2_, connection_0__31__1_, 
        connection_0__31__0_, connection_0__30__31_, connection_0__30__30_, 
        connection_0__30__29_, connection_0__30__28_, connection_0__30__27_, 
        connection_0__30__26_, connection_0__30__25_, connection_0__30__24_, 
        connection_0__30__23_, connection_0__30__22_, connection_0__30__21_, 
        connection_0__30__20_, connection_0__30__19_, connection_0__30__18_, 
        connection_0__30__17_, connection_0__30__16_, connection_0__30__15_, 
        connection_0__30__14_, connection_0__30__13_, connection_0__30__12_, 
        connection_0__30__11_, connection_0__30__10_, connection_0__30__9_, 
        connection_0__30__8_, connection_0__30__7_, connection_0__30__6_, 
        connection_0__30__5_, connection_0__30__4_, connection_0__30__3_, 
        connection_0__30__2_, connection_0__30__1_, connection_0__30__0_}), 
        .i_en(i_en), .i_cmd(i_cmd[31:30]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_128 first_half_stages_0__group_first_half_0__switch_first_half_0__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__2_, 
        connection_valid_0__0_}), .i_data_bus({connection_0__2__31_, 
        connection_0__2__30_, connection_0__2__29_, connection_0__2__28_, 
        connection_0__2__27_, connection_0__2__26_, connection_0__2__25_, 
        connection_0__2__24_, connection_0__2__23_, connection_0__2__22_, 
        connection_0__2__21_, connection_0__2__20_, connection_0__2__19_, 
        connection_0__2__18_, connection_0__2__17_, connection_0__2__16_, 
        connection_0__2__15_, connection_0__2__14_, connection_0__2__13_, 
        connection_0__2__12_, connection_0__2__11_, connection_0__2__10_, 
        connection_0__2__9_, connection_0__2__8_, connection_0__2__7_, 
        connection_0__2__6_, connection_0__2__5_, connection_0__2__4_, 
        connection_0__2__3_, connection_0__2__2_, connection_0__2__1_, 
        connection_0__2__0_, connection_0__0__31_, connection_0__0__30_, 
        connection_0__0__29_, connection_0__0__28_, connection_0__0__27_, 
        connection_0__0__26_, connection_0__0__25_, connection_0__0__24_, 
        connection_0__0__23_, connection_0__0__22_, connection_0__0__21_, 
        connection_0__0__20_, connection_0__0__19_, connection_0__0__18_, 
        connection_0__0__17_, connection_0__0__16_, connection_0__0__15_, 
        connection_0__0__14_, connection_0__0__13_, connection_0__0__12_, 
        connection_0__0__11_, connection_0__0__10_, connection_0__0__9_, 
        connection_0__0__8_, connection_0__0__7_, connection_0__0__6_, 
        connection_0__0__5_, connection_0__0__4_, connection_0__0__3_, 
        connection_0__0__2_, connection_0__0__1_, connection_0__0__0_}), 
        .o_valid({connection_valid_1__1_, connection_valid_1__0_}), 
        .o_data_bus({connection_1__1__31_, connection_1__1__30_, 
        connection_1__1__29_, connection_1__1__28_, connection_1__1__27_, 
        connection_1__1__26_, connection_1__1__25_, connection_1__1__24_, 
        connection_1__1__23_, connection_1__1__22_, connection_1__1__21_, 
        connection_1__1__20_, connection_1__1__19_, connection_1__1__18_, 
        connection_1__1__17_, connection_1__1__16_, connection_1__1__15_, 
        connection_1__1__14_, connection_1__1__13_, connection_1__1__12_, 
        connection_1__1__11_, connection_1__1__10_, connection_1__1__9_, 
        connection_1__1__8_, connection_1__1__7_, connection_1__1__6_, 
        connection_1__1__5_, connection_1__1__4_, connection_1__1__3_, 
        connection_1__1__2_, connection_1__1__1_, connection_1__1__0_, 
        connection_1__0__31_, connection_1__0__30_, connection_1__0__29_, 
        connection_1__0__28_, connection_1__0__27_, connection_1__0__26_, 
        connection_1__0__25_, connection_1__0__24_, connection_1__0__23_, 
        connection_1__0__22_, connection_1__0__21_, connection_1__0__20_, 
        connection_1__0__19_, connection_1__0__18_, connection_1__0__17_, 
        connection_1__0__16_, connection_1__0__15_, connection_1__0__14_, 
        connection_1__0__13_, connection_1__0__12_, connection_1__0__11_, 
        connection_1__0__10_, connection_1__0__9_, connection_1__0__8_, 
        connection_1__0__7_, connection_1__0__6_, connection_1__0__5_, 
        connection_1__0__4_, connection_1__0__3_, connection_1__0__2_, 
        connection_1__0__1_, connection_1__0__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[255:254]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_127 first_half_stages_0__group_first_half_0__switch_first_half_1__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__6_, 
        connection_valid_0__4_}), .i_data_bus({connection_0__6__31_, 
        connection_0__6__30_, connection_0__6__29_, connection_0__6__28_, 
        connection_0__6__27_, connection_0__6__26_, connection_0__6__25_, 
        connection_0__6__24_, connection_0__6__23_, connection_0__6__22_, 
        connection_0__6__21_, connection_0__6__20_, connection_0__6__19_, 
        connection_0__6__18_, connection_0__6__17_, connection_0__6__16_, 
        connection_0__6__15_, connection_0__6__14_, connection_0__6__13_, 
        connection_0__6__12_, connection_0__6__11_, connection_0__6__10_, 
        connection_0__6__9_, connection_0__6__8_, connection_0__6__7_, 
        connection_0__6__6_, connection_0__6__5_, connection_0__6__4_, 
        connection_0__6__3_, connection_0__6__2_, connection_0__6__1_, 
        connection_0__6__0_, connection_0__4__31_, connection_0__4__30_, 
        connection_0__4__29_, connection_0__4__28_, connection_0__4__27_, 
        connection_0__4__26_, connection_0__4__25_, connection_0__4__24_, 
        connection_0__4__23_, connection_0__4__22_, connection_0__4__21_, 
        connection_0__4__20_, connection_0__4__19_, connection_0__4__18_, 
        connection_0__4__17_, connection_0__4__16_, connection_0__4__15_, 
        connection_0__4__14_, connection_0__4__13_, connection_0__4__12_, 
        connection_0__4__11_, connection_0__4__10_, connection_0__4__9_, 
        connection_0__4__8_, connection_0__4__7_, connection_0__4__6_, 
        connection_0__4__5_, connection_0__4__4_, connection_0__4__3_, 
        connection_0__4__2_, connection_0__4__1_, connection_0__4__0_}), 
        .o_valid({connection_valid_1__3_, connection_valid_1__2_}), 
        .o_data_bus({connection_1__3__31_, connection_1__3__30_, 
        connection_1__3__29_, connection_1__3__28_, connection_1__3__27_, 
        connection_1__3__26_, connection_1__3__25_, connection_1__3__24_, 
        connection_1__3__23_, connection_1__3__22_, connection_1__3__21_, 
        connection_1__3__20_, connection_1__3__19_, connection_1__3__18_, 
        connection_1__3__17_, connection_1__3__16_, connection_1__3__15_, 
        connection_1__3__14_, connection_1__3__13_, connection_1__3__12_, 
        connection_1__3__11_, connection_1__3__10_, connection_1__3__9_, 
        connection_1__3__8_, connection_1__3__7_, connection_1__3__6_, 
        connection_1__3__5_, connection_1__3__4_, connection_1__3__3_, 
        connection_1__3__2_, connection_1__3__1_, connection_1__3__0_, 
        connection_1__2__31_, connection_1__2__30_, connection_1__2__29_, 
        connection_1__2__28_, connection_1__2__27_, connection_1__2__26_, 
        connection_1__2__25_, connection_1__2__24_, connection_1__2__23_, 
        connection_1__2__22_, connection_1__2__21_, connection_1__2__20_, 
        connection_1__2__19_, connection_1__2__18_, connection_1__2__17_, 
        connection_1__2__16_, connection_1__2__15_, connection_1__2__14_, 
        connection_1__2__13_, connection_1__2__12_, connection_1__2__11_, 
        connection_1__2__10_, connection_1__2__9_, connection_1__2__8_, 
        connection_1__2__7_, connection_1__2__6_, connection_1__2__5_, 
        connection_1__2__4_, connection_1__2__3_, connection_1__2__2_, 
        connection_1__2__1_, connection_1__2__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[253:252]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_126 first_half_stages_0__group_first_half_0__switch_first_half_2__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__10_, 
        connection_valid_0__8_}), .i_data_bus({connection_0__10__31_, 
        connection_0__10__30_, connection_0__10__29_, connection_0__10__28_, 
        connection_0__10__27_, connection_0__10__26_, connection_0__10__25_, 
        connection_0__10__24_, connection_0__10__23_, connection_0__10__22_, 
        connection_0__10__21_, connection_0__10__20_, connection_0__10__19_, 
        connection_0__10__18_, connection_0__10__17_, connection_0__10__16_, 
        connection_0__10__15_, connection_0__10__14_, connection_0__10__13_, 
        connection_0__10__12_, connection_0__10__11_, connection_0__10__10_, 
        connection_0__10__9_, connection_0__10__8_, connection_0__10__7_, 
        connection_0__10__6_, connection_0__10__5_, connection_0__10__4_, 
        connection_0__10__3_, connection_0__10__2_, connection_0__10__1_, 
        connection_0__10__0_, connection_0__8__31_, connection_0__8__30_, 
        connection_0__8__29_, connection_0__8__28_, connection_0__8__27_, 
        connection_0__8__26_, connection_0__8__25_, connection_0__8__24_, 
        connection_0__8__23_, connection_0__8__22_, connection_0__8__21_, 
        connection_0__8__20_, connection_0__8__19_, connection_0__8__18_, 
        connection_0__8__17_, connection_0__8__16_, connection_0__8__15_, 
        connection_0__8__14_, connection_0__8__13_, connection_0__8__12_, 
        connection_0__8__11_, connection_0__8__10_, connection_0__8__9_, 
        connection_0__8__8_, connection_0__8__7_, connection_0__8__6_, 
        connection_0__8__5_, connection_0__8__4_, connection_0__8__3_, 
        connection_0__8__2_, connection_0__8__1_, connection_0__8__0_}), 
        .o_valid({connection_valid_1__5_, connection_valid_1__4_}), 
        .o_data_bus({connection_1__5__31_, connection_1__5__30_, 
        connection_1__5__29_, connection_1__5__28_, connection_1__5__27_, 
        connection_1__5__26_, connection_1__5__25_, connection_1__5__24_, 
        connection_1__5__23_, connection_1__5__22_, connection_1__5__21_, 
        connection_1__5__20_, connection_1__5__19_, connection_1__5__18_, 
        connection_1__5__17_, connection_1__5__16_, connection_1__5__15_, 
        connection_1__5__14_, connection_1__5__13_, connection_1__5__12_, 
        connection_1__5__11_, connection_1__5__10_, connection_1__5__9_, 
        connection_1__5__8_, connection_1__5__7_, connection_1__5__6_, 
        connection_1__5__5_, connection_1__5__4_, connection_1__5__3_, 
        connection_1__5__2_, connection_1__5__1_, connection_1__5__0_, 
        connection_1__4__31_, connection_1__4__30_, connection_1__4__29_, 
        connection_1__4__28_, connection_1__4__27_, connection_1__4__26_, 
        connection_1__4__25_, connection_1__4__24_, connection_1__4__23_, 
        connection_1__4__22_, connection_1__4__21_, connection_1__4__20_, 
        connection_1__4__19_, connection_1__4__18_, connection_1__4__17_, 
        connection_1__4__16_, connection_1__4__15_, connection_1__4__14_, 
        connection_1__4__13_, connection_1__4__12_, connection_1__4__11_, 
        connection_1__4__10_, connection_1__4__9_, connection_1__4__8_, 
        connection_1__4__7_, connection_1__4__6_, connection_1__4__5_, 
        connection_1__4__4_, connection_1__4__3_, connection_1__4__2_, 
        connection_1__4__1_, connection_1__4__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[251:250]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_125 first_half_stages_0__group_first_half_0__switch_first_half_3__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__14_, 
        connection_valid_0__12_}), .i_data_bus({connection_0__14__31_, 
        connection_0__14__30_, connection_0__14__29_, connection_0__14__28_, 
        connection_0__14__27_, connection_0__14__26_, connection_0__14__25_, 
        connection_0__14__24_, connection_0__14__23_, connection_0__14__22_, 
        connection_0__14__21_, connection_0__14__20_, connection_0__14__19_, 
        connection_0__14__18_, connection_0__14__17_, connection_0__14__16_, 
        connection_0__14__15_, connection_0__14__14_, connection_0__14__13_, 
        connection_0__14__12_, connection_0__14__11_, connection_0__14__10_, 
        connection_0__14__9_, connection_0__14__8_, connection_0__14__7_, 
        connection_0__14__6_, connection_0__14__5_, connection_0__14__4_, 
        connection_0__14__3_, connection_0__14__2_, connection_0__14__1_, 
        connection_0__14__0_, connection_0__12__31_, connection_0__12__30_, 
        connection_0__12__29_, connection_0__12__28_, connection_0__12__27_, 
        connection_0__12__26_, connection_0__12__25_, connection_0__12__24_, 
        connection_0__12__23_, connection_0__12__22_, connection_0__12__21_, 
        connection_0__12__20_, connection_0__12__19_, connection_0__12__18_, 
        connection_0__12__17_, connection_0__12__16_, connection_0__12__15_, 
        connection_0__12__14_, connection_0__12__13_, connection_0__12__12_, 
        connection_0__12__11_, connection_0__12__10_, connection_0__12__9_, 
        connection_0__12__8_, connection_0__12__7_, connection_0__12__6_, 
        connection_0__12__5_, connection_0__12__4_, connection_0__12__3_, 
        connection_0__12__2_, connection_0__12__1_, connection_0__12__0_}), 
        .o_valid({connection_valid_1__7_, connection_valid_1__6_}), 
        .o_data_bus({connection_1__7__31_, connection_1__7__30_, 
        connection_1__7__29_, connection_1__7__28_, connection_1__7__27_, 
        connection_1__7__26_, connection_1__7__25_, connection_1__7__24_, 
        connection_1__7__23_, connection_1__7__22_, connection_1__7__21_, 
        connection_1__7__20_, connection_1__7__19_, connection_1__7__18_, 
        connection_1__7__17_, connection_1__7__16_, connection_1__7__15_, 
        connection_1__7__14_, connection_1__7__13_, connection_1__7__12_, 
        connection_1__7__11_, connection_1__7__10_, connection_1__7__9_, 
        connection_1__7__8_, connection_1__7__7_, connection_1__7__6_, 
        connection_1__7__5_, connection_1__7__4_, connection_1__7__3_, 
        connection_1__7__2_, connection_1__7__1_, connection_1__7__0_, 
        connection_1__6__31_, connection_1__6__30_, connection_1__6__29_, 
        connection_1__6__28_, connection_1__6__27_, connection_1__6__26_, 
        connection_1__6__25_, connection_1__6__24_, connection_1__6__23_, 
        connection_1__6__22_, connection_1__6__21_, connection_1__6__20_, 
        connection_1__6__19_, connection_1__6__18_, connection_1__6__17_, 
        connection_1__6__16_, connection_1__6__15_, connection_1__6__14_, 
        connection_1__6__13_, connection_1__6__12_, connection_1__6__11_, 
        connection_1__6__10_, connection_1__6__9_, connection_1__6__8_, 
        connection_1__6__7_, connection_1__6__6_, connection_1__6__5_, 
        connection_1__6__4_, connection_1__6__3_, connection_1__6__2_, 
        connection_1__6__1_, connection_1__6__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[249:248]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_124 first_half_stages_0__group_first_half_0__switch_first_half_4__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__18_, 
        connection_valid_0__16_}), .i_data_bus({connection_0__18__31_, 
        connection_0__18__30_, connection_0__18__29_, connection_0__18__28_, 
        connection_0__18__27_, connection_0__18__26_, connection_0__18__25_, 
        connection_0__18__24_, connection_0__18__23_, connection_0__18__22_, 
        connection_0__18__21_, connection_0__18__20_, connection_0__18__19_, 
        connection_0__18__18_, connection_0__18__17_, connection_0__18__16_, 
        connection_0__18__15_, connection_0__18__14_, connection_0__18__13_, 
        connection_0__18__12_, connection_0__18__11_, connection_0__18__10_, 
        connection_0__18__9_, connection_0__18__8_, connection_0__18__7_, 
        connection_0__18__6_, connection_0__18__5_, connection_0__18__4_, 
        connection_0__18__3_, connection_0__18__2_, connection_0__18__1_, 
        connection_0__18__0_, connection_0__16__31_, connection_0__16__30_, 
        connection_0__16__29_, connection_0__16__28_, connection_0__16__27_, 
        connection_0__16__26_, connection_0__16__25_, connection_0__16__24_, 
        connection_0__16__23_, connection_0__16__22_, connection_0__16__21_, 
        connection_0__16__20_, connection_0__16__19_, connection_0__16__18_, 
        connection_0__16__17_, connection_0__16__16_, connection_0__16__15_, 
        connection_0__16__14_, connection_0__16__13_, connection_0__16__12_, 
        connection_0__16__11_, connection_0__16__10_, connection_0__16__9_, 
        connection_0__16__8_, connection_0__16__7_, connection_0__16__6_, 
        connection_0__16__5_, connection_0__16__4_, connection_0__16__3_, 
        connection_0__16__2_, connection_0__16__1_, connection_0__16__0_}), 
        .o_valid({connection_valid_1__9_, connection_valid_1__8_}), 
        .o_data_bus({connection_1__9__31_, connection_1__9__30_, 
        connection_1__9__29_, connection_1__9__28_, connection_1__9__27_, 
        connection_1__9__26_, connection_1__9__25_, connection_1__9__24_, 
        connection_1__9__23_, connection_1__9__22_, connection_1__9__21_, 
        connection_1__9__20_, connection_1__9__19_, connection_1__9__18_, 
        connection_1__9__17_, connection_1__9__16_, connection_1__9__15_, 
        connection_1__9__14_, connection_1__9__13_, connection_1__9__12_, 
        connection_1__9__11_, connection_1__9__10_, connection_1__9__9_, 
        connection_1__9__8_, connection_1__9__7_, connection_1__9__6_, 
        connection_1__9__5_, connection_1__9__4_, connection_1__9__3_, 
        connection_1__9__2_, connection_1__9__1_, connection_1__9__0_, 
        connection_1__8__31_, connection_1__8__30_, connection_1__8__29_, 
        connection_1__8__28_, connection_1__8__27_, connection_1__8__26_, 
        connection_1__8__25_, connection_1__8__24_, connection_1__8__23_, 
        connection_1__8__22_, connection_1__8__21_, connection_1__8__20_, 
        connection_1__8__19_, connection_1__8__18_, connection_1__8__17_, 
        connection_1__8__16_, connection_1__8__15_, connection_1__8__14_, 
        connection_1__8__13_, connection_1__8__12_, connection_1__8__11_, 
        connection_1__8__10_, connection_1__8__9_, connection_1__8__8_, 
        connection_1__8__7_, connection_1__8__6_, connection_1__8__5_, 
        connection_1__8__4_, connection_1__8__3_, connection_1__8__2_, 
        connection_1__8__1_, connection_1__8__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[247:246]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_123 first_half_stages_0__group_first_half_0__switch_first_half_5__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__22_, 
        connection_valid_0__20_}), .i_data_bus({connection_0__22__31_, 
        connection_0__22__30_, connection_0__22__29_, connection_0__22__28_, 
        connection_0__22__27_, connection_0__22__26_, connection_0__22__25_, 
        connection_0__22__24_, connection_0__22__23_, connection_0__22__22_, 
        connection_0__22__21_, connection_0__22__20_, connection_0__22__19_, 
        connection_0__22__18_, connection_0__22__17_, connection_0__22__16_, 
        connection_0__22__15_, connection_0__22__14_, connection_0__22__13_, 
        connection_0__22__12_, connection_0__22__11_, connection_0__22__10_, 
        connection_0__22__9_, connection_0__22__8_, connection_0__22__7_, 
        connection_0__22__6_, connection_0__22__5_, connection_0__22__4_, 
        connection_0__22__3_, connection_0__22__2_, connection_0__22__1_, 
        connection_0__22__0_, connection_0__20__31_, connection_0__20__30_, 
        connection_0__20__29_, connection_0__20__28_, connection_0__20__27_, 
        connection_0__20__26_, connection_0__20__25_, connection_0__20__24_, 
        connection_0__20__23_, connection_0__20__22_, connection_0__20__21_, 
        connection_0__20__20_, connection_0__20__19_, connection_0__20__18_, 
        connection_0__20__17_, connection_0__20__16_, connection_0__20__15_, 
        connection_0__20__14_, connection_0__20__13_, connection_0__20__12_, 
        connection_0__20__11_, connection_0__20__10_, connection_0__20__9_, 
        connection_0__20__8_, connection_0__20__7_, connection_0__20__6_, 
        connection_0__20__5_, connection_0__20__4_, connection_0__20__3_, 
        connection_0__20__2_, connection_0__20__1_, connection_0__20__0_}), 
        .o_valid({connection_valid_1__11_, connection_valid_1__10_}), 
        .o_data_bus({connection_1__11__31_, connection_1__11__30_, 
        connection_1__11__29_, connection_1__11__28_, connection_1__11__27_, 
        connection_1__11__26_, connection_1__11__25_, connection_1__11__24_, 
        connection_1__11__23_, connection_1__11__22_, connection_1__11__21_, 
        connection_1__11__20_, connection_1__11__19_, connection_1__11__18_, 
        connection_1__11__17_, connection_1__11__16_, connection_1__11__15_, 
        connection_1__11__14_, connection_1__11__13_, connection_1__11__12_, 
        connection_1__11__11_, connection_1__11__10_, connection_1__11__9_, 
        connection_1__11__8_, connection_1__11__7_, connection_1__11__6_, 
        connection_1__11__5_, connection_1__11__4_, connection_1__11__3_, 
        connection_1__11__2_, connection_1__11__1_, connection_1__11__0_, 
        connection_1__10__31_, connection_1__10__30_, connection_1__10__29_, 
        connection_1__10__28_, connection_1__10__27_, connection_1__10__26_, 
        connection_1__10__25_, connection_1__10__24_, connection_1__10__23_, 
        connection_1__10__22_, connection_1__10__21_, connection_1__10__20_, 
        connection_1__10__19_, connection_1__10__18_, connection_1__10__17_, 
        connection_1__10__16_, connection_1__10__15_, connection_1__10__14_, 
        connection_1__10__13_, connection_1__10__12_, connection_1__10__11_, 
        connection_1__10__10_, connection_1__10__9_, connection_1__10__8_, 
        connection_1__10__7_, connection_1__10__6_, connection_1__10__5_, 
        connection_1__10__4_, connection_1__10__3_, connection_1__10__2_, 
        connection_1__10__1_, connection_1__10__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[245:244]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_122 first_half_stages_0__group_first_half_0__switch_first_half_6__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__26_, 
        connection_valid_0__24_}), .i_data_bus({connection_0__26__31_, 
        connection_0__26__30_, connection_0__26__29_, connection_0__26__28_, 
        connection_0__26__27_, connection_0__26__26_, connection_0__26__25_, 
        connection_0__26__24_, connection_0__26__23_, connection_0__26__22_, 
        connection_0__26__21_, connection_0__26__20_, connection_0__26__19_, 
        connection_0__26__18_, connection_0__26__17_, connection_0__26__16_, 
        connection_0__26__15_, connection_0__26__14_, connection_0__26__13_, 
        connection_0__26__12_, connection_0__26__11_, connection_0__26__10_, 
        connection_0__26__9_, connection_0__26__8_, connection_0__26__7_, 
        connection_0__26__6_, connection_0__26__5_, connection_0__26__4_, 
        connection_0__26__3_, connection_0__26__2_, connection_0__26__1_, 
        connection_0__26__0_, connection_0__24__31_, connection_0__24__30_, 
        connection_0__24__29_, connection_0__24__28_, connection_0__24__27_, 
        connection_0__24__26_, connection_0__24__25_, connection_0__24__24_, 
        connection_0__24__23_, connection_0__24__22_, connection_0__24__21_, 
        connection_0__24__20_, connection_0__24__19_, connection_0__24__18_, 
        connection_0__24__17_, connection_0__24__16_, connection_0__24__15_, 
        connection_0__24__14_, connection_0__24__13_, connection_0__24__12_, 
        connection_0__24__11_, connection_0__24__10_, connection_0__24__9_, 
        connection_0__24__8_, connection_0__24__7_, connection_0__24__6_, 
        connection_0__24__5_, connection_0__24__4_, connection_0__24__3_, 
        connection_0__24__2_, connection_0__24__1_, connection_0__24__0_}), 
        .o_valid({connection_valid_1__13_, connection_valid_1__12_}), 
        .o_data_bus({connection_1__13__31_, connection_1__13__30_, 
        connection_1__13__29_, connection_1__13__28_, connection_1__13__27_, 
        connection_1__13__26_, connection_1__13__25_, connection_1__13__24_, 
        connection_1__13__23_, connection_1__13__22_, connection_1__13__21_, 
        connection_1__13__20_, connection_1__13__19_, connection_1__13__18_, 
        connection_1__13__17_, connection_1__13__16_, connection_1__13__15_, 
        connection_1__13__14_, connection_1__13__13_, connection_1__13__12_, 
        connection_1__13__11_, connection_1__13__10_, connection_1__13__9_, 
        connection_1__13__8_, connection_1__13__7_, connection_1__13__6_, 
        connection_1__13__5_, connection_1__13__4_, connection_1__13__3_, 
        connection_1__13__2_, connection_1__13__1_, connection_1__13__0_, 
        connection_1__12__31_, connection_1__12__30_, connection_1__12__29_, 
        connection_1__12__28_, connection_1__12__27_, connection_1__12__26_, 
        connection_1__12__25_, connection_1__12__24_, connection_1__12__23_, 
        connection_1__12__22_, connection_1__12__21_, connection_1__12__20_, 
        connection_1__12__19_, connection_1__12__18_, connection_1__12__17_, 
        connection_1__12__16_, connection_1__12__15_, connection_1__12__14_, 
        connection_1__12__13_, connection_1__12__12_, connection_1__12__11_, 
        connection_1__12__10_, connection_1__12__9_, connection_1__12__8_, 
        connection_1__12__7_, connection_1__12__6_, connection_1__12__5_, 
        connection_1__12__4_, connection_1__12__3_, connection_1__12__2_, 
        connection_1__12__1_, connection_1__12__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[243:242]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_121 first_half_stages_0__group_first_half_0__switch_first_half_7__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__30_, 
        connection_valid_0__28_}), .i_data_bus({connection_0__30__31_, 
        connection_0__30__30_, connection_0__30__29_, connection_0__30__28_, 
        connection_0__30__27_, connection_0__30__26_, connection_0__30__25_, 
        connection_0__30__24_, connection_0__30__23_, connection_0__30__22_, 
        connection_0__30__21_, connection_0__30__20_, connection_0__30__19_, 
        connection_0__30__18_, connection_0__30__17_, connection_0__30__16_, 
        connection_0__30__15_, connection_0__30__14_, connection_0__30__13_, 
        connection_0__30__12_, connection_0__30__11_, connection_0__30__10_, 
        connection_0__30__9_, connection_0__30__8_, connection_0__30__7_, 
        connection_0__30__6_, connection_0__30__5_, connection_0__30__4_, 
        connection_0__30__3_, connection_0__30__2_, connection_0__30__1_, 
        connection_0__30__0_, connection_0__28__31_, connection_0__28__30_, 
        connection_0__28__29_, connection_0__28__28_, connection_0__28__27_, 
        connection_0__28__26_, connection_0__28__25_, connection_0__28__24_, 
        connection_0__28__23_, connection_0__28__22_, connection_0__28__21_, 
        connection_0__28__20_, connection_0__28__19_, connection_0__28__18_, 
        connection_0__28__17_, connection_0__28__16_, connection_0__28__15_, 
        connection_0__28__14_, connection_0__28__13_, connection_0__28__12_, 
        connection_0__28__11_, connection_0__28__10_, connection_0__28__9_, 
        connection_0__28__8_, connection_0__28__7_, connection_0__28__6_, 
        connection_0__28__5_, connection_0__28__4_, connection_0__28__3_, 
        connection_0__28__2_, connection_0__28__1_, connection_0__28__0_}), 
        .o_valid({connection_valid_1__15_, connection_valid_1__14_}), 
        .o_data_bus({connection_1__15__31_, connection_1__15__30_, 
        connection_1__15__29_, connection_1__15__28_, connection_1__15__27_, 
        connection_1__15__26_, connection_1__15__25_, connection_1__15__24_, 
        connection_1__15__23_, connection_1__15__22_, connection_1__15__21_, 
        connection_1__15__20_, connection_1__15__19_, connection_1__15__18_, 
        connection_1__15__17_, connection_1__15__16_, connection_1__15__15_, 
        connection_1__15__14_, connection_1__15__13_, connection_1__15__12_, 
        connection_1__15__11_, connection_1__15__10_, connection_1__15__9_, 
        connection_1__15__8_, connection_1__15__7_, connection_1__15__6_, 
        connection_1__15__5_, connection_1__15__4_, connection_1__15__3_, 
        connection_1__15__2_, connection_1__15__1_, connection_1__15__0_, 
        connection_1__14__31_, connection_1__14__30_, connection_1__14__29_, 
        connection_1__14__28_, connection_1__14__27_, connection_1__14__26_, 
        connection_1__14__25_, connection_1__14__24_, connection_1__14__23_, 
        connection_1__14__22_, connection_1__14__21_, connection_1__14__20_, 
        connection_1__14__19_, connection_1__14__18_, connection_1__14__17_, 
        connection_1__14__16_, connection_1__14__15_, connection_1__14__14_, 
        connection_1__14__13_, connection_1__14__12_, connection_1__14__11_, 
        connection_1__14__10_, connection_1__14__9_, connection_1__14__8_, 
        connection_1__14__7_, connection_1__14__6_, connection_1__14__5_, 
        connection_1__14__4_, connection_1__14__3_, connection_1__14__2_, 
        connection_1__14__1_, connection_1__14__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[241:240]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_120 first_half_stages_0__group_first_half_0__switch_first_half_8__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__3_, 
        connection_valid_0__1_}), .i_data_bus({connection_0__3__31_, 
        connection_0__3__30_, connection_0__3__29_, connection_0__3__28_, 
        connection_0__3__27_, connection_0__3__26_, connection_0__3__25_, 
        connection_0__3__24_, connection_0__3__23_, connection_0__3__22_, 
        connection_0__3__21_, connection_0__3__20_, connection_0__3__19_, 
        connection_0__3__18_, connection_0__3__17_, connection_0__3__16_, 
        connection_0__3__15_, connection_0__3__14_, connection_0__3__13_, 
        connection_0__3__12_, connection_0__3__11_, connection_0__3__10_, 
        connection_0__3__9_, connection_0__3__8_, connection_0__3__7_, 
        connection_0__3__6_, connection_0__3__5_, connection_0__3__4_, 
        connection_0__3__3_, connection_0__3__2_, connection_0__3__1_, 
        connection_0__3__0_, connection_0__1__31_, connection_0__1__30_, 
        connection_0__1__29_, connection_0__1__28_, connection_0__1__27_, 
        connection_0__1__26_, connection_0__1__25_, connection_0__1__24_, 
        connection_0__1__23_, connection_0__1__22_, connection_0__1__21_, 
        connection_0__1__20_, connection_0__1__19_, connection_0__1__18_, 
        connection_0__1__17_, connection_0__1__16_, connection_0__1__15_, 
        connection_0__1__14_, connection_0__1__13_, connection_0__1__12_, 
        connection_0__1__11_, connection_0__1__10_, connection_0__1__9_, 
        connection_0__1__8_, connection_0__1__7_, connection_0__1__6_, 
        connection_0__1__5_, connection_0__1__4_, connection_0__1__3_, 
        connection_0__1__2_, connection_0__1__1_, connection_0__1__0_}), 
        .o_valid({connection_valid_1__17_, connection_valid_1__16_}), 
        .o_data_bus({connection_1__17__31_, connection_1__17__30_, 
        connection_1__17__29_, connection_1__17__28_, connection_1__17__27_, 
        connection_1__17__26_, connection_1__17__25_, connection_1__17__24_, 
        connection_1__17__23_, connection_1__17__22_, connection_1__17__21_, 
        connection_1__17__20_, connection_1__17__19_, connection_1__17__18_, 
        connection_1__17__17_, connection_1__17__16_, connection_1__17__15_, 
        connection_1__17__14_, connection_1__17__13_, connection_1__17__12_, 
        connection_1__17__11_, connection_1__17__10_, connection_1__17__9_, 
        connection_1__17__8_, connection_1__17__7_, connection_1__17__6_, 
        connection_1__17__5_, connection_1__17__4_, connection_1__17__3_, 
        connection_1__17__2_, connection_1__17__1_, connection_1__17__0_, 
        connection_1__16__31_, connection_1__16__30_, connection_1__16__29_, 
        connection_1__16__28_, connection_1__16__27_, connection_1__16__26_, 
        connection_1__16__25_, connection_1__16__24_, connection_1__16__23_, 
        connection_1__16__22_, connection_1__16__21_, connection_1__16__20_, 
        connection_1__16__19_, connection_1__16__18_, connection_1__16__17_, 
        connection_1__16__16_, connection_1__16__15_, connection_1__16__14_, 
        connection_1__16__13_, connection_1__16__12_, connection_1__16__11_, 
        connection_1__16__10_, connection_1__16__9_, connection_1__16__8_, 
        connection_1__16__7_, connection_1__16__6_, connection_1__16__5_, 
        connection_1__16__4_, connection_1__16__3_, connection_1__16__2_, 
        connection_1__16__1_, connection_1__16__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[239:238]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_119 first_half_stages_0__group_first_half_0__switch_first_half_9__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__7_, 
        connection_valid_0__5_}), .i_data_bus({connection_0__7__31_, 
        connection_0__7__30_, connection_0__7__29_, connection_0__7__28_, 
        connection_0__7__27_, connection_0__7__26_, connection_0__7__25_, 
        connection_0__7__24_, connection_0__7__23_, connection_0__7__22_, 
        connection_0__7__21_, connection_0__7__20_, connection_0__7__19_, 
        connection_0__7__18_, connection_0__7__17_, connection_0__7__16_, 
        connection_0__7__15_, connection_0__7__14_, connection_0__7__13_, 
        connection_0__7__12_, connection_0__7__11_, connection_0__7__10_, 
        connection_0__7__9_, connection_0__7__8_, connection_0__7__7_, 
        connection_0__7__6_, connection_0__7__5_, connection_0__7__4_, 
        connection_0__7__3_, connection_0__7__2_, connection_0__7__1_, 
        connection_0__7__0_, connection_0__5__31_, connection_0__5__30_, 
        connection_0__5__29_, connection_0__5__28_, connection_0__5__27_, 
        connection_0__5__26_, connection_0__5__25_, connection_0__5__24_, 
        connection_0__5__23_, connection_0__5__22_, connection_0__5__21_, 
        connection_0__5__20_, connection_0__5__19_, connection_0__5__18_, 
        connection_0__5__17_, connection_0__5__16_, connection_0__5__15_, 
        connection_0__5__14_, connection_0__5__13_, connection_0__5__12_, 
        connection_0__5__11_, connection_0__5__10_, connection_0__5__9_, 
        connection_0__5__8_, connection_0__5__7_, connection_0__5__6_, 
        connection_0__5__5_, connection_0__5__4_, connection_0__5__3_, 
        connection_0__5__2_, connection_0__5__1_, connection_0__5__0_}), 
        .o_valid({connection_valid_1__19_, connection_valid_1__18_}), 
        .o_data_bus({connection_1__19__31_, connection_1__19__30_, 
        connection_1__19__29_, connection_1__19__28_, connection_1__19__27_, 
        connection_1__19__26_, connection_1__19__25_, connection_1__19__24_, 
        connection_1__19__23_, connection_1__19__22_, connection_1__19__21_, 
        connection_1__19__20_, connection_1__19__19_, connection_1__19__18_, 
        connection_1__19__17_, connection_1__19__16_, connection_1__19__15_, 
        connection_1__19__14_, connection_1__19__13_, connection_1__19__12_, 
        connection_1__19__11_, connection_1__19__10_, connection_1__19__9_, 
        connection_1__19__8_, connection_1__19__7_, connection_1__19__6_, 
        connection_1__19__5_, connection_1__19__4_, connection_1__19__3_, 
        connection_1__19__2_, connection_1__19__1_, connection_1__19__0_, 
        connection_1__18__31_, connection_1__18__30_, connection_1__18__29_, 
        connection_1__18__28_, connection_1__18__27_, connection_1__18__26_, 
        connection_1__18__25_, connection_1__18__24_, connection_1__18__23_, 
        connection_1__18__22_, connection_1__18__21_, connection_1__18__20_, 
        connection_1__18__19_, connection_1__18__18_, connection_1__18__17_, 
        connection_1__18__16_, connection_1__18__15_, connection_1__18__14_, 
        connection_1__18__13_, connection_1__18__12_, connection_1__18__11_, 
        connection_1__18__10_, connection_1__18__9_, connection_1__18__8_, 
        connection_1__18__7_, connection_1__18__6_, connection_1__18__5_, 
        connection_1__18__4_, connection_1__18__3_, connection_1__18__2_, 
        connection_1__18__1_, connection_1__18__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[237:236]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_118 first_half_stages_0__group_first_half_0__switch_first_half_10__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__11_, 
        connection_valid_0__9_}), .i_data_bus({connection_0__11__31_, 
        connection_0__11__30_, connection_0__11__29_, connection_0__11__28_, 
        connection_0__11__27_, connection_0__11__26_, connection_0__11__25_, 
        connection_0__11__24_, connection_0__11__23_, connection_0__11__22_, 
        connection_0__11__21_, connection_0__11__20_, connection_0__11__19_, 
        connection_0__11__18_, connection_0__11__17_, connection_0__11__16_, 
        connection_0__11__15_, connection_0__11__14_, connection_0__11__13_, 
        connection_0__11__12_, connection_0__11__11_, connection_0__11__10_, 
        connection_0__11__9_, connection_0__11__8_, connection_0__11__7_, 
        connection_0__11__6_, connection_0__11__5_, connection_0__11__4_, 
        connection_0__11__3_, connection_0__11__2_, connection_0__11__1_, 
        connection_0__11__0_, connection_0__9__31_, connection_0__9__30_, 
        connection_0__9__29_, connection_0__9__28_, connection_0__9__27_, 
        connection_0__9__26_, connection_0__9__25_, connection_0__9__24_, 
        connection_0__9__23_, connection_0__9__22_, connection_0__9__21_, 
        connection_0__9__20_, connection_0__9__19_, connection_0__9__18_, 
        connection_0__9__17_, connection_0__9__16_, connection_0__9__15_, 
        connection_0__9__14_, connection_0__9__13_, connection_0__9__12_, 
        connection_0__9__11_, connection_0__9__10_, connection_0__9__9_, 
        connection_0__9__8_, connection_0__9__7_, connection_0__9__6_, 
        connection_0__9__5_, connection_0__9__4_, connection_0__9__3_, 
        connection_0__9__2_, connection_0__9__1_, connection_0__9__0_}), 
        .o_valid({connection_valid_1__21_, connection_valid_1__20_}), 
        .o_data_bus({connection_1__21__31_, connection_1__21__30_, 
        connection_1__21__29_, connection_1__21__28_, connection_1__21__27_, 
        connection_1__21__26_, connection_1__21__25_, connection_1__21__24_, 
        connection_1__21__23_, connection_1__21__22_, connection_1__21__21_, 
        connection_1__21__20_, connection_1__21__19_, connection_1__21__18_, 
        connection_1__21__17_, connection_1__21__16_, connection_1__21__15_, 
        connection_1__21__14_, connection_1__21__13_, connection_1__21__12_, 
        connection_1__21__11_, connection_1__21__10_, connection_1__21__9_, 
        connection_1__21__8_, connection_1__21__7_, connection_1__21__6_, 
        connection_1__21__5_, connection_1__21__4_, connection_1__21__3_, 
        connection_1__21__2_, connection_1__21__1_, connection_1__21__0_, 
        connection_1__20__31_, connection_1__20__30_, connection_1__20__29_, 
        connection_1__20__28_, connection_1__20__27_, connection_1__20__26_, 
        connection_1__20__25_, connection_1__20__24_, connection_1__20__23_, 
        connection_1__20__22_, connection_1__20__21_, connection_1__20__20_, 
        connection_1__20__19_, connection_1__20__18_, connection_1__20__17_, 
        connection_1__20__16_, connection_1__20__15_, connection_1__20__14_, 
        connection_1__20__13_, connection_1__20__12_, connection_1__20__11_, 
        connection_1__20__10_, connection_1__20__9_, connection_1__20__8_, 
        connection_1__20__7_, connection_1__20__6_, connection_1__20__5_, 
        connection_1__20__4_, connection_1__20__3_, connection_1__20__2_, 
        connection_1__20__1_, connection_1__20__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[235:234]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_117 first_half_stages_0__group_first_half_0__switch_first_half_11__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__15_, 
        connection_valid_0__13_}), .i_data_bus({connection_0__15__31_, 
        connection_0__15__30_, connection_0__15__29_, connection_0__15__28_, 
        connection_0__15__27_, connection_0__15__26_, connection_0__15__25_, 
        connection_0__15__24_, connection_0__15__23_, connection_0__15__22_, 
        connection_0__15__21_, connection_0__15__20_, connection_0__15__19_, 
        connection_0__15__18_, connection_0__15__17_, connection_0__15__16_, 
        connection_0__15__15_, connection_0__15__14_, connection_0__15__13_, 
        connection_0__15__12_, connection_0__15__11_, connection_0__15__10_, 
        connection_0__15__9_, connection_0__15__8_, connection_0__15__7_, 
        connection_0__15__6_, connection_0__15__5_, connection_0__15__4_, 
        connection_0__15__3_, connection_0__15__2_, connection_0__15__1_, 
        connection_0__15__0_, connection_0__13__31_, connection_0__13__30_, 
        connection_0__13__29_, connection_0__13__28_, connection_0__13__27_, 
        connection_0__13__26_, connection_0__13__25_, connection_0__13__24_, 
        connection_0__13__23_, connection_0__13__22_, connection_0__13__21_, 
        connection_0__13__20_, connection_0__13__19_, connection_0__13__18_, 
        connection_0__13__17_, connection_0__13__16_, connection_0__13__15_, 
        connection_0__13__14_, connection_0__13__13_, connection_0__13__12_, 
        connection_0__13__11_, connection_0__13__10_, connection_0__13__9_, 
        connection_0__13__8_, connection_0__13__7_, connection_0__13__6_, 
        connection_0__13__5_, connection_0__13__4_, connection_0__13__3_, 
        connection_0__13__2_, connection_0__13__1_, connection_0__13__0_}), 
        .o_valid({connection_valid_1__23_, connection_valid_1__22_}), 
        .o_data_bus({connection_1__23__31_, connection_1__23__30_, 
        connection_1__23__29_, connection_1__23__28_, connection_1__23__27_, 
        connection_1__23__26_, connection_1__23__25_, connection_1__23__24_, 
        connection_1__23__23_, connection_1__23__22_, connection_1__23__21_, 
        connection_1__23__20_, connection_1__23__19_, connection_1__23__18_, 
        connection_1__23__17_, connection_1__23__16_, connection_1__23__15_, 
        connection_1__23__14_, connection_1__23__13_, connection_1__23__12_, 
        connection_1__23__11_, connection_1__23__10_, connection_1__23__9_, 
        connection_1__23__8_, connection_1__23__7_, connection_1__23__6_, 
        connection_1__23__5_, connection_1__23__4_, connection_1__23__3_, 
        connection_1__23__2_, connection_1__23__1_, connection_1__23__0_, 
        connection_1__22__31_, connection_1__22__30_, connection_1__22__29_, 
        connection_1__22__28_, connection_1__22__27_, connection_1__22__26_, 
        connection_1__22__25_, connection_1__22__24_, connection_1__22__23_, 
        connection_1__22__22_, connection_1__22__21_, connection_1__22__20_, 
        connection_1__22__19_, connection_1__22__18_, connection_1__22__17_, 
        connection_1__22__16_, connection_1__22__15_, connection_1__22__14_, 
        connection_1__22__13_, connection_1__22__12_, connection_1__22__11_, 
        connection_1__22__10_, connection_1__22__9_, connection_1__22__8_, 
        connection_1__22__7_, connection_1__22__6_, connection_1__22__5_, 
        connection_1__22__4_, connection_1__22__3_, connection_1__22__2_, 
        connection_1__22__1_, connection_1__22__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[233:232]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_116 first_half_stages_0__group_first_half_0__switch_first_half_12__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__19_, 
        connection_valid_0__17_}), .i_data_bus({connection_0__19__31_, 
        connection_0__19__30_, connection_0__19__29_, connection_0__19__28_, 
        connection_0__19__27_, connection_0__19__26_, connection_0__19__25_, 
        connection_0__19__24_, connection_0__19__23_, connection_0__19__22_, 
        connection_0__19__21_, connection_0__19__20_, connection_0__19__19_, 
        connection_0__19__18_, connection_0__19__17_, connection_0__19__16_, 
        connection_0__19__15_, connection_0__19__14_, connection_0__19__13_, 
        connection_0__19__12_, connection_0__19__11_, connection_0__19__10_, 
        connection_0__19__9_, connection_0__19__8_, connection_0__19__7_, 
        connection_0__19__6_, connection_0__19__5_, connection_0__19__4_, 
        connection_0__19__3_, connection_0__19__2_, connection_0__19__1_, 
        connection_0__19__0_, connection_0__17__31_, connection_0__17__30_, 
        connection_0__17__29_, connection_0__17__28_, connection_0__17__27_, 
        connection_0__17__26_, connection_0__17__25_, connection_0__17__24_, 
        connection_0__17__23_, connection_0__17__22_, connection_0__17__21_, 
        connection_0__17__20_, connection_0__17__19_, connection_0__17__18_, 
        connection_0__17__17_, connection_0__17__16_, connection_0__17__15_, 
        connection_0__17__14_, connection_0__17__13_, connection_0__17__12_, 
        connection_0__17__11_, connection_0__17__10_, connection_0__17__9_, 
        connection_0__17__8_, connection_0__17__7_, connection_0__17__6_, 
        connection_0__17__5_, connection_0__17__4_, connection_0__17__3_, 
        connection_0__17__2_, connection_0__17__1_, connection_0__17__0_}), 
        .o_valid({connection_valid_1__25_, connection_valid_1__24_}), 
        .o_data_bus({connection_1__25__31_, connection_1__25__30_, 
        connection_1__25__29_, connection_1__25__28_, connection_1__25__27_, 
        connection_1__25__26_, connection_1__25__25_, connection_1__25__24_, 
        connection_1__25__23_, connection_1__25__22_, connection_1__25__21_, 
        connection_1__25__20_, connection_1__25__19_, connection_1__25__18_, 
        connection_1__25__17_, connection_1__25__16_, connection_1__25__15_, 
        connection_1__25__14_, connection_1__25__13_, connection_1__25__12_, 
        connection_1__25__11_, connection_1__25__10_, connection_1__25__9_, 
        connection_1__25__8_, connection_1__25__7_, connection_1__25__6_, 
        connection_1__25__5_, connection_1__25__4_, connection_1__25__3_, 
        connection_1__25__2_, connection_1__25__1_, connection_1__25__0_, 
        connection_1__24__31_, connection_1__24__30_, connection_1__24__29_, 
        connection_1__24__28_, connection_1__24__27_, connection_1__24__26_, 
        connection_1__24__25_, connection_1__24__24_, connection_1__24__23_, 
        connection_1__24__22_, connection_1__24__21_, connection_1__24__20_, 
        connection_1__24__19_, connection_1__24__18_, connection_1__24__17_, 
        connection_1__24__16_, connection_1__24__15_, connection_1__24__14_, 
        connection_1__24__13_, connection_1__24__12_, connection_1__24__11_, 
        connection_1__24__10_, connection_1__24__9_, connection_1__24__8_, 
        connection_1__24__7_, connection_1__24__6_, connection_1__24__5_, 
        connection_1__24__4_, connection_1__24__3_, connection_1__24__2_, 
        connection_1__24__1_, connection_1__24__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[231:230]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_115 first_half_stages_0__group_first_half_0__switch_first_half_13__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__23_, 
        connection_valid_0__21_}), .i_data_bus({connection_0__23__31_, 
        connection_0__23__30_, connection_0__23__29_, connection_0__23__28_, 
        connection_0__23__27_, connection_0__23__26_, connection_0__23__25_, 
        connection_0__23__24_, connection_0__23__23_, connection_0__23__22_, 
        connection_0__23__21_, connection_0__23__20_, connection_0__23__19_, 
        connection_0__23__18_, connection_0__23__17_, connection_0__23__16_, 
        connection_0__23__15_, connection_0__23__14_, connection_0__23__13_, 
        connection_0__23__12_, connection_0__23__11_, connection_0__23__10_, 
        connection_0__23__9_, connection_0__23__8_, connection_0__23__7_, 
        connection_0__23__6_, connection_0__23__5_, connection_0__23__4_, 
        connection_0__23__3_, connection_0__23__2_, connection_0__23__1_, 
        connection_0__23__0_, connection_0__21__31_, connection_0__21__30_, 
        connection_0__21__29_, connection_0__21__28_, connection_0__21__27_, 
        connection_0__21__26_, connection_0__21__25_, connection_0__21__24_, 
        connection_0__21__23_, connection_0__21__22_, connection_0__21__21_, 
        connection_0__21__20_, connection_0__21__19_, connection_0__21__18_, 
        connection_0__21__17_, connection_0__21__16_, connection_0__21__15_, 
        connection_0__21__14_, connection_0__21__13_, connection_0__21__12_, 
        connection_0__21__11_, connection_0__21__10_, connection_0__21__9_, 
        connection_0__21__8_, connection_0__21__7_, connection_0__21__6_, 
        connection_0__21__5_, connection_0__21__4_, connection_0__21__3_, 
        connection_0__21__2_, connection_0__21__1_, connection_0__21__0_}), 
        .o_valid({connection_valid_1__27_, connection_valid_1__26_}), 
        .o_data_bus({connection_1__27__31_, connection_1__27__30_, 
        connection_1__27__29_, connection_1__27__28_, connection_1__27__27_, 
        connection_1__27__26_, connection_1__27__25_, connection_1__27__24_, 
        connection_1__27__23_, connection_1__27__22_, connection_1__27__21_, 
        connection_1__27__20_, connection_1__27__19_, connection_1__27__18_, 
        connection_1__27__17_, connection_1__27__16_, connection_1__27__15_, 
        connection_1__27__14_, connection_1__27__13_, connection_1__27__12_, 
        connection_1__27__11_, connection_1__27__10_, connection_1__27__9_, 
        connection_1__27__8_, connection_1__27__7_, connection_1__27__6_, 
        connection_1__27__5_, connection_1__27__4_, connection_1__27__3_, 
        connection_1__27__2_, connection_1__27__1_, connection_1__27__0_, 
        connection_1__26__31_, connection_1__26__30_, connection_1__26__29_, 
        connection_1__26__28_, connection_1__26__27_, connection_1__26__26_, 
        connection_1__26__25_, connection_1__26__24_, connection_1__26__23_, 
        connection_1__26__22_, connection_1__26__21_, connection_1__26__20_, 
        connection_1__26__19_, connection_1__26__18_, connection_1__26__17_, 
        connection_1__26__16_, connection_1__26__15_, connection_1__26__14_, 
        connection_1__26__13_, connection_1__26__12_, connection_1__26__11_, 
        connection_1__26__10_, connection_1__26__9_, connection_1__26__8_, 
        connection_1__26__7_, connection_1__26__6_, connection_1__26__5_, 
        connection_1__26__4_, connection_1__26__3_, connection_1__26__2_, 
        connection_1__26__1_, connection_1__26__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[229:228]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_114 first_half_stages_0__group_first_half_0__switch_first_half_14__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__27_, 
        connection_valid_0__25_}), .i_data_bus({connection_0__27__31_, 
        connection_0__27__30_, connection_0__27__29_, connection_0__27__28_, 
        connection_0__27__27_, connection_0__27__26_, connection_0__27__25_, 
        connection_0__27__24_, connection_0__27__23_, connection_0__27__22_, 
        connection_0__27__21_, connection_0__27__20_, connection_0__27__19_, 
        connection_0__27__18_, connection_0__27__17_, connection_0__27__16_, 
        connection_0__27__15_, connection_0__27__14_, connection_0__27__13_, 
        connection_0__27__12_, connection_0__27__11_, connection_0__27__10_, 
        connection_0__27__9_, connection_0__27__8_, connection_0__27__7_, 
        connection_0__27__6_, connection_0__27__5_, connection_0__27__4_, 
        connection_0__27__3_, connection_0__27__2_, connection_0__27__1_, 
        connection_0__27__0_, connection_0__25__31_, connection_0__25__30_, 
        connection_0__25__29_, connection_0__25__28_, connection_0__25__27_, 
        connection_0__25__26_, connection_0__25__25_, connection_0__25__24_, 
        connection_0__25__23_, connection_0__25__22_, connection_0__25__21_, 
        connection_0__25__20_, connection_0__25__19_, connection_0__25__18_, 
        connection_0__25__17_, connection_0__25__16_, connection_0__25__15_, 
        connection_0__25__14_, connection_0__25__13_, connection_0__25__12_, 
        connection_0__25__11_, connection_0__25__10_, connection_0__25__9_, 
        connection_0__25__8_, connection_0__25__7_, connection_0__25__6_, 
        connection_0__25__5_, connection_0__25__4_, connection_0__25__3_, 
        connection_0__25__2_, connection_0__25__1_, connection_0__25__0_}), 
        .o_valid({connection_valid_1__29_, connection_valid_1__28_}), 
        .o_data_bus({connection_1__29__31_, connection_1__29__30_, 
        connection_1__29__29_, connection_1__29__28_, connection_1__29__27_, 
        connection_1__29__26_, connection_1__29__25_, connection_1__29__24_, 
        connection_1__29__23_, connection_1__29__22_, connection_1__29__21_, 
        connection_1__29__20_, connection_1__29__19_, connection_1__29__18_, 
        connection_1__29__17_, connection_1__29__16_, connection_1__29__15_, 
        connection_1__29__14_, connection_1__29__13_, connection_1__29__12_, 
        connection_1__29__11_, connection_1__29__10_, connection_1__29__9_, 
        connection_1__29__8_, connection_1__29__7_, connection_1__29__6_, 
        connection_1__29__5_, connection_1__29__4_, connection_1__29__3_, 
        connection_1__29__2_, connection_1__29__1_, connection_1__29__0_, 
        connection_1__28__31_, connection_1__28__30_, connection_1__28__29_, 
        connection_1__28__28_, connection_1__28__27_, connection_1__28__26_, 
        connection_1__28__25_, connection_1__28__24_, connection_1__28__23_, 
        connection_1__28__22_, connection_1__28__21_, connection_1__28__20_, 
        connection_1__28__19_, connection_1__28__18_, connection_1__28__17_, 
        connection_1__28__16_, connection_1__28__15_, connection_1__28__14_, 
        connection_1__28__13_, connection_1__28__12_, connection_1__28__11_, 
        connection_1__28__10_, connection_1__28__9_, connection_1__28__8_, 
        connection_1__28__7_, connection_1__28__6_, connection_1__28__5_, 
        connection_1__28__4_, connection_1__28__3_, connection_1__28__2_, 
        connection_1__28__1_, connection_1__28__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[227:226]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_113 first_half_stages_0__group_first_half_0__switch_first_half_15__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__31_, 
        connection_valid_0__29_}), .i_data_bus({connection_0__31__31_, 
        connection_0__31__30_, connection_0__31__29_, connection_0__31__28_, 
        connection_0__31__27_, connection_0__31__26_, connection_0__31__25_, 
        connection_0__31__24_, connection_0__31__23_, connection_0__31__22_, 
        connection_0__31__21_, connection_0__31__20_, connection_0__31__19_, 
        connection_0__31__18_, connection_0__31__17_, connection_0__31__16_, 
        connection_0__31__15_, connection_0__31__14_, connection_0__31__13_, 
        connection_0__31__12_, connection_0__31__11_, connection_0__31__10_, 
        connection_0__31__9_, connection_0__31__8_, connection_0__31__7_, 
        connection_0__31__6_, connection_0__31__5_, connection_0__31__4_, 
        connection_0__31__3_, connection_0__31__2_, connection_0__31__1_, 
        connection_0__31__0_, connection_0__29__31_, connection_0__29__30_, 
        connection_0__29__29_, connection_0__29__28_, connection_0__29__27_, 
        connection_0__29__26_, connection_0__29__25_, connection_0__29__24_, 
        connection_0__29__23_, connection_0__29__22_, connection_0__29__21_, 
        connection_0__29__20_, connection_0__29__19_, connection_0__29__18_, 
        connection_0__29__17_, connection_0__29__16_, connection_0__29__15_, 
        connection_0__29__14_, connection_0__29__13_, connection_0__29__12_, 
        connection_0__29__11_, connection_0__29__10_, connection_0__29__9_, 
        connection_0__29__8_, connection_0__29__7_, connection_0__29__6_, 
        connection_0__29__5_, connection_0__29__4_, connection_0__29__3_, 
        connection_0__29__2_, connection_0__29__1_, connection_0__29__0_}), 
        .o_valid({connection_valid_1__31_, connection_valid_1__30_}), 
        .o_data_bus({connection_1__31__31_, connection_1__31__30_, 
        connection_1__31__29_, connection_1__31__28_, connection_1__31__27_, 
        connection_1__31__26_, connection_1__31__25_, connection_1__31__24_, 
        connection_1__31__23_, connection_1__31__22_, connection_1__31__21_, 
        connection_1__31__20_, connection_1__31__19_, connection_1__31__18_, 
        connection_1__31__17_, connection_1__31__16_, connection_1__31__15_, 
        connection_1__31__14_, connection_1__31__13_, connection_1__31__12_, 
        connection_1__31__11_, connection_1__31__10_, connection_1__31__9_, 
        connection_1__31__8_, connection_1__31__7_, connection_1__31__6_, 
        connection_1__31__5_, connection_1__31__4_, connection_1__31__3_, 
        connection_1__31__2_, connection_1__31__1_, connection_1__31__0_, 
        connection_1__30__31_, connection_1__30__30_, connection_1__30__29_, 
        connection_1__30__28_, connection_1__30__27_, connection_1__30__26_, 
        connection_1__30__25_, connection_1__30__24_, connection_1__30__23_, 
        connection_1__30__22_, connection_1__30__21_, connection_1__30__20_, 
        connection_1__30__19_, connection_1__30__18_, connection_1__30__17_, 
        connection_1__30__16_, connection_1__30__15_, connection_1__30__14_, 
        connection_1__30__13_, connection_1__30__12_, connection_1__30__11_, 
        connection_1__30__10_, connection_1__30__9_, connection_1__30__8_, 
        connection_1__30__7_, connection_1__30__6_, connection_1__30__5_, 
        connection_1__30__4_, connection_1__30__3_, connection_1__30__2_, 
        connection_1__30__1_, connection_1__30__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[225:224]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_112 first_half_stages_1__group_first_half_0__switch_first_half_0__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_1__2_, 
        connection_valid_1__0_}), .i_data_bus({connection_1__2__31_, 
        connection_1__2__30_, connection_1__2__29_, connection_1__2__28_, 
        connection_1__2__27_, connection_1__2__26_, connection_1__2__25_, 
        connection_1__2__24_, connection_1__2__23_, connection_1__2__22_, 
        connection_1__2__21_, connection_1__2__20_, connection_1__2__19_, 
        connection_1__2__18_, connection_1__2__17_, connection_1__2__16_, 
        connection_1__2__15_, connection_1__2__14_, connection_1__2__13_, 
        connection_1__2__12_, connection_1__2__11_, connection_1__2__10_, 
        connection_1__2__9_, connection_1__2__8_, connection_1__2__7_, 
        connection_1__2__6_, connection_1__2__5_, connection_1__2__4_, 
        connection_1__2__3_, connection_1__2__2_, connection_1__2__1_, 
        connection_1__2__0_, connection_1__0__31_, connection_1__0__30_, 
        connection_1__0__29_, connection_1__0__28_, connection_1__0__27_, 
        connection_1__0__26_, connection_1__0__25_, connection_1__0__24_, 
        connection_1__0__23_, connection_1__0__22_, connection_1__0__21_, 
        connection_1__0__20_, connection_1__0__19_, connection_1__0__18_, 
        connection_1__0__17_, connection_1__0__16_, connection_1__0__15_, 
        connection_1__0__14_, connection_1__0__13_, connection_1__0__12_, 
        connection_1__0__11_, connection_1__0__10_, connection_1__0__9_, 
        connection_1__0__8_, connection_1__0__7_, connection_1__0__6_, 
        connection_1__0__5_, connection_1__0__4_, connection_1__0__3_, 
        connection_1__0__2_, connection_1__0__1_, connection_1__0__0_}), 
        .o_valid({connection_valid_2__1_, connection_valid_2__0_}), 
        .o_data_bus({connection_2__1__31_, connection_2__1__30_, 
        connection_2__1__29_, connection_2__1__28_, connection_2__1__27_, 
        connection_2__1__26_, connection_2__1__25_, connection_2__1__24_, 
        connection_2__1__23_, connection_2__1__22_, connection_2__1__21_, 
        connection_2__1__20_, connection_2__1__19_, connection_2__1__18_, 
        connection_2__1__17_, connection_2__1__16_, connection_2__1__15_, 
        connection_2__1__14_, connection_2__1__13_, connection_2__1__12_, 
        connection_2__1__11_, connection_2__1__10_, connection_2__1__9_, 
        connection_2__1__8_, connection_2__1__7_, connection_2__1__6_, 
        connection_2__1__5_, connection_2__1__4_, connection_2__1__3_, 
        connection_2__1__2_, connection_2__1__1_, connection_2__1__0_, 
        connection_2__0__31_, connection_2__0__30_, connection_2__0__29_, 
        connection_2__0__28_, connection_2__0__27_, connection_2__0__26_, 
        connection_2__0__25_, connection_2__0__24_, connection_2__0__23_, 
        connection_2__0__22_, connection_2__0__21_, connection_2__0__20_, 
        connection_2__0__19_, connection_2__0__18_, connection_2__0__17_, 
        connection_2__0__16_, connection_2__0__15_, connection_2__0__14_, 
        connection_2__0__13_, connection_2__0__12_, connection_2__0__11_, 
        connection_2__0__10_, connection_2__0__9_, connection_2__0__8_, 
        connection_2__0__7_, connection_2__0__6_, connection_2__0__5_, 
        connection_2__0__4_, connection_2__0__3_, connection_2__0__2_, 
        connection_2__0__1_, connection_2__0__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[223:222]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_111 first_half_stages_1__group_first_half_0__switch_first_half_1__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_1__6_, 
        connection_valid_1__4_}), .i_data_bus({connection_1__6__31_, 
        connection_1__6__30_, connection_1__6__29_, connection_1__6__28_, 
        connection_1__6__27_, connection_1__6__26_, connection_1__6__25_, 
        connection_1__6__24_, connection_1__6__23_, connection_1__6__22_, 
        connection_1__6__21_, connection_1__6__20_, connection_1__6__19_, 
        connection_1__6__18_, connection_1__6__17_, connection_1__6__16_, 
        connection_1__6__15_, connection_1__6__14_, connection_1__6__13_, 
        connection_1__6__12_, connection_1__6__11_, connection_1__6__10_, 
        connection_1__6__9_, connection_1__6__8_, connection_1__6__7_, 
        connection_1__6__6_, connection_1__6__5_, connection_1__6__4_, 
        connection_1__6__3_, connection_1__6__2_, connection_1__6__1_, 
        connection_1__6__0_, connection_1__4__31_, connection_1__4__30_, 
        connection_1__4__29_, connection_1__4__28_, connection_1__4__27_, 
        connection_1__4__26_, connection_1__4__25_, connection_1__4__24_, 
        connection_1__4__23_, connection_1__4__22_, connection_1__4__21_, 
        connection_1__4__20_, connection_1__4__19_, connection_1__4__18_, 
        connection_1__4__17_, connection_1__4__16_, connection_1__4__15_, 
        connection_1__4__14_, connection_1__4__13_, connection_1__4__12_, 
        connection_1__4__11_, connection_1__4__10_, connection_1__4__9_, 
        connection_1__4__8_, connection_1__4__7_, connection_1__4__6_, 
        connection_1__4__5_, connection_1__4__4_, connection_1__4__3_, 
        connection_1__4__2_, connection_1__4__1_, connection_1__4__0_}), 
        .o_valid({connection_valid_2__3_, connection_valid_2__2_}), 
        .o_data_bus({connection_2__3__31_, connection_2__3__30_, 
        connection_2__3__29_, connection_2__3__28_, connection_2__3__27_, 
        connection_2__3__26_, connection_2__3__25_, connection_2__3__24_, 
        connection_2__3__23_, connection_2__3__22_, connection_2__3__21_, 
        connection_2__3__20_, connection_2__3__19_, connection_2__3__18_, 
        connection_2__3__17_, connection_2__3__16_, connection_2__3__15_, 
        connection_2__3__14_, connection_2__3__13_, connection_2__3__12_, 
        connection_2__3__11_, connection_2__3__10_, connection_2__3__9_, 
        connection_2__3__8_, connection_2__3__7_, connection_2__3__6_, 
        connection_2__3__5_, connection_2__3__4_, connection_2__3__3_, 
        connection_2__3__2_, connection_2__3__1_, connection_2__3__0_, 
        connection_2__2__31_, connection_2__2__30_, connection_2__2__29_, 
        connection_2__2__28_, connection_2__2__27_, connection_2__2__26_, 
        connection_2__2__25_, connection_2__2__24_, connection_2__2__23_, 
        connection_2__2__22_, connection_2__2__21_, connection_2__2__20_, 
        connection_2__2__19_, connection_2__2__18_, connection_2__2__17_, 
        connection_2__2__16_, connection_2__2__15_, connection_2__2__14_, 
        connection_2__2__13_, connection_2__2__12_, connection_2__2__11_, 
        connection_2__2__10_, connection_2__2__9_, connection_2__2__8_, 
        connection_2__2__7_, connection_2__2__6_, connection_2__2__5_, 
        connection_2__2__4_, connection_2__2__3_, connection_2__2__2_, 
        connection_2__2__1_, connection_2__2__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[221:220]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_110 first_half_stages_1__group_first_half_0__switch_first_half_2__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_1__10_, 
        connection_valid_1__8_}), .i_data_bus({connection_1__10__31_, 
        connection_1__10__30_, connection_1__10__29_, connection_1__10__28_, 
        connection_1__10__27_, connection_1__10__26_, connection_1__10__25_, 
        connection_1__10__24_, connection_1__10__23_, connection_1__10__22_, 
        connection_1__10__21_, connection_1__10__20_, connection_1__10__19_, 
        connection_1__10__18_, connection_1__10__17_, connection_1__10__16_, 
        connection_1__10__15_, connection_1__10__14_, connection_1__10__13_, 
        connection_1__10__12_, connection_1__10__11_, connection_1__10__10_, 
        connection_1__10__9_, connection_1__10__8_, connection_1__10__7_, 
        connection_1__10__6_, connection_1__10__5_, connection_1__10__4_, 
        connection_1__10__3_, connection_1__10__2_, connection_1__10__1_, 
        connection_1__10__0_, connection_1__8__31_, connection_1__8__30_, 
        connection_1__8__29_, connection_1__8__28_, connection_1__8__27_, 
        connection_1__8__26_, connection_1__8__25_, connection_1__8__24_, 
        connection_1__8__23_, connection_1__8__22_, connection_1__8__21_, 
        connection_1__8__20_, connection_1__8__19_, connection_1__8__18_, 
        connection_1__8__17_, connection_1__8__16_, connection_1__8__15_, 
        connection_1__8__14_, connection_1__8__13_, connection_1__8__12_, 
        connection_1__8__11_, connection_1__8__10_, connection_1__8__9_, 
        connection_1__8__8_, connection_1__8__7_, connection_1__8__6_, 
        connection_1__8__5_, connection_1__8__4_, connection_1__8__3_, 
        connection_1__8__2_, connection_1__8__1_, connection_1__8__0_}), 
        .o_valid({connection_valid_2__5_, connection_valid_2__4_}), 
        .o_data_bus({connection_2__5__31_, connection_2__5__30_, 
        connection_2__5__29_, connection_2__5__28_, connection_2__5__27_, 
        connection_2__5__26_, connection_2__5__25_, connection_2__5__24_, 
        connection_2__5__23_, connection_2__5__22_, connection_2__5__21_, 
        connection_2__5__20_, connection_2__5__19_, connection_2__5__18_, 
        connection_2__5__17_, connection_2__5__16_, connection_2__5__15_, 
        connection_2__5__14_, connection_2__5__13_, connection_2__5__12_, 
        connection_2__5__11_, connection_2__5__10_, connection_2__5__9_, 
        connection_2__5__8_, connection_2__5__7_, connection_2__5__6_, 
        connection_2__5__5_, connection_2__5__4_, connection_2__5__3_, 
        connection_2__5__2_, connection_2__5__1_, connection_2__5__0_, 
        connection_2__4__31_, connection_2__4__30_, connection_2__4__29_, 
        connection_2__4__28_, connection_2__4__27_, connection_2__4__26_, 
        connection_2__4__25_, connection_2__4__24_, connection_2__4__23_, 
        connection_2__4__22_, connection_2__4__21_, connection_2__4__20_, 
        connection_2__4__19_, connection_2__4__18_, connection_2__4__17_, 
        connection_2__4__16_, connection_2__4__15_, connection_2__4__14_, 
        connection_2__4__13_, connection_2__4__12_, connection_2__4__11_, 
        connection_2__4__10_, connection_2__4__9_, connection_2__4__8_, 
        connection_2__4__7_, connection_2__4__6_, connection_2__4__5_, 
        connection_2__4__4_, connection_2__4__3_, connection_2__4__2_, 
        connection_2__4__1_, connection_2__4__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[219:218]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_109 first_half_stages_1__group_first_half_0__switch_first_half_3__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_1__14_, 
        connection_valid_1__12_}), .i_data_bus({connection_1__14__31_, 
        connection_1__14__30_, connection_1__14__29_, connection_1__14__28_, 
        connection_1__14__27_, connection_1__14__26_, connection_1__14__25_, 
        connection_1__14__24_, connection_1__14__23_, connection_1__14__22_, 
        connection_1__14__21_, connection_1__14__20_, connection_1__14__19_, 
        connection_1__14__18_, connection_1__14__17_, connection_1__14__16_, 
        connection_1__14__15_, connection_1__14__14_, connection_1__14__13_, 
        connection_1__14__12_, connection_1__14__11_, connection_1__14__10_, 
        connection_1__14__9_, connection_1__14__8_, connection_1__14__7_, 
        connection_1__14__6_, connection_1__14__5_, connection_1__14__4_, 
        connection_1__14__3_, connection_1__14__2_, connection_1__14__1_, 
        connection_1__14__0_, connection_1__12__31_, connection_1__12__30_, 
        connection_1__12__29_, connection_1__12__28_, connection_1__12__27_, 
        connection_1__12__26_, connection_1__12__25_, connection_1__12__24_, 
        connection_1__12__23_, connection_1__12__22_, connection_1__12__21_, 
        connection_1__12__20_, connection_1__12__19_, connection_1__12__18_, 
        connection_1__12__17_, connection_1__12__16_, connection_1__12__15_, 
        connection_1__12__14_, connection_1__12__13_, connection_1__12__12_, 
        connection_1__12__11_, connection_1__12__10_, connection_1__12__9_, 
        connection_1__12__8_, connection_1__12__7_, connection_1__12__6_, 
        connection_1__12__5_, connection_1__12__4_, connection_1__12__3_, 
        connection_1__12__2_, connection_1__12__1_, connection_1__12__0_}), 
        .o_valid({connection_valid_2__7_, connection_valid_2__6_}), 
        .o_data_bus({connection_2__7__31_, connection_2__7__30_, 
        connection_2__7__29_, connection_2__7__28_, connection_2__7__27_, 
        connection_2__7__26_, connection_2__7__25_, connection_2__7__24_, 
        connection_2__7__23_, connection_2__7__22_, connection_2__7__21_, 
        connection_2__7__20_, connection_2__7__19_, connection_2__7__18_, 
        connection_2__7__17_, connection_2__7__16_, connection_2__7__15_, 
        connection_2__7__14_, connection_2__7__13_, connection_2__7__12_, 
        connection_2__7__11_, connection_2__7__10_, connection_2__7__9_, 
        connection_2__7__8_, connection_2__7__7_, connection_2__7__6_, 
        connection_2__7__5_, connection_2__7__4_, connection_2__7__3_, 
        connection_2__7__2_, connection_2__7__1_, connection_2__7__0_, 
        connection_2__6__31_, connection_2__6__30_, connection_2__6__29_, 
        connection_2__6__28_, connection_2__6__27_, connection_2__6__26_, 
        connection_2__6__25_, connection_2__6__24_, connection_2__6__23_, 
        connection_2__6__22_, connection_2__6__21_, connection_2__6__20_, 
        connection_2__6__19_, connection_2__6__18_, connection_2__6__17_, 
        connection_2__6__16_, connection_2__6__15_, connection_2__6__14_, 
        connection_2__6__13_, connection_2__6__12_, connection_2__6__11_, 
        connection_2__6__10_, connection_2__6__9_, connection_2__6__8_, 
        connection_2__6__7_, connection_2__6__6_, connection_2__6__5_, 
        connection_2__6__4_, connection_2__6__3_, connection_2__6__2_, 
        connection_2__6__1_, connection_2__6__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[217:216]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_108 first_half_stages_1__group_first_half_0__switch_first_half_4__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_1__3_, 
        connection_valid_1__1_}), .i_data_bus({connection_1__3__31_, 
        connection_1__3__30_, connection_1__3__29_, connection_1__3__28_, 
        connection_1__3__27_, connection_1__3__26_, connection_1__3__25_, 
        connection_1__3__24_, connection_1__3__23_, connection_1__3__22_, 
        connection_1__3__21_, connection_1__3__20_, connection_1__3__19_, 
        connection_1__3__18_, connection_1__3__17_, connection_1__3__16_, 
        connection_1__3__15_, connection_1__3__14_, connection_1__3__13_, 
        connection_1__3__12_, connection_1__3__11_, connection_1__3__10_, 
        connection_1__3__9_, connection_1__3__8_, connection_1__3__7_, 
        connection_1__3__6_, connection_1__3__5_, connection_1__3__4_, 
        connection_1__3__3_, connection_1__3__2_, connection_1__3__1_, 
        connection_1__3__0_, connection_1__1__31_, connection_1__1__30_, 
        connection_1__1__29_, connection_1__1__28_, connection_1__1__27_, 
        connection_1__1__26_, connection_1__1__25_, connection_1__1__24_, 
        connection_1__1__23_, connection_1__1__22_, connection_1__1__21_, 
        connection_1__1__20_, connection_1__1__19_, connection_1__1__18_, 
        connection_1__1__17_, connection_1__1__16_, connection_1__1__15_, 
        connection_1__1__14_, connection_1__1__13_, connection_1__1__12_, 
        connection_1__1__11_, connection_1__1__10_, connection_1__1__9_, 
        connection_1__1__8_, connection_1__1__7_, connection_1__1__6_, 
        connection_1__1__5_, connection_1__1__4_, connection_1__1__3_, 
        connection_1__1__2_, connection_1__1__1_, connection_1__1__0_}), 
        .o_valid({connection_valid_2__9_, connection_valid_2__8_}), 
        .o_data_bus({connection_2__9__31_, connection_2__9__30_, 
        connection_2__9__29_, connection_2__9__28_, connection_2__9__27_, 
        connection_2__9__26_, connection_2__9__25_, connection_2__9__24_, 
        connection_2__9__23_, connection_2__9__22_, connection_2__9__21_, 
        connection_2__9__20_, connection_2__9__19_, connection_2__9__18_, 
        connection_2__9__17_, connection_2__9__16_, connection_2__9__15_, 
        connection_2__9__14_, connection_2__9__13_, connection_2__9__12_, 
        connection_2__9__11_, connection_2__9__10_, connection_2__9__9_, 
        connection_2__9__8_, connection_2__9__7_, connection_2__9__6_, 
        connection_2__9__5_, connection_2__9__4_, connection_2__9__3_, 
        connection_2__9__2_, connection_2__9__1_, connection_2__9__0_, 
        connection_2__8__31_, connection_2__8__30_, connection_2__8__29_, 
        connection_2__8__28_, connection_2__8__27_, connection_2__8__26_, 
        connection_2__8__25_, connection_2__8__24_, connection_2__8__23_, 
        connection_2__8__22_, connection_2__8__21_, connection_2__8__20_, 
        connection_2__8__19_, connection_2__8__18_, connection_2__8__17_, 
        connection_2__8__16_, connection_2__8__15_, connection_2__8__14_, 
        connection_2__8__13_, connection_2__8__12_, connection_2__8__11_, 
        connection_2__8__10_, connection_2__8__9_, connection_2__8__8_, 
        connection_2__8__7_, connection_2__8__6_, connection_2__8__5_, 
        connection_2__8__4_, connection_2__8__3_, connection_2__8__2_, 
        connection_2__8__1_, connection_2__8__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[215:214]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_107 first_half_stages_1__group_first_half_0__switch_first_half_5__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_1__7_, 
        connection_valid_1__5_}), .i_data_bus({connection_1__7__31_, 
        connection_1__7__30_, connection_1__7__29_, connection_1__7__28_, 
        connection_1__7__27_, connection_1__7__26_, connection_1__7__25_, 
        connection_1__7__24_, connection_1__7__23_, connection_1__7__22_, 
        connection_1__7__21_, connection_1__7__20_, connection_1__7__19_, 
        connection_1__7__18_, connection_1__7__17_, connection_1__7__16_, 
        connection_1__7__15_, connection_1__7__14_, connection_1__7__13_, 
        connection_1__7__12_, connection_1__7__11_, connection_1__7__10_, 
        connection_1__7__9_, connection_1__7__8_, connection_1__7__7_, 
        connection_1__7__6_, connection_1__7__5_, connection_1__7__4_, 
        connection_1__7__3_, connection_1__7__2_, connection_1__7__1_, 
        connection_1__7__0_, connection_1__5__31_, connection_1__5__30_, 
        connection_1__5__29_, connection_1__5__28_, connection_1__5__27_, 
        connection_1__5__26_, connection_1__5__25_, connection_1__5__24_, 
        connection_1__5__23_, connection_1__5__22_, connection_1__5__21_, 
        connection_1__5__20_, connection_1__5__19_, connection_1__5__18_, 
        connection_1__5__17_, connection_1__5__16_, connection_1__5__15_, 
        connection_1__5__14_, connection_1__5__13_, connection_1__5__12_, 
        connection_1__5__11_, connection_1__5__10_, connection_1__5__9_, 
        connection_1__5__8_, connection_1__5__7_, connection_1__5__6_, 
        connection_1__5__5_, connection_1__5__4_, connection_1__5__3_, 
        connection_1__5__2_, connection_1__5__1_, connection_1__5__0_}), 
        .o_valid({connection_valid_2__11_, connection_valid_2__10_}), 
        .o_data_bus({connection_2__11__31_, connection_2__11__30_, 
        connection_2__11__29_, connection_2__11__28_, connection_2__11__27_, 
        connection_2__11__26_, connection_2__11__25_, connection_2__11__24_, 
        connection_2__11__23_, connection_2__11__22_, connection_2__11__21_, 
        connection_2__11__20_, connection_2__11__19_, connection_2__11__18_, 
        connection_2__11__17_, connection_2__11__16_, connection_2__11__15_, 
        connection_2__11__14_, connection_2__11__13_, connection_2__11__12_, 
        connection_2__11__11_, connection_2__11__10_, connection_2__11__9_, 
        connection_2__11__8_, connection_2__11__7_, connection_2__11__6_, 
        connection_2__11__5_, connection_2__11__4_, connection_2__11__3_, 
        connection_2__11__2_, connection_2__11__1_, connection_2__11__0_, 
        connection_2__10__31_, connection_2__10__30_, connection_2__10__29_, 
        connection_2__10__28_, connection_2__10__27_, connection_2__10__26_, 
        connection_2__10__25_, connection_2__10__24_, connection_2__10__23_, 
        connection_2__10__22_, connection_2__10__21_, connection_2__10__20_, 
        connection_2__10__19_, connection_2__10__18_, connection_2__10__17_, 
        connection_2__10__16_, connection_2__10__15_, connection_2__10__14_, 
        connection_2__10__13_, connection_2__10__12_, connection_2__10__11_, 
        connection_2__10__10_, connection_2__10__9_, connection_2__10__8_, 
        connection_2__10__7_, connection_2__10__6_, connection_2__10__5_, 
        connection_2__10__4_, connection_2__10__3_, connection_2__10__2_, 
        connection_2__10__1_, connection_2__10__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[213:212]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_106 first_half_stages_1__group_first_half_0__switch_first_half_6__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_1__11_, 
        connection_valid_1__9_}), .i_data_bus({connection_1__11__31_, 
        connection_1__11__30_, connection_1__11__29_, connection_1__11__28_, 
        connection_1__11__27_, connection_1__11__26_, connection_1__11__25_, 
        connection_1__11__24_, connection_1__11__23_, connection_1__11__22_, 
        connection_1__11__21_, connection_1__11__20_, connection_1__11__19_, 
        connection_1__11__18_, connection_1__11__17_, connection_1__11__16_, 
        connection_1__11__15_, connection_1__11__14_, connection_1__11__13_, 
        connection_1__11__12_, connection_1__11__11_, connection_1__11__10_, 
        connection_1__11__9_, connection_1__11__8_, connection_1__11__7_, 
        connection_1__11__6_, connection_1__11__5_, connection_1__11__4_, 
        connection_1__11__3_, connection_1__11__2_, connection_1__11__1_, 
        connection_1__11__0_, connection_1__9__31_, connection_1__9__30_, 
        connection_1__9__29_, connection_1__9__28_, connection_1__9__27_, 
        connection_1__9__26_, connection_1__9__25_, connection_1__9__24_, 
        connection_1__9__23_, connection_1__9__22_, connection_1__9__21_, 
        connection_1__9__20_, connection_1__9__19_, connection_1__9__18_, 
        connection_1__9__17_, connection_1__9__16_, connection_1__9__15_, 
        connection_1__9__14_, connection_1__9__13_, connection_1__9__12_, 
        connection_1__9__11_, connection_1__9__10_, connection_1__9__9_, 
        connection_1__9__8_, connection_1__9__7_, connection_1__9__6_, 
        connection_1__9__5_, connection_1__9__4_, connection_1__9__3_, 
        connection_1__9__2_, connection_1__9__1_, connection_1__9__0_}), 
        .o_valid({connection_valid_2__13_, connection_valid_2__12_}), 
        .o_data_bus({connection_2__13__31_, connection_2__13__30_, 
        connection_2__13__29_, connection_2__13__28_, connection_2__13__27_, 
        connection_2__13__26_, connection_2__13__25_, connection_2__13__24_, 
        connection_2__13__23_, connection_2__13__22_, connection_2__13__21_, 
        connection_2__13__20_, connection_2__13__19_, connection_2__13__18_, 
        connection_2__13__17_, connection_2__13__16_, connection_2__13__15_, 
        connection_2__13__14_, connection_2__13__13_, connection_2__13__12_, 
        connection_2__13__11_, connection_2__13__10_, connection_2__13__9_, 
        connection_2__13__8_, connection_2__13__7_, connection_2__13__6_, 
        connection_2__13__5_, connection_2__13__4_, connection_2__13__3_, 
        connection_2__13__2_, connection_2__13__1_, connection_2__13__0_, 
        connection_2__12__31_, connection_2__12__30_, connection_2__12__29_, 
        connection_2__12__28_, connection_2__12__27_, connection_2__12__26_, 
        connection_2__12__25_, connection_2__12__24_, connection_2__12__23_, 
        connection_2__12__22_, connection_2__12__21_, connection_2__12__20_, 
        connection_2__12__19_, connection_2__12__18_, connection_2__12__17_, 
        connection_2__12__16_, connection_2__12__15_, connection_2__12__14_, 
        connection_2__12__13_, connection_2__12__12_, connection_2__12__11_, 
        connection_2__12__10_, connection_2__12__9_, connection_2__12__8_, 
        connection_2__12__7_, connection_2__12__6_, connection_2__12__5_, 
        connection_2__12__4_, connection_2__12__3_, connection_2__12__2_, 
        connection_2__12__1_, connection_2__12__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[211:210]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_105 first_half_stages_1__group_first_half_0__switch_first_half_7__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_1__15_, 
        connection_valid_1__13_}), .i_data_bus({connection_1__15__31_, 
        connection_1__15__30_, connection_1__15__29_, connection_1__15__28_, 
        connection_1__15__27_, connection_1__15__26_, connection_1__15__25_, 
        connection_1__15__24_, connection_1__15__23_, connection_1__15__22_, 
        connection_1__15__21_, connection_1__15__20_, connection_1__15__19_, 
        connection_1__15__18_, connection_1__15__17_, connection_1__15__16_, 
        connection_1__15__15_, connection_1__15__14_, connection_1__15__13_, 
        connection_1__15__12_, connection_1__15__11_, connection_1__15__10_, 
        connection_1__15__9_, connection_1__15__8_, connection_1__15__7_, 
        connection_1__15__6_, connection_1__15__5_, connection_1__15__4_, 
        connection_1__15__3_, connection_1__15__2_, connection_1__15__1_, 
        connection_1__15__0_, connection_1__13__31_, connection_1__13__30_, 
        connection_1__13__29_, connection_1__13__28_, connection_1__13__27_, 
        connection_1__13__26_, connection_1__13__25_, connection_1__13__24_, 
        connection_1__13__23_, connection_1__13__22_, connection_1__13__21_, 
        connection_1__13__20_, connection_1__13__19_, connection_1__13__18_, 
        connection_1__13__17_, connection_1__13__16_, connection_1__13__15_, 
        connection_1__13__14_, connection_1__13__13_, connection_1__13__12_, 
        connection_1__13__11_, connection_1__13__10_, connection_1__13__9_, 
        connection_1__13__8_, connection_1__13__7_, connection_1__13__6_, 
        connection_1__13__5_, connection_1__13__4_, connection_1__13__3_, 
        connection_1__13__2_, connection_1__13__1_, connection_1__13__0_}), 
        .o_valid({connection_valid_2__15_, connection_valid_2__14_}), 
        .o_data_bus({connection_2__15__31_, connection_2__15__30_, 
        connection_2__15__29_, connection_2__15__28_, connection_2__15__27_, 
        connection_2__15__26_, connection_2__15__25_, connection_2__15__24_, 
        connection_2__15__23_, connection_2__15__22_, connection_2__15__21_, 
        connection_2__15__20_, connection_2__15__19_, connection_2__15__18_, 
        connection_2__15__17_, connection_2__15__16_, connection_2__15__15_, 
        connection_2__15__14_, connection_2__15__13_, connection_2__15__12_, 
        connection_2__15__11_, connection_2__15__10_, connection_2__15__9_, 
        connection_2__15__8_, connection_2__15__7_, connection_2__15__6_, 
        connection_2__15__5_, connection_2__15__4_, connection_2__15__3_, 
        connection_2__15__2_, connection_2__15__1_, connection_2__15__0_, 
        connection_2__14__31_, connection_2__14__30_, connection_2__14__29_, 
        connection_2__14__28_, connection_2__14__27_, connection_2__14__26_, 
        connection_2__14__25_, connection_2__14__24_, connection_2__14__23_, 
        connection_2__14__22_, connection_2__14__21_, connection_2__14__20_, 
        connection_2__14__19_, connection_2__14__18_, connection_2__14__17_, 
        connection_2__14__16_, connection_2__14__15_, connection_2__14__14_, 
        connection_2__14__13_, connection_2__14__12_, connection_2__14__11_, 
        connection_2__14__10_, connection_2__14__9_, connection_2__14__8_, 
        connection_2__14__7_, connection_2__14__6_, connection_2__14__5_, 
        connection_2__14__4_, connection_2__14__3_, connection_2__14__2_, 
        connection_2__14__1_, connection_2__14__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[209:208]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_104 first_half_stages_1__group_first_half_1__switch_first_half_0__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_1__18_, 
        connection_valid_1__16_}), .i_data_bus({connection_1__18__31_, 
        connection_1__18__30_, connection_1__18__29_, connection_1__18__28_, 
        connection_1__18__27_, connection_1__18__26_, connection_1__18__25_, 
        connection_1__18__24_, connection_1__18__23_, connection_1__18__22_, 
        connection_1__18__21_, connection_1__18__20_, connection_1__18__19_, 
        connection_1__18__18_, connection_1__18__17_, connection_1__18__16_, 
        connection_1__18__15_, connection_1__18__14_, connection_1__18__13_, 
        connection_1__18__12_, connection_1__18__11_, connection_1__18__10_, 
        connection_1__18__9_, connection_1__18__8_, connection_1__18__7_, 
        connection_1__18__6_, connection_1__18__5_, connection_1__18__4_, 
        connection_1__18__3_, connection_1__18__2_, connection_1__18__1_, 
        connection_1__18__0_, connection_1__16__31_, connection_1__16__30_, 
        connection_1__16__29_, connection_1__16__28_, connection_1__16__27_, 
        connection_1__16__26_, connection_1__16__25_, connection_1__16__24_, 
        connection_1__16__23_, connection_1__16__22_, connection_1__16__21_, 
        connection_1__16__20_, connection_1__16__19_, connection_1__16__18_, 
        connection_1__16__17_, connection_1__16__16_, connection_1__16__15_, 
        connection_1__16__14_, connection_1__16__13_, connection_1__16__12_, 
        connection_1__16__11_, connection_1__16__10_, connection_1__16__9_, 
        connection_1__16__8_, connection_1__16__7_, connection_1__16__6_, 
        connection_1__16__5_, connection_1__16__4_, connection_1__16__3_, 
        connection_1__16__2_, connection_1__16__1_, connection_1__16__0_}), 
        .o_valid({connection_valid_2__17_, connection_valid_2__16_}), 
        .o_data_bus({connection_2__17__31_, connection_2__17__30_, 
        connection_2__17__29_, connection_2__17__28_, connection_2__17__27_, 
        connection_2__17__26_, connection_2__17__25_, connection_2__17__24_, 
        connection_2__17__23_, connection_2__17__22_, connection_2__17__21_, 
        connection_2__17__20_, connection_2__17__19_, connection_2__17__18_, 
        connection_2__17__17_, connection_2__17__16_, connection_2__17__15_, 
        connection_2__17__14_, connection_2__17__13_, connection_2__17__12_, 
        connection_2__17__11_, connection_2__17__10_, connection_2__17__9_, 
        connection_2__17__8_, connection_2__17__7_, connection_2__17__6_, 
        connection_2__17__5_, connection_2__17__4_, connection_2__17__3_, 
        connection_2__17__2_, connection_2__17__1_, connection_2__17__0_, 
        connection_2__16__31_, connection_2__16__30_, connection_2__16__29_, 
        connection_2__16__28_, connection_2__16__27_, connection_2__16__26_, 
        connection_2__16__25_, connection_2__16__24_, connection_2__16__23_, 
        connection_2__16__22_, connection_2__16__21_, connection_2__16__20_, 
        connection_2__16__19_, connection_2__16__18_, connection_2__16__17_, 
        connection_2__16__16_, connection_2__16__15_, connection_2__16__14_, 
        connection_2__16__13_, connection_2__16__12_, connection_2__16__11_, 
        connection_2__16__10_, connection_2__16__9_, connection_2__16__8_, 
        connection_2__16__7_, connection_2__16__6_, connection_2__16__5_, 
        connection_2__16__4_, connection_2__16__3_, connection_2__16__2_, 
        connection_2__16__1_, connection_2__16__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[207:206]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_103 first_half_stages_1__group_first_half_1__switch_first_half_1__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_1__22_, 
        connection_valid_1__20_}), .i_data_bus({connection_1__22__31_, 
        connection_1__22__30_, connection_1__22__29_, connection_1__22__28_, 
        connection_1__22__27_, connection_1__22__26_, connection_1__22__25_, 
        connection_1__22__24_, connection_1__22__23_, connection_1__22__22_, 
        connection_1__22__21_, connection_1__22__20_, connection_1__22__19_, 
        connection_1__22__18_, connection_1__22__17_, connection_1__22__16_, 
        connection_1__22__15_, connection_1__22__14_, connection_1__22__13_, 
        connection_1__22__12_, connection_1__22__11_, connection_1__22__10_, 
        connection_1__22__9_, connection_1__22__8_, connection_1__22__7_, 
        connection_1__22__6_, connection_1__22__5_, connection_1__22__4_, 
        connection_1__22__3_, connection_1__22__2_, connection_1__22__1_, 
        connection_1__22__0_, connection_1__20__31_, connection_1__20__30_, 
        connection_1__20__29_, connection_1__20__28_, connection_1__20__27_, 
        connection_1__20__26_, connection_1__20__25_, connection_1__20__24_, 
        connection_1__20__23_, connection_1__20__22_, connection_1__20__21_, 
        connection_1__20__20_, connection_1__20__19_, connection_1__20__18_, 
        connection_1__20__17_, connection_1__20__16_, connection_1__20__15_, 
        connection_1__20__14_, connection_1__20__13_, connection_1__20__12_, 
        connection_1__20__11_, connection_1__20__10_, connection_1__20__9_, 
        connection_1__20__8_, connection_1__20__7_, connection_1__20__6_, 
        connection_1__20__5_, connection_1__20__4_, connection_1__20__3_, 
        connection_1__20__2_, connection_1__20__1_, connection_1__20__0_}), 
        .o_valid({connection_valid_2__19_, connection_valid_2__18_}), 
        .o_data_bus({connection_2__19__31_, connection_2__19__30_, 
        connection_2__19__29_, connection_2__19__28_, connection_2__19__27_, 
        connection_2__19__26_, connection_2__19__25_, connection_2__19__24_, 
        connection_2__19__23_, connection_2__19__22_, connection_2__19__21_, 
        connection_2__19__20_, connection_2__19__19_, connection_2__19__18_, 
        connection_2__19__17_, connection_2__19__16_, connection_2__19__15_, 
        connection_2__19__14_, connection_2__19__13_, connection_2__19__12_, 
        connection_2__19__11_, connection_2__19__10_, connection_2__19__9_, 
        connection_2__19__8_, connection_2__19__7_, connection_2__19__6_, 
        connection_2__19__5_, connection_2__19__4_, connection_2__19__3_, 
        connection_2__19__2_, connection_2__19__1_, connection_2__19__0_, 
        connection_2__18__31_, connection_2__18__30_, connection_2__18__29_, 
        connection_2__18__28_, connection_2__18__27_, connection_2__18__26_, 
        connection_2__18__25_, connection_2__18__24_, connection_2__18__23_, 
        connection_2__18__22_, connection_2__18__21_, connection_2__18__20_, 
        connection_2__18__19_, connection_2__18__18_, connection_2__18__17_, 
        connection_2__18__16_, connection_2__18__15_, connection_2__18__14_, 
        connection_2__18__13_, connection_2__18__12_, connection_2__18__11_, 
        connection_2__18__10_, connection_2__18__9_, connection_2__18__8_, 
        connection_2__18__7_, connection_2__18__6_, connection_2__18__5_, 
        connection_2__18__4_, connection_2__18__3_, connection_2__18__2_, 
        connection_2__18__1_, connection_2__18__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[205:204]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_102 first_half_stages_1__group_first_half_1__switch_first_half_2__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_1__26_, 
        connection_valid_1__24_}), .i_data_bus({connection_1__26__31_, 
        connection_1__26__30_, connection_1__26__29_, connection_1__26__28_, 
        connection_1__26__27_, connection_1__26__26_, connection_1__26__25_, 
        connection_1__26__24_, connection_1__26__23_, connection_1__26__22_, 
        connection_1__26__21_, connection_1__26__20_, connection_1__26__19_, 
        connection_1__26__18_, connection_1__26__17_, connection_1__26__16_, 
        connection_1__26__15_, connection_1__26__14_, connection_1__26__13_, 
        connection_1__26__12_, connection_1__26__11_, connection_1__26__10_, 
        connection_1__26__9_, connection_1__26__8_, connection_1__26__7_, 
        connection_1__26__6_, connection_1__26__5_, connection_1__26__4_, 
        connection_1__26__3_, connection_1__26__2_, connection_1__26__1_, 
        connection_1__26__0_, connection_1__24__31_, connection_1__24__30_, 
        connection_1__24__29_, connection_1__24__28_, connection_1__24__27_, 
        connection_1__24__26_, connection_1__24__25_, connection_1__24__24_, 
        connection_1__24__23_, connection_1__24__22_, connection_1__24__21_, 
        connection_1__24__20_, connection_1__24__19_, connection_1__24__18_, 
        connection_1__24__17_, connection_1__24__16_, connection_1__24__15_, 
        connection_1__24__14_, connection_1__24__13_, connection_1__24__12_, 
        connection_1__24__11_, connection_1__24__10_, connection_1__24__9_, 
        connection_1__24__8_, connection_1__24__7_, connection_1__24__6_, 
        connection_1__24__5_, connection_1__24__4_, connection_1__24__3_, 
        connection_1__24__2_, connection_1__24__1_, connection_1__24__0_}), 
        .o_valid({connection_valid_2__21_, connection_valid_2__20_}), 
        .o_data_bus({connection_2__21__31_, connection_2__21__30_, 
        connection_2__21__29_, connection_2__21__28_, connection_2__21__27_, 
        connection_2__21__26_, connection_2__21__25_, connection_2__21__24_, 
        connection_2__21__23_, connection_2__21__22_, connection_2__21__21_, 
        connection_2__21__20_, connection_2__21__19_, connection_2__21__18_, 
        connection_2__21__17_, connection_2__21__16_, connection_2__21__15_, 
        connection_2__21__14_, connection_2__21__13_, connection_2__21__12_, 
        connection_2__21__11_, connection_2__21__10_, connection_2__21__9_, 
        connection_2__21__8_, connection_2__21__7_, connection_2__21__6_, 
        connection_2__21__5_, connection_2__21__4_, connection_2__21__3_, 
        connection_2__21__2_, connection_2__21__1_, connection_2__21__0_, 
        connection_2__20__31_, connection_2__20__30_, connection_2__20__29_, 
        connection_2__20__28_, connection_2__20__27_, connection_2__20__26_, 
        connection_2__20__25_, connection_2__20__24_, connection_2__20__23_, 
        connection_2__20__22_, connection_2__20__21_, connection_2__20__20_, 
        connection_2__20__19_, connection_2__20__18_, connection_2__20__17_, 
        connection_2__20__16_, connection_2__20__15_, connection_2__20__14_, 
        connection_2__20__13_, connection_2__20__12_, connection_2__20__11_, 
        connection_2__20__10_, connection_2__20__9_, connection_2__20__8_, 
        connection_2__20__7_, connection_2__20__6_, connection_2__20__5_, 
        connection_2__20__4_, connection_2__20__3_, connection_2__20__2_, 
        connection_2__20__1_, connection_2__20__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[203:202]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_101 first_half_stages_1__group_first_half_1__switch_first_half_3__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_1__30_, 
        connection_valid_1__28_}), .i_data_bus({connection_1__30__31_, 
        connection_1__30__30_, connection_1__30__29_, connection_1__30__28_, 
        connection_1__30__27_, connection_1__30__26_, connection_1__30__25_, 
        connection_1__30__24_, connection_1__30__23_, connection_1__30__22_, 
        connection_1__30__21_, connection_1__30__20_, connection_1__30__19_, 
        connection_1__30__18_, connection_1__30__17_, connection_1__30__16_, 
        connection_1__30__15_, connection_1__30__14_, connection_1__30__13_, 
        connection_1__30__12_, connection_1__30__11_, connection_1__30__10_, 
        connection_1__30__9_, connection_1__30__8_, connection_1__30__7_, 
        connection_1__30__6_, connection_1__30__5_, connection_1__30__4_, 
        connection_1__30__3_, connection_1__30__2_, connection_1__30__1_, 
        connection_1__30__0_, connection_1__28__31_, connection_1__28__30_, 
        connection_1__28__29_, connection_1__28__28_, connection_1__28__27_, 
        connection_1__28__26_, connection_1__28__25_, connection_1__28__24_, 
        connection_1__28__23_, connection_1__28__22_, connection_1__28__21_, 
        connection_1__28__20_, connection_1__28__19_, connection_1__28__18_, 
        connection_1__28__17_, connection_1__28__16_, connection_1__28__15_, 
        connection_1__28__14_, connection_1__28__13_, connection_1__28__12_, 
        connection_1__28__11_, connection_1__28__10_, connection_1__28__9_, 
        connection_1__28__8_, connection_1__28__7_, connection_1__28__6_, 
        connection_1__28__5_, connection_1__28__4_, connection_1__28__3_, 
        connection_1__28__2_, connection_1__28__1_, connection_1__28__0_}), 
        .o_valid({connection_valid_2__23_, connection_valid_2__22_}), 
        .o_data_bus({connection_2__23__31_, connection_2__23__30_, 
        connection_2__23__29_, connection_2__23__28_, connection_2__23__27_, 
        connection_2__23__26_, connection_2__23__25_, connection_2__23__24_, 
        connection_2__23__23_, connection_2__23__22_, connection_2__23__21_, 
        connection_2__23__20_, connection_2__23__19_, connection_2__23__18_, 
        connection_2__23__17_, connection_2__23__16_, connection_2__23__15_, 
        connection_2__23__14_, connection_2__23__13_, connection_2__23__12_, 
        connection_2__23__11_, connection_2__23__10_, connection_2__23__9_, 
        connection_2__23__8_, connection_2__23__7_, connection_2__23__6_, 
        connection_2__23__5_, connection_2__23__4_, connection_2__23__3_, 
        connection_2__23__2_, connection_2__23__1_, connection_2__23__0_, 
        connection_2__22__31_, connection_2__22__30_, connection_2__22__29_, 
        connection_2__22__28_, connection_2__22__27_, connection_2__22__26_, 
        connection_2__22__25_, connection_2__22__24_, connection_2__22__23_, 
        connection_2__22__22_, connection_2__22__21_, connection_2__22__20_, 
        connection_2__22__19_, connection_2__22__18_, connection_2__22__17_, 
        connection_2__22__16_, connection_2__22__15_, connection_2__22__14_, 
        connection_2__22__13_, connection_2__22__12_, connection_2__22__11_, 
        connection_2__22__10_, connection_2__22__9_, connection_2__22__8_, 
        connection_2__22__7_, connection_2__22__6_, connection_2__22__5_, 
        connection_2__22__4_, connection_2__22__3_, connection_2__22__2_, 
        connection_2__22__1_, connection_2__22__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[201:200]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_100 first_half_stages_1__group_first_half_1__switch_first_half_4__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_1__19_, 
        connection_valid_1__17_}), .i_data_bus({connection_1__19__31_, 
        connection_1__19__30_, connection_1__19__29_, connection_1__19__28_, 
        connection_1__19__27_, connection_1__19__26_, connection_1__19__25_, 
        connection_1__19__24_, connection_1__19__23_, connection_1__19__22_, 
        connection_1__19__21_, connection_1__19__20_, connection_1__19__19_, 
        connection_1__19__18_, connection_1__19__17_, connection_1__19__16_, 
        connection_1__19__15_, connection_1__19__14_, connection_1__19__13_, 
        connection_1__19__12_, connection_1__19__11_, connection_1__19__10_, 
        connection_1__19__9_, connection_1__19__8_, connection_1__19__7_, 
        connection_1__19__6_, connection_1__19__5_, connection_1__19__4_, 
        connection_1__19__3_, connection_1__19__2_, connection_1__19__1_, 
        connection_1__19__0_, connection_1__17__31_, connection_1__17__30_, 
        connection_1__17__29_, connection_1__17__28_, connection_1__17__27_, 
        connection_1__17__26_, connection_1__17__25_, connection_1__17__24_, 
        connection_1__17__23_, connection_1__17__22_, connection_1__17__21_, 
        connection_1__17__20_, connection_1__17__19_, connection_1__17__18_, 
        connection_1__17__17_, connection_1__17__16_, connection_1__17__15_, 
        connection_1__17__14_, connection_1__17__13_, connection_1__17__12_, 
        connection_1__17__11_, connection_1__17__10_, connection_1__17__9_, 
        connection_1__17__8_, connection_1__17__7_, connection_1__17__6_, 
        connection_1__17__5_, connection_1__17__4_, connection_1__17__3_, 
        connection_1__17__2_, connection_1__17__1_, connection_1__17__0_}), 
        .o_valid({connection_valid_2__25_, connection_valid_2__24_}), 
        .o_data_bus({connection_2__25__31_, connection_2__25__30_, 
        connection_2__25__29_, connection_2__25__28_, connection_2__25__27_, 
        connection_2__25__26_, connection_2__25__25_, connection_2__25__24_, 
        connection_2__25__23_, connection_2__25__22_, connection_2__25__21_, 
        connection_2__25__20_, connection_2__25__19_, connection_2__25__18_, 
        connection_2__25__17_, connection_2__25__16_, connection_2__25__15_, 
        connection_2__25__14_, connection_2__25__13_, connection_2__25__12_, 
        connection_2__25__11_, connection_2__25__10_, connection_2__25__9_, 
        connection_2__25__8_, connection_2__25__7_, connection_2__25__6_, 
        connection_2__25__5_, connection_2__25__4_, connection_2__25__3_, 
        connection_2__25__2_, connection_2__25__1_, connection_2__25__0_, 
        connection_2__24__31_, connection_2__24__30_, connection_2__24__29_, 
        connection_2__24__28_, connection_2__24__27_, connection_2__24__26_, 
        connection_2__24__25_, connection_2__24__24_, connection_2__24__23_, 
        connection_2__24__22_, connection_2__24__21_, connection_2__24__20_, 
        connection_2__24__19_, connection_2__24__18_, connection_2__24__17_, 
        connection_2__24__16_, connection_2__24__15_, connection_2__24__14_, 
        connection_2__24__13_, connection_2__24__12_, connection_2__24__11_, 
        connection_2__24__10_, connection_2__24__9_, connection_2__24__8_, 
        connection_2__24__7_, connection_2__24__6_, connection_2__24__5_, 
        connection_2__24__4_, connection_2__24__3_, connection_2__24__2_, 
        connection_2__24__1_, connection_2__24__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[199:198]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_99 first_half_stages_1__group_first_half_1__switch_first_half_5__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_1__23_, 
        connection_valid_1__21_}), .i_data_bus({connection_1__23__31_, 
        connection_1__23__30_, connection_1__23__29_, connection_1__23__28_, 
        connection_1__23__27_, connection_1__23__26_, connection_1__23__25_, 
        connection_1__23__24_, connection_1__23__23_, connection_1__23__22_, 
        connection_1__23__21_, connection_1__23__20_, connection_1__23__19_, 
        connection_1__23__18_, connection_1__23__17_, connection_1__23__16_, 
        connection_1__23__15_, connection_1__23__14_, connection_1__23__13_, 
        connection_1__23__12_, connection_1__23__11_, connection_1__23__10_, 
        connection_1__23__9_, connection_1__23__8_, connection_1__23__7_, 
        connection_1__23__6_, connection_1__23__5_, connection_1__23__4_, 
        connection_1__23__3_, connection_1__23__2_, connection_1__23__1_, 
        connection_1__23__0_, connection_1__21__31_, connection_1__21__30_, 
        connection_1__21__29_, connection_1__21__28_, connection_1__21__27_, 
        connection_1__21__26_, connection_1__21__25_, connection_1__21__24_, 
        connection_1__21__23_, connection_1__21__22_, connection_1__21__21_, 
        connection_1__21__20_, connection_1__21__19_, connection_1__21__18_, 
        connection_1__21__17_, connection_1__21__16_, connection_1__21__15_, 
        connection_1__21__14_, connection_1__21__13_, connection_1__21__12_, 
        connection_1__21__11_, connection_1__21__10_, connection_1__21__9_, 
        connection_1__21__8_, connection_1__21__7_, connection_1__21__6_, 
        connection_1__21__5_, connection_1__21__4_, connection_1__21__3_, 
        connection_1__21__2_, connection_1__21__1_, connection_1__21__0_}), 
        .o_valid({connection_valid_2__27_, connection_valid_2__26_}), 
        .o_data_bus({connection_2__27__31_, connection_2__27__30_, 
        connection_2__27__29_, connection_2__27__28_, connection_2__27__27_, 
        connection_2__27__26_, connection_2__27__25_, connection_2__27__24_, 
        connection_2__27__23_, connection_2__27__22_, connection_2__27__21_, 
        connection_2__27__20_, connection_2__27__19_, connection_2__27__18_, 
        connection_2__27__17_, connection_2__27__16_, connection_2__27__15_, 
        connection_2__27__14_, connection_2__27__13_, connection_2__27__12_, 
        connection_2__27__11_, connection_2__27__10_, connection_2__27__9_, 
        connection_2__27__8_, connection_2__27__7_, connection_2__27__6_, 
        connection_2__27__5_, connection_2__27__4_, connection_2__27__3_, 
        connection_2__27__2_, connection_2__27__1_, connection_2__27__0_, 
        connection_2__26__31_, connection_2__26__30_, connection_2__26__29_, 
        connection_2__26__28_, connection_2__26__27_, connection_2__26__26_, 
        connection_2__26__25_, connection_2__26__24_, connection_2__26__23_, 
        connection_2__26__22_, connection_2__26__21_, connection_2__26__20_, 
        connection_2__26__19_, connection_2__26__18_, connection_2__26__17_, 
        connection_2__26__16_, connection_2__26__15_, connection_2__26__14_, 
        connection_2__26__13_, connection_2__26__12_, connection_2__26__11_, 
        connection_2__26__10_, connection_2__26__9_, connection_2__26__8_, 
        connection_2__26__7_, connection_2__26__6_, connection_2__26__5_, 
        connection_2__26__4_, connection_2__26__3_, connection_2__26__2_, 
        connection_2__26__1_, connection_2__26__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[197:196]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_98 first_half_stages_1__group_first_half_1__switch_first_half_6__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_1__27_, 
        connection_valid_1__25_}), .i_data_bus({connection_1__27__31_, 
        connection_1__27__30_, connection_1__27__29_, connection_1__27__28_, 
        connection_1__27__27_, connection_1__27__26_, connection_1__27__25_, 
        connection_1__27__24_, connection_1__27__23_, connection_1__27__22_, 
        connection_1__27__21_, connection_1__27__20_, connection_1__27__19_, 
        connection_1__27__18_, connection_1__27__17_, connection_1__27__16_, 
        connection_1__27__15_, connection_1__27__14_, connection_1__27__13_, 
        connection_1__27__12_, connection_1__27__11_, connection_1__27__10_, 
        connection_1__27__9_, connection_1__27__8_, connection_1__27__7_, 
        connection_1__27__6_, connection_1__27__5_, connection_1__27__4_, 
        connection_1__27__3_, connection_1__27__2_, connection_1__27__1_, 
        connection_1__27__0_, connection_1__25__31_, connection_1__25__30_, 
        connection_1__25__29_, connection_1__25__28_, connection_1__25__27_, 
        connection_1__25__26_, connection_1__25__25_, connection_1__25__24_, 
        connection_1__25__23_, connection_1__25__22_, connection_1__25__21_, 
        connection_1__25__20_, connection_1__25__19_, connection_1__25__18_, 
        connection_1__25__17_, connection_1__25__16_, connection_1__25__15_, 
        connection_1__25__14_, connection_1__25__13_, connection_1__25__12_, 
        connection_1__25__11_, connection_1__25__10_, connection_1__25__9_, 
        connection_1__25__8_, connection_1__25__7_, connection_1__25__6_, 
        connection_1__25__5_, connection_1__25__4_, connection_1__25__3_, 
        connection_1__25__2_, connection_1__25__1_, connection_1__25__0_}), 
        .o_valid({connection_valid_2__29_, connection_valid_2__28_}), 
        .o_data_bus({connection_2__29__31_, connection_2__29__30_, 
        connection_2__29__29_, connection_2__29__28_, connection_2__29__27_, 
        connection_2__29__26_, connection_2__29__25_, connection_2__29__24_, 
        connection_2__29__23_, connection_2__29__22_, connection_2__29__21_, 
        connection_2__29__20_, connection_2__29__19_, connection_2__29__18_, 
        connection_2__29__17_, connection_2__29__16_, connection_2__29__15_, 
        connection_2__29__14_, connection_2__29__13_, connection_2__29__12_, 
        connection_2__29__11_, connection_2__29__10_, connection_2__29__9_, 
        connection_2__29__8_, connection_2__29__7_, connection_2__29__6_, 
        connection_2__29__5_, connection_2__29__4_, connection_2__29__3_, 
        connection_2__29__2_, connection_2__29__1_, connection_2__29__0_, 
        connection_2__28__31_, connection_2__28__30_, connection_2__28__29_, 
        connection_2__28__28_, connection_2__28__27_, connection_2__28__26_, 
        connection_2__28__25_, connection_2__28__24_, connection_2__28__23_, 
        connection_2__28__22_, connection_2__28__21_, connection_2__28__20_, 
        connection_2__28__19_, connection_2__28__18_, connection_2__28__17_, 
        connection_2__28__16_, connection_2__28__15_, connection_2__28__14_, 
        connection_2__28__13_, connection_2__28__12_, connection_2__28__11_, 
        connection_2__28__10_, connection_2__28__9_, connection_2__28__8_, 
        connection_2__28__7_, connection_2__28__6_, connection_2__28__5_, 
        connection_2__28__4_, connection_2__28__3_, connection_2__28__2_, 
        connection_2__28__1_, connection_2__28__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[195:194]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_97 first_half_stages_1__group_first_half_1__switch_first_half_7__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_1__31_, 
        connection_valid_1__29_}), .i_data_bus({connection_1__31__31_, 
        connection_1__31__30_, connection_1__31__29_, connection_1__31__28_, 
        connection_1__31__27_, connection_1__31__26_, connection_1__31__25_, 
        connection_1__31__24_, connection_1__31__23_, connection_1__31__22_, 
        connection_1__31__21_, connection_1__31__20_, connection_1__31__19_, 
        connection_1__31__18_, connection_1__31__17_, connection_1__31__16_, 
        connection_1__31__15_, connection_1__31__14_, connection_1__31__13_, 
        connection_1__31__12_, connection_1__31__11_, connection_1__31__10_, 
        connection_1__31__9_, connection_1__31__8_, connection_1__31__7_, 
        connection_1__31__6_, connection_1__31__5_, connection_1__31__4_, 
        connection_1__31__3_, connection_1__31__2_, connection_1__31__1_, 
        connection_1__31__0_, connection_1__29__31_, connection_1__29__30_, 
        connection_1__29__29_, connection_1__29__28_, connection_1__29__27_, 
        connection_1__29__26_, connection_1__29__25_, connection_1__29__24_, 
        connection_1__29__23_, connection_1__29__22_, connection_1__29__21_, 
        connection_1__29__20_, connection_1__29__19_, connection_1__29__18_, 
        connection_1__29__17_, connection_1__29__16_, connection_1__29__15_, 
        connection_1__29__14_, connection_1__29__13_, connection_1__29__12_, 
        connection_1__29__11_, connection_1__29__10_, connection_1__29__9_, 
        connection_1__29__8_, connection_1__29__7_, connection_1__29__6_, 
        connection_1__29__5_, connection_1__29__4_, connection_1__29__3_, 
        connection_1__29__2_, connection_1__29__1_, connection_1__29__0_}), 
        .o_valid({connection_valid_2__31_, connection_valid_2__30_}), 
        .o_data_bus({connection_2__31__31_, connection_2__31__30_, 
        connection_2__31__29_, connection_2__31__28_, connection_2__31__27_, 
        connection_2__31__26_, connection_2__31__25_, connection_2__31__24_, 
        connection_2__31__23_, connection_2__31__22_, connection_2__31__21_, 
        connection_2__31__20_, connection_2__31__19_, connection_2__31__18_, 
        connection_2__31__17_, connection_2__31__16_, connection_2__31__15_, 
        connection_2__31__14_, connection_2__31__13_, connection_2__31__12_, 
        connection_2__31__11_, connection_2__31__10_, connection_2__31__9_, 
        connection_2__31__8_, connection_2__31__7_, connection_2__31__6_, 
        connection_2__31__5_, connection_2__31__4_, connection_2__31__3_, 
        connection_2__31__2_, connection_2__31__1_, connection_2__31__0_, 
        connection_2__30__31_, connection_2__30__30_, connection_2__30__29_, 
        connection_2__30__28_, connection_2__30__27_, connection_2__30__26_, 
        connection_2__30__25_, connection_2__30__24_, connection_2__30__23_, 
        connection_2__30__22_, connection_2__30__21_, connection_2__30__20_, 
        connection_2__30__19_, connection_2__30__18_, connection_2__30__17_, 
        connection_2__30__16_, connection_2__30__15_, connection_2__30__14_, 
        connection_2__30__13_, connection_2__30__12_, connection_2__30__11_, 
        connection_2__30__10_, connection_2__30__9_, connection_2__30__8_, 
        connection_2__30__7_, connection_2__30__6_, connection_2__30__5_, 
        connection_2__30__4_, connection_2__30__3_, connection_2__30__2_, 
        connection_2__30__1_, connection_2__30__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[193:192]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_96 first_half_stages_2__group_first_half_0__switch_first_half_0__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__2_, 
        connection_valid_2__0_}), .i_data_bus({connection_2__2__31_, 
        connection_2__2__30_, connection_2__2__29_, connection_2__2__28_, 
        connection_2__2__27_, connection_2__2__26_, connection_2__2__25_, 
        connection_2__2__24_, connection_2__2__23_, connection_2__2__22_, 
        connection_2__2__21_, connection_2__2__20_, connection_2__2__19_, 
        connection_2__2__18_, connection_2__2__17_, connection_2__2__16_, 
        connection_2__2__15_, connection_2__2__14_, connection_2__2__13_, 
        connection_2__2__12_, connection_2__2__11_, connection_2__2__10_, 
        connection_2__2__9_, connection_2__2__8_, connection_2__2__7_, 
        connection_2__2__6_, connection_2__2__5_, connection_2__2__4_, 
        connection_2__2__3_, connection_2__2__2_, connection_2__2__1_, 
        connection_2__2__0_, connection_2__0__31_, connection_2__0__30_, 
        connection_2__0__29_, connection_2__0__28_, connection_2__0__27_, 
        connection_2__0__26_, connection_2__0__25_, connection_2__0__24_, 
        connection_2__0__23_, connection_2__0__22_, connection_2__0__21_, 
        connection_2__0__20_, connection_2__0__19_, connection_2__0__18_, 
        connection_2__0__17_, connection_2__0__16_, connection_2__0__15_, 
        connection_2__0__14_, connection_2__0__13_, connection_2__0__12_, 
        connection_2__0__11_, connection_2__0__10_, connection_2__0__9_, 
        connection_2__0__8_, connection_2__0__7_, connection_2__0__6_, 
        connection_2__0__5_, connection_2__0__4_, connection_2__0__3_, 
        connection_2__0__2_, connection_2__0__1_, connection_2__0__0_}), 
        .o_valid({connection_valid_3__1_, connection_valid_3__0_}), 
        .o_data_bus({connection_3__1__31_, connection_3__1__30_, 
        connection_3__1__29_, connection_3__1__28_, connection_3__1__27_, 
        connection_3__1__26_, connection_3__1__25_, connection_3__1__24_, 
        connection_3__1__23_, connection_3__1__22_, connection_3__1__21_, 
        connection_3__1__20_, connection_3__1__19_, connection_3__1__18_, 
        connection_3__1__17_, connection_3__1__16_, connection_3__1__15_, 
        connection_3__1__14_, connection_3__1__13_, connection_3__1__12_, 
        connection_3__1__11_, connection_3__1__10_, connection_3__1__9_, 
        connection_3__1__8_, connection_3__1__7_, connection_3__1__6_, 
        connection_3__1__5_, connection_3__1__4_, connection_3__1__3_, 
        connection_3__1__2_, connection_3__1__1_, connection_3__1__0_, 
        connection_3__0__31_, connection_3__0__30_, connection_3__0__29_, 
        connection_3__0__28_, connection_3__0__27_, connection_3__0__26_, 
        connection_3__0__25_, connection_3__0__24_, connection_3__0__23_, 
        connection_3__0__22_, connection_3__0__21_, connection_3__0__20_, 
        connection_3__0__19_, connection_3__0__18_, connection_3__0__17_, 
        connection_3__0__16_, connection_3__0__15_, connection_3__0__14_, 
        connection_3__0__13_, connection_3__0__12_, connection_3__0__11_, 
        connection_3__0__10_, connection_3__0__9_, connection_3__0__8_, 
        connection_3__0__7_, connection_3__0__6_, connection_3__0__5_, 
        connection_3__0__4_, connection_3__0__3_, connection_3__0__2_, 
        connection_3__0__1_, connection_3__0__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[191:190]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_95 first_half_stages_2__group_first_half_0__switch_first_half_1__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__6_, 
        connection_valid_2__4_}), .i_data_bus({connection_2__6__31_, 
        connection_2__6__30_, connection_2__6__29_, connection_2__6__28_, 
        connection_2__6__27_, connection_2__6__26_, connection_2__6__25_, 
        connection_2__6__24_, connection_2__6__23_, connection_2__6__22_, 
        connection_2__6__21_, connection_2__6__20_, connection_2__6__19_, 
        connection_2__6__18_, connection_2__6__17_, connection_2__6__16_, 
        connection_2__6__15_, connection_2__6__14_, connection_2__6__13_, 
        connection_2__6__12_, connection_2__6__11_, connection_2__6__10_, 
        connection_2__6__9_, connection_2__6__8_, connection_2__6__7_, 
        connection_2__6__6_, connection_2__6__5_, connection_2__6__4_, 
        connection_2__6__3_, connection_2__6__2_, connection_2__6__1_, 
        connection_2__6__0_, connection_2__4__31_, connection_2__4__30_, 
        connection_2__4__29_, connection_2__4__28_, connection_2__4__27_, 
        connection_2__4__26_, connection_2__4__25_, connection_2__4__24_, 
        connection_2__4__23_, connection_2__4__22_, connection_2__4__21_, 
        connection_2__4__20_, connection_2__4__19_, connection_2__4__18_, 
        connection_2__4__17_, connection_2__4__16_, connection_2__4__15_, 
        connection_2__4__14_, connection_2__4__13_, connection_2__4__12_, 
        connection_2__4__11_, connection_2__4__10_, connection_2__4__9_, 
        connection_2__4__8_, connection_2__4__7_, connection_2__4__6_, 
        connection_2__4__5_, connection_2__4__4_, connection_2__4__3_, 
        connection_2__4__2_, connection_2__4__1_, connection_2__4__0_}), 
        .o_valid({connection_valid_3__3_, connection_valid_3__2_}), 
        .o_data_bus({connection_3__3__31_, connection_3__3__30_, 
        connection_3__3__29_, connection_3__3__28_, connection_3__3__27_, 
        connection_3__3__26_, connection_3__3__25_, connection_3__3__24_, 
        connection_3__3__23_, connection_3__3__22_, connection_3__3__21_, 
        connection_3__3__20_, connection_3__3__19_, connection_3__3__18_, 
        connection_3__3__17_, connection_3__3__16_, connection_3__3__15_, 
        connection_3__3__14_, connection_3__3__13_, connection_3__3__12_, 
        connection_3__3__11_, connection_3__3__10_, connection_3__3__9_, 
        connection_3__3__8_, connection_3__3__7_, connection_3__3__6_, 
        connection_3__3__5_, connection_3__3__4_, connection_3__3__3_, 
        connection_3__3__2_, connection_3__3__1_, connection_3__3__0_, 
        connection_3__2__31_, connection_3__2__30_, connection_3__2__29_, 
        connection_3__2__28_, connection_3__2__27_, connection_3__2__26_, 
        connection_3__2__25_, connection_3__2__24_, connection_3__2__23_, 
        connection_3__2__22_, connection_3__2__21_, connection_3__2__20_, 
        connection_3__2__19_, connection_3__2__18_, connection_3__2__17_, 
        connection_3__2__16_, connection_3__2__15_, connection_3__2__14_, 
        connection_3__2__13_, connection_3__2__12_, connection_3__2__11_, 
        connection_3__2__10_, connection_3__2__9_, connection_3__2__8_, 
        connection_3__2__7_, connection_3__2__6_, connection_3__2__5_, 
        connection_3__2__4_, connection_3__2__3_, connection_3__2__2_, 
        connection_3__2__1_, connection_3__2__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[189:188]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_94 first_half_stages_2__group_first_half_0__switch_first_half_2__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__3_, 
        connection_valid_2__1_}), .i_data_bus({connection_2__3__31_, 
        connection_2__3__30_, connection_2__3__29_, connection_2__3__28_, 
        connection_2__3__27_, connection_2__3__26_, connection_2__3__25_, 
        connection_2__3__24_, connection_2__3__23_, connection_2__3__22_, 
        connection_2__3__21_, connection_2__3__20_, connection_2__3__19_, 
        connection_2__3__18_, connection_2__3__17_, connection_2__3__16_, 
        connection_2__3__15_, connection_2__3__14_, connection_2__3__13_, 
        connection_2__3__12_, connection_2__3__11_, connection_2__3__10_, 
        connection_2__3__9_, connection_2__3__8_, connection_2__3__7_, 
        connection_2__3__6_, connection_2__3__5_, connection_2__3__4_, 
        connection_2__3__3_, connection_2__3__2_, connection_2__3__1_, 
        connection_2__3__0_, connection_2__1__31_, connection_2__1__30_, 
        connection_2__1__29_, connection_2__1__28_, connection_2__1__27_, 
        connection_2__1__26_, connection_2__1__25_, connection_2__1__24_, 
        connection_2__1__23_, connection_2__1__22_, connection_2__1__21_, 
        connection_2__1__20_, connection_2__1__19_, connection_2__1__18_, 
        connection_2__1__17_, connection_2__1__16_, connection_2__1__15_, 
        connection_2__1__14_, connection_2__1__13_, connection_2__1__12_, 
        connection_2__1__11_, connection_2__1__10_, connection_2__1__9_, 
        connection_2__1__8_, connection_2__1__7_, connection_2__1__6_, 
        connection_2__1__5_, connection_2__1__4_, connection_2__1__3_, 
        connection_2__1__2_, connection_2__1__1_, connection_2__1__0_}), 
        .o_valid({connection_valid_3__5_, connection_valid_3__4_}), 
        .o_data_bus({connection_3__5__31_, connection_3__5__30_, 
        connection_3__5__29_, connection_3__5__28_, connection_3__5__27_, 
        connection_3__5__26_, connection_3__5__25_, connection_3__5__24_, 
        connection_3__5__23_, connection_3__5__22_, connection_3__5__21_, 
        connection_3__5__20_, connection_3__5__19_, connection_3__5__18_, 
        connection_3__5__17_, connection_3__5__16_, connection_3__5__15_, 
        connection_3__5__14_, connection_3__5__13_, connection_3__5__12_, 
        connection_3__5__11_, connection_3__5__10_, connection_3__5__9_, 
        connection_3__5__8_, connection_3__5__7_, connection_3__5__6_, 
        connection_3__5__5_, connection_3__5__4_, connection_3__5__3_, 
        connection_3__5__2_, connection_3__5__1_, connection_3__5__0_, 
        connection_3__4__31_, connection_3__4__30_, connection_3__4__29_, 
        connection_3__4__28_, connection_3__4__27_, connection_3__4__26_, 
        connection_3__4__25_, connection_3__4__24_, connection_3__4__23_, 
        connection_3__4__22_, connection_3__4__21_, connection_3__4__20_, 
        connection_3__4__19_, connection_3__4__18_, connection_3__4__17_, 
        connection_3__4__16_, connection_3__4__15_, connection_3__4__14_, 
        connection_3__4__13_, connection_3__4__12_, connection_3__4__11_, 
        connection_3__4__10_, connection_3__4__9_, connection_3__4__8_, 
        connection_3__4__7_, connection_3__4__6_, connection_3__4__5_, 
        connection_3__4__4_, connection_3__4__3_, connection_3__4__2_, 
        connection_3__4__1_, connection_3__4__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[187:186]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_93 first_half_stages_2__group_first_half_0__switch_first_half_3__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__7_, 
        connection_valid_2__5_}), .i_data_bus({connection_2__7__31_, 
        connection_2__7__30_, connection_2__7__29_, connection_2__7__28_, 
        connection_2__7__27_, connection_2__7__26_, connection_2__7__25_, 
        connection_2__7__24_, connection_2__7__23_, connection_2__7__22_, 
        connection_2__7__21_, connection_2__7__20_, connection_2__7__19_, 
        connection_2__7__18_, connection_2__7__17_, connection_2__7__16_, 
        connection_2__7__15_, connection_2__7__14_, connection_2__7__13_, 
        connection_2__7__12_, connection_2__7__11_, connection_2__7__10_, 
        connection_2__7__9_, connection_2__7__8_, connection_2__7__7_, 
        connection_2__7__6_, connection_2__7__5_, connection_2__7__4_, 
        connection_2__7__3_, connection_2__7__2_, connection_2__7__1_, 
        connection_2__7__0_, connection_2__5__31_, connection_2__5__30_, 
        connection_2__5__29_, connection_2__5__28_, connection_2__5__27_, 
        connection_2__5__26_, connection_2__5__25_, connection_2__5__24_, 
        connection_2__5__23_, connection_2__5__22_, connection_2__5__21_, 
        connection_2__5__20_, connection_2__5__19_, connection_2__5__18_, 
        connection_2__5__17_, connection_2__5__16_, connection_2__5__15_, 
        connection_2__5__14_, connection_2__5__13_, connection_2__5__12_, 
        connection_2__5__11_, connection_2__5__10_, connection_2__5__9_, 
        connection_2__5__8_, connection_2__5__7_, connection_2__5__6_, 
        connection_2__5__5_, connection_2__5__4_, connection_2__5__3_, 
        connection_2__5__2_, connection_2__5__1_, connection_2__5__0_}), 
        .o_valid({connection_valid_3__7_, connection_valid_3__6_}), 
        .o_data_bus({connection_3__7__31_, connection_3__7__30_, 
        connection_3__7__29_, connection_3__7__28_, connection_3__7__27_, 
        connection_3__7__26_, connection_3__7__25_, connection_3__7__24_, 
        connection_3__7__23_, connection_3__7__22_, connection_3__7__21_, 
        connection_3__7__20_, connection_3__7__19_, connection_3__7__18_, 
        connection_3__7__17_, connection_3__7__16_, connection_3__7__15_, 
        connection_3__7__14_, connection_3__7__13_, connection_3__7__12_, 
        connection_3__7__11_, connection_3__7__10_, connection_3__7__9_, 
        connection_3__7__8_, connection_3__7__7_, connection_3__7__6_, 
        connection_3__7__5_, connection_3__7__4_, connection_3__7__3_, 
        connection_3__7__2_, connection_3__7__1_, connection_3__7__0_, 
        connection_3__6__31_, connection_3__6__30_, connection_3__6__29_, 
        connection_3__6__28_, connection_3__6__27_, connection_3__6__26_, 
        connection_3__6__25_, connection_3__6__24_, connection_3__6__23_, 
        connection_3__6__22_, connection_3__6__21_, connection_3__6__20_, 
        connection_3__6__19_, connection_3__6__18_, connection_3__6__17_, 
        connection_3__6__16_, connection_3__6__15_, connection_3__6__14_, 
        connection_3__6__13_, connection_3__6__12_, connection_3__6__11_, 
        connection_3__6__10_, connection_3__6__9_, connection_3__6__8_, 
        connection_3__6__7_, connection_3__6__6_, connection_3__6__5_, 
        connection_3__6__4_, connection_3__6__3_, connection_3__6__2_, 
        connection_3__6__1_, connection_3__6__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[185:184]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_92 first_half_stages_2__group_first_half_1__switch_first_half_0__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__10_, 
        connection_valid_2__8_}), .i_data_bus({connection_2__10__31_, 
        connection_2__10__30_, connection_2__10__29_, connection_2__10__28_, 
        connection_2__10__27_, connection_2__10__26_, connection_2__10__25_, 
        connection_2__10__24_, connection_2__10__23_, connection_2__10__22_, 
        connection_2__10__21_, connection_2__10__20_, connection_2__10__19_, 
        connection_2__10__18_, connection_2__10__17_, connection_2__10__16_, 
        connection_2__10__15_, connection_2__10__14_, connection_2__10__13_, 
        connection_2__10__12_, connection_2__10__11_, connection_2__10__10_, 
        connection_2__10__9_, connection_2__10__8_, connection_2__10__7_, 
        connection_2__10__6_, connection_2__10__5_, connection_2__10__4_, 
        connection_2__10__3_, connection_2__10__2_, connection_2__10__1_, 
        connection_2__10__0_, connection_2__8__31_, connection_2__8__30_, 
        connection_2__8__29_, connection_2__8__28_, connection_2__8__27_, 
        connection_2__8__26_, connection_2__8__25_, connection_2__8__24_, 
        connection_2__8__23_, connection_2__8__22_, connection_2__8__21_, 
        connection_2__8__20_, connection_2__8__19_, connection_2__8__18_, 
        connection_2__8__17_, connection_2__8__16_, connection_2__8__15_, 
        connection_2__8__14_, connection_2__8__13_, connection_2__8__12_, 
        connection_2__8__11_, connection_2__8__10_, connection_2__8__9_, 
        connection_2__8__8_, connection_2__8__7_, connection_2__8__6_, 
        connection_2__8__5_, connection_2__8__4_, connection_2__8__3_, 
        connection_2__8__2_, connection_2__8__1_, connection_2__8__0_}), 
        .o_valid({connection_valid_3__9_, connection_valid_3__8_}), 
        .o_data_bus({connection_3__9__31_, connection_3__9__30_, 
        connection_3__9__29_, connection_3__9__28_, connection_3__9__27_, 
        connection_3__9__26_, connection_3__9__25_, connection_3__9__24_, 
        connection_3__9__23_, connection_3__9__22_, connection_3__9__21_, 
        connection_3__9__20_, connection_3__9__19_, connection_3__9__18_, 
        connection_3__9__17_, connection_3__9__16_, connection_3__9__15_, 
        connection_3__9__14_, connection_3__9__13_, connection_3__9__12_, 
        connection_3__9__11_, connection_3__9__10_, connection_3__9__9_, 
        connection_3__9__8_, connection_3__9__7_, connection_3__9__6_, 
        connection_3__9__5_, connection_3__9__4_, connection_3__9__3_, 
        connection_3__9__2_, connection_3__9__1_, connection_3__9__0_, 
        connection_3__8__31_, connection_3__8__30_, connection_3__8__29_, 
        connection_3__8__28_, connection_3__8__27_, connection_3__8__26_, 
        connection_3__8__25_, connection_3__8__24_, connection_3__8__23_, 
        connection_3__8__22_, connection_3__8__21_, connection_3__8__20_, 
        connection_3__8__19_, connection_3__8__18_, connection_3__8__17_, 
        connection_3__8__16_, connection_3__8__15_, connection_3__8__14_, 
        connection_3__8__13_, connection_3__8__12_, connection_3__8__11_, 
        connection_3__8__10_, connection_3__8__9_, connection_3__8__8_, 
        connection_3__8__7_, connection_3__8__6_, connection_3__8__5_, 
        connection_3__8__4_, connection_3__8__3_, connection_3__8__2_, 
        connection_3__8__1_, connection_3__8__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[183:182]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_91 first_half_stages_2__group_first_half_1__switch_first_half_1__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__14_, 
        connection_valid_2__12_}), .i_data_bus({connection_2__14__31_, 
        connection_2__14__30_, connection_2__14__29_, connection_2__14__28_, 
        connection_2__14__27_, connection_2__14__26_, connection_2__14__25_, 
        connection_2__14__24_, connection_2__14__23_, connection_2__14__22_, 
        connection_2__14__21_, connection_2__14__20_, connection_2__14__19_, 
        connection_2__14__18_, connection_2__14__17_, connection_2__14__16_, 
        connection_2__14__15_, connection_2__14__14_, connection_2__14__13_, 
        connection_2__14__12_, connection_2__14__11_, connection_2__14__10_, 
        connection_2__14__9_, connection_2__14__8_, connection_2__14__7_, 
        connection_2__14__6_, connection_2__14__5_, connection_2__14__4_, 
        connection_2__14__3_, connection_2__14__2_, connection_2__14__1_, 
        connection_2__14__0_, connection_2__12__31_, connection_2__12__30_, 
        connection_2__12__29_, connection_2__12__28_, connection_2__12__27_, 
        connection_2__12__26_, connection_2__12__25_, connection_2__12__24_, 
        connection_2__12__23_, connection_2__12__22_, connection_2__12__21_, 
        connection_2__12__20_, connection_2__12__19_, connection_2__12__18_, 
        connection_2__12__17_, connection_2__12__16_, connection_2__12__15_, 
        connection_2__12__14_, connection_2__12__13_, connection_2__12__12_, 
        connection_2__12__11_, connection_2__12__10_, connection_2__12__9_, 
        connection_2__12__8_, connection_2__12__7_, connection_2__12__6_, 
        connection_2__12__5_, connection_2__12__4_, connection_2__12__3_, 
        connection_2__12__2_, connection_2__12__1_, connection_2__12__0_}), 
        .o_valid({connection_valid_3__11_, connection_valid_3__10_}), 
        .o_data_bus({connection_3__11__31_, connection_3__11__30_, 
        connection_3__11__29_, connection_3__11__28_, connection_3__11__27_, 
        connection_3__11__26_, connection_3__11__25_, connection_3__11__24_, 
        connection_3__11__23_, connection_3__11__22_, connection_3__11__21_, 
        connection_3__11__20_, connection_3__11__19_, connection_3__11__18_, 
        connection_3__11__17_, connection_3__11__16_, connection_3__11__15_, 
        connection_3__11__14_, connection_3__11__13_, connection_3__11__12_, 
        connection_3__11__11_, connection_3__11__10_, connection_3__11__9_, 
        connection_3__11__8_, connection_3__11__7_, connection_3__11__6_, 
        connection_3__11__5_, connection_3__11__4_, connection_3__11__3_, 
        connection_3__11__2_, connection_3__11__1_, connection_3__11__0_, 
        connection_3__10__31_, connection_3__10__30_, connection_3__10__29_, 
        connection_3__10__28_, connection_3__10__27_, connection_3__10__26_, 
        connection_3__10__25_, connection_3__10__24_, connection_3__10__23_, 
        connection_3__10__22_, connection_3__10__21_, connection_3__10__20_, 
        connection_3__10__19_, connection_3__10__18_, connection_3__10__17_, 
        connection_3__10__16_, connection_3__10__15_, connection_3__10__14_, 
        connection_3__10__13_, connection_3__10__12_, connection_3__10__11_, 
        connection_3__10__10_, connection_3__10__9_, connection_3__10__8_, 
        connection_3__10__7_, connection_3__10__6_, connection_3__10__5_, 
        connection_3__10__4_, connection_3__10__3_, connection_3__10__2_, 
        connection_3__10__1_, connection_3__10__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[181:180]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_90 first_half_stages_2__group_first_half_1__switch_first_half_2__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__11_, 
        connection_valid_2__9_}), .i_data_bus({connection_2__11__31_, 
        connection_2__11__30_, connection_2__11__29_, connection_2__11__28_, 
        connection_2__11__27_, connection_2__11__26_, connection_2__11__25_, 
        connection_2__11__24_, connection_2__11__23_, connection_2__11__22_, 
        connection_2__11__21_, connection_2__11__20_, connection_2__11__19_, 
        connection_2__11__18_, connection_2__11__17_, connection_2__11__16_, 
        connection_2__11__15_, connection_2__11__14_, connection_2__11__13_, 
        connection_2__11__12_, connection_2__11__11_, connection_2__11__10_, 
        connection_2__11__9_, connection_2__11__8_, connection_2__11__7_, 
        connection_2__11__6_, connection_2__11__5_, connection_2__11__4_, 
        connection_2__11__3_, connection_2__11__2_, connection_2__11__1_, 
        connection_2__11__0_, connection_2__9__31_, connection_2__9__30_, 
        connection_2__9__29_, connection_2__9__28_, connection_2__9__27_, 
        connection_2__9__26_, connection_2__9__25_, connection_2__9__24_, 
        connection_2__9__23_, connection_2__9__22_, connection_2__9__21_, 
        connection_2__9__20_, connection_2__9__19_, connection_2__9__18_, 
        connection_2__9__17_, connection_2__9__16_, connection_2__9__15_, 
        connection_2__9__14_, connection_2__9__13_, connection_2__9__12_, 
        connection_2__9__11_, connection_2__9__10_, connection_2__9__9_, 
        connection_2__9__8_, connection_2__9__7_, connection_2__9__6_, 
        connection_2__9__5_, connection_2__9__4_, connection_2__9__3_, 
        connection_2__9__2_, connection_2__9__1_, connection_2__9__0_}), 
        .o_valid({connection_valid_3__13_, connection_valid_3__12_}), 
        .o_data_bus({connection_3__13__31_, connection_3__13__30_, 
        connection_3__13__29_, connection_3__13__28_, connection_3__13__27_, 
        connection_3__13__26_, connection_3__13__25_, connection_3__13__24_, 
        connection_3__13__23_, connection_3__13__22_, connection_3__13__21_, 
        connection_3__13__20_, connection_3__13__19_, connection_3__13__18_, 
        connection_3__13__17_, connection_3__13__16_, connection_3__13__15_, 
        connection_3__13__14_, connection_3__13__13_, connection_3__13__12_, 
        connection_3__13__11_, connection_3__13__10_, connection_3__13__9_, 
        connection_3__13__8_, connection_3__13__7_, connection_3__13__6_, 
        connection_3__13__5_, connection_3__13__4_, connection_3__13__3_, 
        connection_3__13__2_, connection_3__13__1_, connection_3__13__0_, 
        connection_3__12__31_, connection_3__12__30_, connection_3__12__29_, 
        connection_3__12__28_, connection_3__12__27_, connection_3__12__26_, 
        connection_3__12__25_, connection_3__12__24_, connection_3__12__23_, 
        connection_3__12__22_, connection_3__12__21_, connection_3__12__20_, 
        connection_3__12__19_, connection_3__12__18_, connection_3__12__17_, 
        connection_3__12__16_, connection_3__12__15_, connection_3__12__14_, 
        connection_3__12__13_, connection_3__12__12_, connection_3__12__11_, 
        connection_3__12__10_, connection_3__12__9_, connection_3__12__8_, 
        connection_3__12__7_, connection_3__12__6_, connection_3__12__5_, 
        connection_3__12__4_, connection_3__12__3_, connection_3__12__2_, 
        connection_3__12__1_, connection_3__12__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[179:178]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_89 first_half_stages_2__group_first_half_1__switch_first_half_3__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__15_, 
        connection_valid_2__13_}), .i_data_bus({connection_2__15__31_, 
        connection_2__15__30_, connection_2__15__29_, connection_2__15__28_, 
        connection_2__15__27_, connection_2__15__26_, connection_2__15__25_, 
        connection_2__15__24_, connection_2__15__23_, connection_2__15__22_, 
        connection_2__15__21_, connection_2__15__20_, connection_2__15__19_, 
        connection_2__15__18_, connection_2__15__17_, connection_2__15__16_, 
        connection_2__15__15_, connection_2__15__14_, connection_2__15__13_, 
        connection_2__15__12_, connection_2__15__11_, connection_2__15__10_, 
        connection_2__15__9_, connection_2__15__8_, connection_2__15__7_, 
        connection_2__15__6_, connection_2__15__5_, connection_2__15__4_, 
        connection_2__15__3_, connection_2__15__2_, connection_2__15__1_, 
        connection_2__15__0_, connection_2__13__31_, connection_2__13__30_, 
        connection_2__13__29_, connection_2__13__28_, connection_2__13__27_, 
        connection_2__13__26_, connection_2__13__25_, connection_2__13__24_, 
        connection_2__13__23_, connection_2__13__22_, connection_2__13__21_, 
        connection_2__13__20_, connection_2__13__19_, connection_2__13__18_, 
        connection_2__13__17_, connection_2__13__16_, connection_2__13__15_, 
        connection_2__13__14_, connection_2__13__13_, connection_2__13__12_, 
        connection_2__13__11_, connection_2__13__10_, connection_2__13__9_, 
        connection_2__13__8_, connection_2__13__7_, connection_2__13__6_, 
        connection_2__13__5_, connection_2__13__4_, connection_2__13__3_, 
        connection_2__13__2_, connection_2__13__1_, connection_2__13__0_}), 
        .o_valid({connection_valid_3__15_, connection_valid_3__14_}), 
        .o_data_bus({connection_3__15__31_, connection_3__15__30_, 
        connection_3__15__29_, connection_3__15__28_, connection_3__15__27_, 
        connection_3__15__26_, connection_3__15__25_, connection_3__15__24_, 
        connection_3__15__23_, connection_3__15__22_, connection_3__15__21_, 
        connection_3__15__20_, connection_3__15__19_, connection_3__15__18_, 
        connection_3__15__17_, connection_3__15__16_, connection_3__15__15_, 
        connection_3__15__14_, connection_3__15__13_, connection_3__15__12_, 
        connection_3__15__11_, connection_3__15__10_, connection_3__15__9_, 
        connection_3__15__8_, connection_3__15__7_, connection_3__15__6_, 
        connection_3__15__5_, connection_3__15__4_, connection_3__15__3_, 
        connection_3__15__2_, connection_3__15__1_, connection_3__15__0_, 
        connection_3__14__31_, connection_3__14__30_, connection_3__14__29_, 
        connection_3__14__28_, connection_3__14__27_, connection_3__14__26_, 
        connection_3__14__25_, connection_3__14__24_, connection_3__14__23_, 
        connection_3__14__22_, connection_3__14__21_, connection_3__14__20_, 
        connection_3__14__19_, connection_3__14__18_, connection_3__14__17_, 
        connection_3__14__16_, connection_3__14__15_, connection_3__14__14_, 
        connection_3__14__13_, connection_3__14__12_, connection_3__14__11_, 
        connection_3__14__10_, connection_3__14__9_, connection_3__14__8_, 
        connection_3__14__7_, connection_3__14__6_, connection_3__14__5_, 
        connection_3__14__4_, connection_3__14__3_, connection_3__14__2_, 
        connection_3__14__1_, connection_3__14__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[177:176]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_88 first_half_stages_2__group_first_half_2__switch_first_half_0__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__18_, 
        connection_valid_2__16_}), .i_data_bus({connection_2__18__31_, 
        connection_2__18__30_, connection_2__18__29_, connection_2__18__28_, 
        connection_2__18__27_, connection_2__18__26_, connection_2__18__25_, 
        connection_2__18__24_, connection_2__18__23_, connection_2__18__22_, 
        connection_2__18__21_, connection_2__18__20_, connection_2__18__19_, 
        connection_2__18__18_, connection_2__18__17_, connection_2__18__16_, 
        connection_2__18__15_, connection_2__18__14_, connection_2__18__13_, 
        connection_2__18__12_, connection_2__18__11_, connection_2__18__10_, 
        connection_2__18__9_, connection_2__18__8_, connection_2__18__7_, 
        connection_2__18__6_, connection_2__18__5_, connection_2__18__4_, 
        connection_2__18__3_, connection_2__18__2_, connection_2__18__1_, 
        connection_2__18__0_, connection_2__16__31_, connection_2__16__30_, 
        connection_2__16__29_, connection_2__16__28_, connection_2__16__27_, 
        connection_2__16__26_, connection_2__16__25_, connection_2__16__24_, 
        connection_2__16__23_, connection_2__16__22_, connection_2__16__21_, 
        connection_2__16__20_, connection_2__16__19_, connection_2__16__18_, 
        connection_2__16__17_, connection_2__16__16_, connection_2__16__15_, 
        connection_2__16__14_, connection_2__16__13_, connection_2__16__12_, 
        connection_2__16__11_, connection_2__16__10_, connection_2__16__9_, 
        connection_2__16__8_, connection_2__16__7_, connection_2__16__6_, 
        connection_2__16__5_, connection_2__16__4_, connection_2__16__3_, 
        connection_2__16__2_, connection_2__16__1_, connection_2__16__0_}), 
        .o_valid({connection_valid_3__17_, connection_valid_3__16_}), 
        .o_data_bus({connection_3__17__31_, connection_3__17__30_, 
        connection_3__17__29_, connection_3__17__28_, connection_3__17__27_, 
        connection_3__17__26_, connection_3__17__25_, connection_3__17__24_, 
        connection_3__17__23_, connection_3__17__22_, connection_3__17__21_, 
        connection_3__17__20_, connection_3__17__19_, connection_3__17__18_, 
        connection_3__17__17_, connection_3__17__16_, connection_3__17__15_, 
        connection_3__17__14_, connection_3__17__13_, connection_3__17__12_, 
        connection_3__17__11_, connection_3__17__10_, connection_3__17__9_, 
        connection_3__17__8_, connection_3__17__7_, connection_3__17__6_, 
        connection_3__17__5_, connection_3__17__4_, connection_3__17__3_, 
        connection_3__17__2_, connection_3__17__1_, connection_3__17__0_, 
        connection_3__16__31_, connection_3__16__30_, connection_3__16__29_, 
        connection_3__16__28_, connection_3__16__27_, connection_3__16__26_, 
        connection_3__16__25_, connection_3__16__24_, connection_3__16__23_, 
        connection_3__16__22_, connection_3__16__21_, connection_3__16__20_, 
        connection_3__16__19_, connection_3__16__18_, connection_3__16__17_, 
        connection_3__16__16_, connection_3__16__15_, connection_3__16__14_, 
        connection_3__16__13_, connection_3__16__12_, connection_3__16__11_, 
        connection_3__16__10_, connection_3__16__9_, connection_3__16__8_, 
        connection_3__16__7_, connection_3__16__6_, connection_3__16__5_, 
        connection_3__16__4_, connection_3__16__3_, connection_3__16__2_, 
        connection_3__16__1_, connection_3__16__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[175:174]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_87 first_half_stages_2__group_first_half_2__switch_first_half_1__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__22_, 
        connection_valid_2__20_}), .i_data_bus({connection_2__22__31_, 
        connection_2__22__30_, connection_2__22__29_, connection_2__22__28_, 
        connection_2__22__27_, connection_2__22__26_, connection_2__22__25_, 
        connection_2__22__24_, connection_2__22__23_, connection_2__22__22_, 
        connection_2__22__21_, connection_2__22__20_, connection_2__22__19_, 
        connection_2__22__18_, connection_2__22__17_, connection_2__22__16_, 
        connection_2__22__15_, connection_2__22__14_, connection_2__22__13_, 
        connection_2__22__12_, connection_2__22__11_, connection_2__22__10_, 
        connection_2__22__9_, connection_2__22__8_, connection_2__22__7_, 
        connection_2__22__6_, connection_2__22__5_, connection_2__22__4_, 
        connection_2__22__3_, connection_2__22__2_, connection_2__22__1_, 
        connection_2__22__0_, connection_2__20__31_, connection_2__20__30_, 
        connection_2__20__29_, connection_2__20__28_, connection_2__20__27_, 
        connection_2__20__26_, connection_2__20__25_, connection_2__20__24_, 
        connection_2__20__23_, connection_2__20__22_, connection_2__20__21_, 
        connection_2__20__20_, connection_2__20__19_, connection_2__20__18_, 
        connection_2__20__17_, connection_2__20__16_, connection_2__20__15_, 
        connection_2__20__14_, connection_2__20__13_, connection_2__20__12_, 
        connection_2__20__11_, connection_2__20__10_, connection_2__20__9_, 
        connection_2__20__8_, connection_2__20__7_, connection_2__20__6_, 
        connection_2__20__5_, connection_2__20__4_, connection_2__20__3_, 
        connection_2__20__2_, connection_2__20__1_, connection_2__20__0_}), 
        .o_valid({connection_valid_3__19_, connection_valid_3__18_}), 
        .o_data_bus({connection_3__19__31_, connection_3__19__30_, 
        connection_3__19__29_, connection_3__19__28_, connection_3__19__27_, 
        connection_3__19__26_, connection_3__19__25_, connection_3__19__24_, 
        connection_3__19__23_, connection_3__19__22_, connection_3__19__21_, 
        connection_3__19__20_, connection_3__19__19_, connection_3__19__18_, 
        connection_3__19__17_, connection_3__19__16_, connection_3__19__15_, 
        connection_3__19__14_, connection_3__19__13_, connection_3__19__12_, 
        connection_3__19__11_, connection_3__19__10_, connection_3__19__9_, 
        connection_3__19__8_, connection_3__19__7_, connection_3__19__6_, 
        connection_3__19__5_, connection_3__19__4_, connection_3__19__3_, 
        connection_3__19__2_, connection_3__19__1_, connection_3__19__0_, 
        connection_3__18__31_, connection_3__18__30_, connection_3__18__29_, 
        connection_3__18__28_, connection_3__18__27_, connection_3__18__26_, 
        connection_3__18__25_, connection_3__18__24_, connection_3__18__23_, 
        connection_3__18__22_, connection_3__18__21_, connection_3__18__20_, 
        connection_3__18__19_, connection_3__18__18_, connection_3__18__17_, 
        connection_3__18__16_, connection_3__18__15_, connection_3__18__14_, 
        connection_3__18__13_, connection_3__18__12_, connection_3__18__11_, 
        connection_3__18__10_, connection_3__18__9_, connection_3__18__8_, 
        connection_3__18__7_, connection_3__18__6_, connection_3__18__5_, 
        connection_3__18__4_, connection_3__18__3_, connection_3__18__2_, 
        connection_3__18__1_, connection_3__18__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[173:172]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_86 first_half_stages_2__group_first_half_2__switch_first_half_2__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__19_, 
        connection_valid_2__17_}), .i_data_bus({connection_2__19__31_, 
        connection_2__19__30_, connection_2__19__29_, connection_2__19__28_, 
        connection_2__19__27_, connection_2__19__26_, connection_2__19__25_, 
        connection_2__19__24_, connection_2__19__23_, connection_2__19__22_, 
        connection_2__19__21_, connection_2__19__20_, connection_2__19__19_, 
        connection_2__19__18_, connection_2__19__17_, connection_2__19__16_, 
        connection_2__19__15_, connection_2__19__14_, connection_2__19__13_, 
        connection_2__19__12_, connection_2__19__11_, connection_2__19__10_, 
        connection_2__19__9_, connection_2__19__8_, connection_2__19__7_, 
        connection_2__19__6_, connection_2__19__5_, connection_2__19__4_, 
        connection_2__19__3_, connection_2__19__2_, connection_2__19__1_, 
        connection_2__19__0_, connection_2__17__31_, connection_2__17__30_, 
        connection_2__17__29_, connection_2__17__28_, connection_2__17__27_, 
        connection_2__17__26_, connection_2__17__25_, connection_2__17__24_, 
        connection_2__17__23_, connection_2__17__22_, connection_2__17__21_, 
        connection_2__17__20_, connection_2__17__19_, connection_2__17__18_, 
        connection_2__17__17_, connection_2__17__16_, connection_2__17__15_, 
        connection_2__17__14_, connection_2__17__13_, connection_2__17__12_, 
        connection_2__17__11_, connection_2__17__10_, connection_2__17__9_, 
        connection_2__17__8_, connection_2__17__7_, connection_2__17__6_, 
        connection_2__17__5_, connection_2__17__4_, connection_2__17__3_, 
        connection_2__17__2_, connection_2__17__1_, connection_2__17__0_}), 
        .o_valid({connection_valid_3__21_, connection_valid_3__20_}), 
        .o_data_bus({connection_3__21__31_, connection_3__21__30_, 
        connection_3__21__29_, connection_3__21__28_, connection_3__21__27_, 
        connection_3__21__26_, connection_3__21__25_, connection_3__21__24_, 
        connection_3__21__23_, connection_3__21__22_, connection_3__21__21_, 
        connection_3__21__20_, connection_3__21__19_, connection_3__21__18_, 
        connection_3__21__17_, connection_3__21__16_, connection_3__21__15_, 
        connection_3__21__14_, connection_3__21__13_, connection_3__21__12_, 
        connection_3__21__11_, connection_3__21__10_, connection_3__21__9_, 
        connection_3__21__8_, connection_3__21__7_, connection_3__21__6_, 
        connection_3__21__5_, connection_3__21__4_, connection_3__21__3_, 
        connection_3__21__2_, connection_3__21__1_, connection_3__21__0_, 
        connection_3__20__31_, connection_3__20__30_, connection_3__20__29_, 
        connection_3__20__28_, connection_3__20__27_, connection_3__20__26_, 
        connection_3__20__25_, connection_3__20__24_, connection_3__20__23_, 
        connection_3__20__22_, connection_3__20__21_, connection_3__20__20_, 
        connection_3__20__19_, connection_3__20__18_, connection_3__20__17_, 
        connection_3__20__16_, connection_3__20__15_, connection_3__20__14_, 
        connection_3__20__13_, connection_3__20__12_, connection_3__20__11_, 
        connection_3__20__10_, connection_3__20__9_, connection_3__20__8_, 
        connection_3__20__7_, connection_3__20__6_, connection_3__20__5_, 
        connection_3__20__4_, connection_3__20__3_, connection_3__20__2_, 
        connection_3__20__1_, connection_3__20__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[171:170]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_85 first_half_stages_2__group_first_half_2__switch_first_half_3__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__23_, 
        connection_valid_2__21_}), .i_data_bus({connection_2__23__31_, 
        connection_2__23__30_, connection_2__23__29_, connection_2__23__28_, 
        connection_2__23__27_, connection_2__23__26_, connection_2__23__25_, 
        connection_2__23__24_, connection_2__23__23_, connection_2__23__22_, 
        connection_2__23__21_, connection_2__23__20_, connection_2__23__19_, 
        connection_2__23__18_, connection_2__23__17_, connection_2__23__16_, 
        connection_2__23__15_, connection_2__23__14_, connection_2__23__13_, 
        connection_2__23__12_, connection_2__23__11_, connection_2__23__10_, 
        connection_2__23__9_, connection_2__23__8_, connection_2__23__7_, 
        connection_2__23__6_, connection_2__23__5_, connection_2__23__4_, 
        connection_2__23__3_, connection_2__23__2_, connection_2__23__1_, 
        connection_2__23__0_, connection_2__21__31_, connection_2__21__30_, 
        connection_2__21__29_, connection_2__21__28_, connection_2__21__27_, 
        connection_2__21__26_, connection_2__21__25_, connection_2__21__24_, 
        connection_2__21__23_, connection_2__21__22_, connection_2__21__21_, 
        connection_2__21__20_, connection_2__21__19_, connection_2__21__18_, 
        connection_2__21__17_, connection_2__21__16_, connection_2__21__15_, 
        connection_2__21__14_, connection_2__21__13_, connection_2__21__12_, 
        connection_2__21__11_, connection_2__21__10_, connection_2__21__9_, 
        connection_2__21__8_, connection_2__21__7_, connection_2__21__6_, 
        connection_2__21__5_, connection_2__21__4_, connection_2__21__3_, 
        connection_2__21__2_, connection_2__21__1_, connection_2__21__0_}), 
        .o_valid({connection_valid_3__23_, connection_valid_3__22_}), 
        .o_data_bus({connection_3__23__31_, connection_3__23__30_, 
        connection_3__23__29_, connection_3__23__28_, connection_3__23__27_, 
        connection_3__23__26_, connection_3__23__25_, connection_3__23__24_, 
        connection_3__23__23_, connection_3__23__22_, connection_3__23__21_, 
        connection_3__23__20_, connection_3__23__19_, connection_3__23__18_, 
        connection_3__23__17_, connection_3__23__16_, connection_3__23__15_, 
        connection_3__23__14_, connection_3__23__13_, connection_3__23__12_, 
        connection_3__23__11_, connection_3__23__10_, connection_3__23__9_, 
        connection_3__23__8_, connection_3__23__7_, connection_3__23__6_, 
        connection_3__23__5_, connection_3__23__4_, connection_3__23__3_, 
        connection_3__23__2_, connection_3__23__1_, connection_3__23__0_, 
        connection_3__22__31_, connection_3__22__30_, connection_3__22__29_, 
        connection_3__22__28_, connection_3__22__27_, connection_3__22__26_, 
        connection_3__22__25_, connection_3__22__24_, connection_3__22__23_, 
        connection_3__22__22_, connection_3__22__21_, connection_3__22__20_, 
        connection_3__22__19_, connection_3__22__18_, connection_3__22__17_, 
        connection_3__22__16_, connection_3__22__15_, connection_3__22__14_, 
        connection_3__22__13_, connection_3__22__12_, connection_3__22__11_, 
        connection_3__22__10_, connection_3__22__9_, connection_3__22__8_, 
        connection_3__22__7_, connection_3__22__6_, connection_3__22__5_, 
        connection_3__22__4_, connection_3__22__3_, connection_3__22__2_, 
        connection_3__22__1_, connection_3__22__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[169:168]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_84 first_half_stages_2__group_first_half_3__switch_first_half_0__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__26_, 
        connection_valid_2__24_}), .i_data_bus({connection_2__26__31_, 
        connection_2__26__30_, connection_2__26__29_, connection_2__26__28_, 
        connection_2__26__27_, connection_2__26__26_, connection_2__26__25_, 
        connection_2__26__24_, connection_2__26__23_, connection_2__26__22_, 
        connection_2__26__21_, connection_2__26__20_, connection_2__26__19_, 
        connection_2__26__18_, connection_2__26__17_, connection_2__26__16_, 
        connection_2__26__15_, connection_2__26__14_, connection_2__26__13_, 
        connection_2__26__12_, connection_2__26__11_, connection_2__26__10_, 
        connection_2__26__9_, connection_2__26__8_, connection_2__26__7_, 
        connection_2__26__6_, connection_2__26__5_, connection_2__26__4_, 
        connection_2__26__3_, connection_2__26__2_, connection_2__26__1_, 
        connection_2__26__0_, connection_2__24__31_, connection_2__24__30_, 
        connection_2__24__29_, connection_2__24__28_, connection_2__24__27_, 
        connection_2__24__26_, connection_2__24__25_, connection_2__24__24_, 
        connection_2__24__23_, connection_2__24__22_, connection_2__24__21_, 
        connection_2__24__20_, connection_2__24__19_, connection_2__24__18_, 
        connection_2__24__17_, connection_2__24__16_, connection_2__24__15_, 
        connection_2__24__14_, connection_2__24__13_, connection_2__24__12_, 
        connection_2__24__11_, connection_2__24__10_, connection_2__24__9_, 
        connection_2__24__8_, connection_2__24__7_, connection_2__24__6_, 
        connection_2__24__5_, connection_2__24__4_, connection_2__24__3_, 
        connection_2__24__2_, connection_2__24__1_, connection_2__24__0_}), 
        .o_valid({connection_valid_3__25_, connection_valid_3__24_}), 
        .o_data_bus({connection_3__25__31_, connection_3__25__30_, 
        connection_3__25__29_, connection_3__25__28_, connection_3__25__27_, 
        connection_3__25__26_, connection_3__25__25_, connection_3__25__24_, 
        connection_3__25__23_, connection_3__25__22_, connection_3__25__21_, 
        connection_3__25__20_, connection_3__25__19_, connection_3__25__18_, 
        connection_3__25__17_, connection_3__25__16_, connection_3__25__15_, 
        connection_3__25__14_, connection_3__25__13_, connection_3__25__12_, 
        connection_3__25__11_, connection_3__25__10_, connection_3__25__9_, 
        connection_3__25__8_, connection_3__25__7_, connection_3__25__6_, 
        connection_3__25__5_, connection_3__25__4_, connection_3__25__3_, 
        connection_3__25__2_, connection_3__25__1_, connection_3__25__0_, 
        connection_3__24__31_, connection_3__24__30_, connection_3__24__29_, 
        connection_3__24__28_, connection_3__24__27_, connection_3__24__26_, 
        connection_3__24__25_, connection_3__24__24_, connection_3__24__23_, 
        connection_3__24__22_, connection_3__24__21_, connection_3__24__20_, 
        connection_3__24__19_, connection_3__24__18_, connection_3__24__17_, 
        connection_3__24__16_, connection_3__24__15_, connection_3__24__14_, 
        connection_3__24__13_, connection_3__24__12_, connection_3__24__11_, 
        connection_3__24__10_, connection_3__24__9_, connection_3__24__8_, 
        connection_3__24__7_, connection_3__24__6_, connection_3__24__5_, 
        connection_3__24__4_, connection_3__24__3_, connection_3__24__2_, 
        connection_3__24__1_, connection_3__24__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[167:166]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_83 first_half_stages_2__group_first_half_3__switch_first_half_1__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__30_, 
        connection_valid_2__28_}), .i_data_bus({connection_2__30__31_, 
        connection_2__30__30_, connection_2__30__29_, connection_2__30__28_, 
        connection_2__30__27_, connection_2__30__26_, connection_2__30__25_, 
        connection_2__30__24_, connection_2__30__23_, connection_2__30__22_, 
        connection_2__30__21_, connection_2__30__20_, connection_2__30__19_, 
        connection_2__30__18_, connection_2__30__17_, connection_2__30__16_, 
        connection_2__30__15_, connection_2__30__14_, connection_2__30__13_, 
        connection_2__30__12_, connection_2__30__11_, connection_2__30__10_, 
        connection_2__30__9_, connection_2__30__8_, connection_2__30__7_, 
        connection_2__30__6_, connection_2__30__5_, connection_2__30__4_, 
        connection_2__30__3_, connection_2__30__2_, connection_2__30__1_, 
        connection_2__30__0_, connection_2__28__31_, connection_2__28__30_, 
        connection_2__28__29_, connection_2__28__28_, connection_2__28__27_, 
        connection_2__28__26_, connection_2__28__25_, connection_2__28__24_, 
        connection_2__28__23_, connection_2__28__22_, connection_2__28__21_, 
        connection_2__28__20_, connection_2__28__19_, connection_2__28__18_, 
        connection_2__28__17_, connection_2__28__16_, connection_2__28__15_, 
        connection_2__28__14_, connection_2__28__13_, connection_2__28__12_, 
        connection_2__28__11_, connection_2__28__10_, connection_2__28__9_, 
        connection_2__28__8_, connection_2__28__7_, connection_2__28__6_, 
        connection_2__28__5_, connection_2__28__4_, connection_2__28__3_, 
        connection_2__28__2_, connection_2__28__1_, connection_2__28__0_}), 
        .o_valid({connection_valid_3__27_, connection_valid_3__26_}), 
        .o_data_bus({connection_3__27__31_, connection_3__27__30_, 
        connection_3__27__29_, connection_3__27__28_, connection_3__27__27_, 
        connection_3__27__26_, connection_3__27__25_, connection_3__27__24_, 
        connection_3__27__23_, connection_3__27__22_, connection_3__27__21_, 
        connection_3__27__20_, connection_3__27__19_, connection_3__27__18_, 
        connection_3__27__17_, connection_3__27__16_, connection_3__27__15_, 
        connection_3__27__14_, connection_3__27__13_, connection_3__27__12_, 
        connection_3__27__11_, connection_3__27__10_, connection_3__27__9_, 
        connection_3__27__8_, connection_3__27__7_, connection_3__27__6_, 
        connection_3__27__5_, connection_3__27__4_, connection_3__27__3_, 
        connection_3__27__2_, connection_3__27__1_, connection_3__27__0_, 
        connection_3__26__31_, connection_3__26__30_, connection_3__26__29_, 
        connection_3__26__28_, connection_3__26__27_, connection_3__26__26_, 
        connection_3__26__25_, connection_3__26__24_, connection_3__26__23_, 
        connection_3__26__22_, connection_3__26__21_, connection_3__26__20_, 
        connection_3__26__19_, connection_3__26__18_, connection_3__26__17_, 
        connection_3__26__16_, connection_3__26__15_, connection_3__26__14_, 
        connection_3__26__13_, connection_3__26__12_, connection_3__26__11_, 
        connection_3__26__10_, connection_3__26__9_, connection_3__26__8_, 
        connection_3__26__7_, connection_3__26__6_, connection_3__26__5_, 
        connection_3__26__4_, connection_3__26__3_, connection_3__26__2_, 
        connection_3__26__1_, connection_3__26__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[165:164]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_82 first_half_stages_2__group_first_half_3__switch_first_half_2__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__27_, 
        connection_valid_2__25_}), .i_data_bus({connection_2__27__31_, 
        connection_2__27__30_, connection_2__27__29_, connection_2__27__28_, 
        connection_2__27__27_, connection_2__27__26_, connection_2__27__25_, 
        connection_2__27__24_, connection_2__27__23_, connection_2__27__22_, 
        connection_2__27__21_, connection_2__27__20_, connection_2__27__19_, 
        connection_2__27__18_, connection_2__27__17_, connection_2__27__16_, 
        connection_2__27__15_, connection_2__27__14_, connection_2__27__13_, 
        connection_2__27__12_, connection_2__27__11_, connection_2__27__10_, 
        connection_2__27__9_, connection_2__27__8_, connection_2__27__7_, 
        connection_2__27__6_, connection_2__27__5_, connection_2__27__4_, 
        connection_2__27__3_, connection_2__27__2_, connection_2__27__1_, 
        connection_2__27__0_, connection_2__25__31_, connection_2__25__30_, 
        connection_2__25__29_, connection_2__25__28_, connection_2__25__27_, 
        connection_2__25__26_, connection_2__25__25_, connection_2__25__24_, 
        connection_2__25__23_, connection_2__25__22_, connection_2__25__21_, 
        connection_2__25__20_, connection_2__25__19_, connection_2__25__18_, 
        connection_2__25__17_, connection_2__25__16_, connection_2__25__15_, 
        connection_2__25__14_, connection_2__25__13_, connection_2__25__12_, 
        connection_2__25__11_, connection_2__25__10_, connection_2__25__9_, 
        connection_2__25__8_, connection_2__25__7_, connection_2__25__6_, 
        connection_2__25__5_, connection_2__25__4_, connection_2__25__3_, 
        connection_2__25__2_, connection_2__25__1_, connection_2__25__0_}), 
        .o_valid({connection_valid_3__29_, connection_valid_3__28_}), 
        .o_data_bus({connection_3__29__31_, connection_3__29__30_, 
        connection_3__29__29_, connection_3__29__28_, connection_3__29__27_, 
        connection_3__29__26_, connection_3__29__25_, connection_3__29__24_, 
        connection_3__29__23_, connection_3__29__22_, connection_3__29__21_, 
        connection_3__29__20_, connection_3__29__19_, connection_3__29__18_, 
        connection_3__29__17_, connection_3__29__16_, connection_3__29__15_, 
        connection_3__29__14_, connection_3__29__13_, connection_3__29__12_, 
        connection_3__29__11_, connection_3__29__10_, connection_3__29__9_, 
        connection_3__29__8_, connection_3__29__7_, connection_3__29__6_, 
        connection_3__29__5_, connection_3__29__4_, connection_3__29__3_, 
        connection_3__29__2_, connection_3__29__1_, connection_3__29__0_, 
        connection_3__28__31_, connection_3__28__30_, connection_3__28__29_, 
        connection_3__28__28_, connection_3__28__27_, connection_3__28__26_, 
        connection_3__28__25_, connection_3__28__24_, connection_3__28__23_, 
        connection_3__28__22_, connection_3__28__21_, connection_3__28__20_, 
        connection_3__28__19_, connection_3__28__18_, connection_3__28__17_, 
        connection_3__28__16_, connection_3__28__15_, connection_3__28__14_, 
        connection_3__28__13_, connection_3__28__12_, connection_3__28__11_, 
        connection_3__28__10_, connection_3__28__9_, connection_3__28__8_, 
        connection_3__28__7_, connection_3__28__6_, connection_3__28__5_, 
        connection_3__28__4_, connection_3__28__3_, connection_3__28__2_, 
        connection_3__28__1_, connection_3__28__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[163:162]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_81 first_half_stages_2__group_first_half_3__switch_first_half_3__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__31_, 
        connection_valid_2__29_}), .i_data_bus({connection_2__31__31_, 
        connection_2__31__30_, connection_2__31__29_, connection_2__31__28_, 
        connection_2__31__27_, connection_2__31__26_, connection_2__31__25_, 
        connection_2__31__24_, connection_2__31__23_, connection_2__31__22_, 
        connection_2__31__21_, connection_2__31__20_, connection_2__31__19_, 
        connection_2__31__18_, connection_2__31__17_, connection_2__31__16_, 
        connection_2__31__15_, connection_2__31__14_, connection_2__31__13_, 
        connection_2__31__12_, connection_2__31__11_, connection_2__31__10_, 
        connection_2__31__9_, connection_2__31__8_, connection_2__31__7_, 
        connection_2__31__6_, connection_2__31__5_, connection_2__31__4_, 
        connection_2__31__3_, connection_2__31__2_, connection_2__31__1_, 
        connection_2__31__0_, connection_2__29__31_, connection_2__29__30_, 
        connection_2__29__29_, connection_2__29__28_, connection_2__29__27_, 
        connection_2__29__26_, connection_2__29__25_, connection_2__29__24_, 
        connection_2__29__23_, connection_2__29__22_, connection_2__29__21_, 
        connection_2__29__20_, connection_2__29__19_, connection_2__29__18_, 
        connection_2__29__17_, connection_2__29__16_, connection_2__29__15_, 
        connection_2__29__14_, connection_2__29__13_, connection_2__29__12_, 
        connection_2__29__11_, connection_2__29__10_, connection_2__29__9_, 
        connection_2__29__8_, connection_2__29__7_, connection_2__29__6_, 
        connection_2__29__5_, connection_2__29__4_, connection_2__29__3_, 
        connection_2__29__2_, connection_2__29__1_, connection_2__29__0_}), 
        .o_valid({connection_valid_3__31_, connection_valid_3__30_}), 
        .o_data_bus({connection_3__31__31_, connection_3__31__30_, 
        connection_3__31__29_, connection_3__31__28_, connection_3__31__27_, 
        connection_3__31__26_, connection_3__31__25_, connection_3__31__24_, 
        connection_3__31__23_, connection_3__31__22_, connection_3__31__21_, 
        connection_3__31__20_, connection_3__31__19_, connection_3__31__18_, 
        connection_3__31__17_, connection_3__31__16_, connection_3__31__15_, 
        connection_3__31__14_, connection_3__31__13_, connection_3__31__12_, 
        connection_3__31__11_, connection_3__31__10_, connection_3__31__9_, 
        connection_3__31__8_, connection_3__31__7_, connection_3__31__6_, 
        connection_3__31__5_, connection_3__31__4_, connection_3__31__3_, 
        connection_3__31__2_, connection_3__31__1_, connection_3__31__0_, 
        connection_3__30__31_, connection_3__30__30_, connection_3__30__29_, 
        connection_3__30__28_, connection_3__30__27_, connection_3__30__26_, 
        connection_3__30__25_, connection_3__30__24_, connection_3__30__23_, 
        connection_3__30__22_, connection_3__30__21_, connection_3__30__20_, 
        connection_3__30__19_, connection_3__30__18_, connection_3__30__17_, 
        connection_3__30__16_, connection_3__30__15_, connection_3__30__14_, 
        connection_3__30__13_, connection_3__30__12_, connection_3__30__11_, 
        connection_3__30__10_, connection_3__30__9_, connection_3__30__8_, 
        connection_3__30__7_, connection_3__30__6_, connection_3__30__5_, 
        connection_3__30__4_, connection_3__30__3_, connection_3__30__2_, 
        connection_3__30__1_, connection_3__30__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[161:160]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_80 first_half_stages_3__group_first_half_0__switch_first_half_0__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__2_, 
        connection_valid_3__0_}), .i_data_bus({connection_3__2__31_, 
        connection_3__2__30_, connection_3__2__29_, connection_3__2__28_, 
        connection_3__2__27_, connection_3__2__26_, connection_3__2__25_, 
        connection_3__2__24_, connection_3__2__23_, connection_3__2__22_, 
        connection_3__2__21_, connection_3__2__20_, connection_3__2__19_, 
        connection_3__2__18_, connection_3__2__17_, connection_3__2__16_, 
        connection_3__2__15_, connection_3__2__14_, connection_3__2__13_, 
        connection_3__2__12_, connection_3__2__11_, connection_3__2__10_, 
        connection_3__2__9_, connection_3__2__8_, connection_3__2__7_, 
        connection_3__2__6_, connection_3__2__5_, connection_3__2__4_, 
        connection_3__2__3_, connection_3__2__2_, connection_3__2__1_, 
        connection_3__2__0_, connection_3__0__31_, connection_3__0__30_, 
        connection_3__0__29_, connection_3__0__28_, connection_3__0__27_, 
        connection_3__0__26_, connection_3__0__25_, connection_3__0__24_, 
        connection_3__0__23_, connection_3__0__22_, connection_3__0__21_, 
        connection_3__0__20_, connection_3__0__19_, connection_3__0__18_, 
        connection_3__0__17_, connection_3__0__16_, connection_3__0__15_, 
        connection_3__0__14_, connection_3__0__13_, connection_3__0__12_, 
        connection_3__0__11_, connection_3__0__10_, connection_3__0__9_, 
        connection_3__0__8_, connection_3__0__7_, connection_3__0__6_, 
        connection_3__0__5_, connection_3__0__4_, connection_3__0__3_, 
        connection_3__0__2_, connection_3__0__1_, connection_3__0__0_}), 
        .o_valid({connection_valid_4__1_, connection_valid_4__0_}), 
        .o_data_bus({connection_4__1__31_, connection_4__1__30_, 
        connection_4__1__29_, connection_4__1__28_, connection_4__1__27_, 
        connection_4__1__26_, connection_4__1__25_, connection_4__1__24_, 
        connection_4__1__23_, connection_4__1__22_, connection_4__1__21_, 
        connection_4__1__20_, connection_4__1__19_, connection_4__1__18_, 
        connection_4__1__17_, connection_4__1__16_, connection_4__1__15_, 
        connection_4__1__14_, connection_4__1__13_, connection_4__1__12_, 
        connection_4__1__11_, connection_4__1__10_, connection_4__1__9_, 
        connection_4__1__8_, connection_4__1__7_, connection_4__1__6_, 
        connection_4__1__5_, connection_4__1__4_, connection_4__1__3_, 
        connection_4__1__2_, connection_4__1__1_, connection_4__1__0_, 
        connection_4__0__31_, connection_4__0__30_, connection_4__0__29_, 
        connection_4__0__28_, connection_4__0__27_, connection_4__0__26_, 
        connection_4__0__25_, connection_4__0__24_, connection_4__0__23_, 
        connection_4__0__22_, connection_4__0__21_, connection_4__0__20_, 
        connection_4__0__19_, connection_4__0__18_, connection_4__0__17_, 
        connection_4__0__16_, connection_4__0__15_, connection_4__0__14_, 
        connection_4__0__13_, connection_4__0__12_, connection_4__0__11_, 
        connection_4__0__10_, connection_4__0__9_, connection_4__0__8_, 
        connection_4__0__7_, connection_4__0__6_, connection_4__0__5_, 
        connection_4__0__4_, connection_4__0__3_, connection_4__0__2_, 
        connection_4__0__1_, connection_4__0__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[159:158]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_79 first_half_stages_3__group_first_half_0__switch_first_half_1__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__3_, 
        connection_valid_3__1_}), .i_data_bus({connection_3__3__31_, 
        connection_3__3__30_, connection_3__3__29_, connection_3__3__28_, 
        connection_3__3__27_, connection_3__3__26_, connection_3__3__25_, 
        connection_3__3__24_, connection_3__3__23_, connection_3__3__22_, 
        connection_3__3__21_, connection_3__3__20_, connection_3__3__19_, 
        connection_3__3__18_, connection_3__3__17_, connection_3__3__16_, 
        connection_3__3__15_, connection_3__3__14_, connection_3__3__13_, 
        connection_3__3__12_, connection_3__3__11_, connection_3__3__10_, 
        connection_3__3__9_, connection_3__3__8_, connection_3__3__7_, 
        connection_3__3__6_, connection_3__3__5_, connection_3__3__4_, 
        connection_3__3__3_, connection_3__3__2_, connection_3__3__1_, 
        connection_3__3__0_, connection_3__1__31_, connection_3__1__30_, 
        connection_3__1__29_, connection_3__1__28_, connection_3__1__27_, 
        connection_3__1__26_, connection_3__1__25_, connection_3__1__24_, 
        connection_3__1__23_, connection_3__1__22_, connection_3__1__21_, 
        connection_3__1__20_, connection_3__1__19_, connection_3__1__18_, 
        connection_3__1__17_, connection_3__1__16_, connection_3__1__15_, 
        connection_3__1__14_, connection_3__1__13_, connection_3__1__12_, 
        connection_3__1__11_, connection_3__1__10_, connection_3__1__9_, 
        connection_3__1__8_, connection_3__1__7_, connection_3__1__6_, 
        connection_3__1__5_, connection_3__1__4_, connection_3__1__3_, 
        connection_3__1__2_, connection_3__1__1_, connection_3__1__0_}), 
        .o_valid({connection_valid_4__3_, connection_valid_4__2_}), 
        .o_data_bus({connection_4__3__31_, connection_4__3__30_, 
        connection_4__3__29_, connection_4__3__28_, connection_4__3__27_, 
        connection_4__3__26_, connection_4__3__25_, connection_4__3__24_, 
        connection_4__3__23_, connection_4__3__22_, connection_4__3__21_, 
        connection_4__3__20_, connection_4__3__19_, connection_4__3__18_, 
        connection_4__3__17_, connection_4__3__16_, connection_4__3__15_, 
        connection_4__3__14_, connection_4__3__13_, connection_4__3__12_, 
        connection_4__3__11_, connection_4__3__10_, connection_4__3__9_, 
        connection_4__3__8_, connection_4__3__7_, connection_4__3__6_, 
        connection_4__3__5_, connection_4__3__4_, connection_4__3__3_, 
        connection_4__3__2_, connection_4__3__1_, connection_4__3__0_, 
        connection_4__2__31_, connection_4__2__30_, connection_4__2__29_, 
        connection_4__2__28_, connection_4__2__27_, connection_4__2__26_, 
        connection_4__2__25_, connection_4__2__24_, connection_4__2__23_, 
        connection_4__2__22_, connection_4__2__21_, connection_4__2__20_, 
        connection_4__2__19_, connection_4__2__18_, connection_4__2__17_, 
        connection_4__2__16_, connection_4__2__15_, connection_4__2__14_, 
        connection_4__2__13_, connection_4__2__12_, connection_4__2__11_, 
        connection_4__2__10_, connection_4__2__9_, connection_4__2__8_, 
        connection_4__2__7_, connection_4__2__6_, connection_4__2__5_, 
        connection_4__2__4_, connection_4__2__3_, connection_4__2__2_, 
        connection_4__2__1_, connection_4__2__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[157:156]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_78 first_half_stages_3__group_first_half_1__switch_first_half_0__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__6_, 
        connection_valid_3__4_}), .i_data_bus({connection_3__6__31_, 
        connection_3__6__30_, connection_3__6__29_, connection_3__6__28_, 
        connection_3__6__27_, connection_3__6__26_, connection_3__6__25_, 
        connection_3__6__24_, connection_3__6__23_, connection_3__6__22_, 
        connection_3__6__21_, connection_3__6__20_, connection_3__6__19_, 
        connection_3__6__18_, connection_3__6__17_, connection_3__6__16_, 
        connection_3__6__15_, connection_3__6__14_, connection_3__6__13_, 
        connection_3__6__12_, connection_3__6__11_, connection_3__6__10_, 
        connection_3__6__9_, connection_3__6__8_, connection_3__6__7_, 
        connection_3__6__6_, connection_3__6__5_, connection_3__6__4_, 
        connection_3__6__3_, connection_3__6__2_, connection_3__6__1_, 
        connection_3__6__0_, connection_3__4__31_, connection_3__4__30_, 
        connection_3__4__29_, connection_3__4__28_, connection_3__4__27_, 
        connection_3__4__26_, connection_3__4__25_, connection_3__4__24_, 
        connection_3__4__23_, connection_3__4__22_, connection_3__4__21_, 
        connection_3__4__20_, connection_3__4__19_, connection_3__4__18_, 
        connection_3__4__17_, connection_3__4__16_, connection_3__4__15_, 
        connection_3__4__14_, connection_3__4__13_, connection_3__4__12_, 
        connection_3__4__11_, connection_3__4__10_, connection_3__4__9_, 
        connection_3__4__8_, connection_3__4__7_, connection_3__4__6_, 
        connection_3__4__5_, connection_3__4__4_, connection_3__4__3_, 
        connection_3__4__2_, connection_3__4__1_, connection_3__4__0_}), 
        .o_valid({connection_valid_4__5_, connection_valid_4__4_}), 
        .o_data_bus({connection_4__5__31_, connection_4__5__30_, 
        connection_4__5__29_, connection_4__5__28_, connection_4__5__27_, 
        connection_4__5__26_, connection_4__5__25_, connection_4__5__24_, 
        connection_4__5__23_, connection_4__5__22_, connection_4__5__21_, 
        connection_4__5__20_, connection_4__5__19_, connection_4__5__18_, 
        connection_4__5__17_, connection_4__5__16_, connection_4__5__15_, 
        connection_4__5__14_, connection_4__5__13_, connection_4__5__12_, 
        connection_4__5__11_, connection_4__5__10_, connection_4__5__9_, 
        connection_4__5__8_, connection_4__5__7_, connection_4__5__6_, 
        connection_4__5__5_, connection_4__5__4_, connection_4__5__3_, 
        connection_4__5__2_, connection_4__5__1_, connection_4__5__0_, 
        connection_4__4__31_, connection_4__4__30_, connection_4__4__29_, 
        connection_4__4__28_, connection_4__4__27_, connection_4__4__26_, 
        connection_4__4__25_, connection_4__4__24_, connection_4__4__23_, 
        connection_4__4__22_, connection_4__4__21_, connection_4__4__20_, 
        connection_4__4__19_, connection_4__4__18_, connection_4__4__17_, 
        connection_4__4__16_, connection_4__4__15_, connection_4__4__14_, 
        connection_4__4__13_, connection_4__4__12_, connection_4__4__11_, 
        connection_4__4__10_, connection_4__4__9_, connection_4__4__8_, 
        connection_4__4__7_, connection_4__4__6_, connection_4__4__5_, 
        connection_4__4__4_, connection_4__4__3_, connection_4__4__2_, 
        connection_4__4__1_, connection_4__4__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[155:154]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_77 first_half_stages_3__group_first_half_1__switch_first_half_1__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__7_, 
        connection_valid_3__5_}), .i_data_bus({connection_3__7__31_, 
        connection_3__7__30_, connection_3__7__29_, connection_3__7__28_, 
        connection_3__7__27_, connection_3__7__26_, connection_3__7__25_, 
        connection_3__7__24_, connection_3__7__23_, connection_3__7__22_, 
        connection_3__7__21_, connection_3__7__20_, connection_3__7__19_, 
        connection_3__7__18_, connection_3__7__17_, connection_3__7__16_, 
        connection_3__7__15_, connection_3__7__14_, connection_3__7__13_, 
        connection_3__7__12_, connection_3__7__11_, connection_3__7__10_, 
        connection_3__7__9_, connection_3__7__8_, connection_3__7__7_, 
        connection_3__7__6_, connection_3__7__5_, connection_3__7__4_, 
        connection_3__7__3_, connection_3__7__2_, connection_3__7__1_, 
        connection_3__7__0_, connection_3__5__31_, connection_3__5__30_, 
        connection_3__5__29_, connection_3__5__28_, connection_3__5__27_, 
        connection_3__5__26_, connection_3__5__25_, connection_3__5__24_, 
        connection_3__5__23_, connection_3__5__22_, connection_3__5__21_, 
        connection_3__5__20_, connection_3__5__19_, connection_3__5__18_, 
        connection_3__5__17_, connection_3__5__16_, connection_3__5__15_, 
        connection_3__5__14_, connection_3__5__13_, connection_3__5__12_, 
        connection_3__5__11_, connection_3__5__10_, connection_3__5__9_, 
        connection_3__5__8_, connection_3__5__7_, connection_3__5__6_, 
        connection_3__5__5_, connection_3__5__4_, connection_3__5__3_, 
        connection_3__5__2_, connection_3__5__1_, connection_3__5__0_}), 
        .o_valid({connection_valid_4__7_, connection_valid_4__6_}), 
        .o_data_bus({connection_4__7__31_, connection_4__7__30_, 
        connection_4__7__29_, connection_4__7__28_, connection_4__7__27_, 
        connection_4__7__26_, connection_4__7__25_, connection_4__7__24_, 
        connection_4__7__23_, connection_4__7__22_, connection_4__7__21_, 
        connection_4__7__20_, connection_4__7__19_, connection_4__7__18_, 
        connection_4__7__17_, connection_4__7__16_, connection_4__7__15_, 
        connection_4__7__14_, connection_4__7__13_, connection_4__7__12_, 
        connection_4__7__11_, connection_4__7__10_, connection_4__7__9_, 
        connection_4__7__8_, connection_4__7__7_, connection_4__7__6_, 
        connection_4__7__5_, connection_4__7__4_, connection_4__7__3_, 
        connection_4__7__2_, connection_4__7__1_, connection_4__7__0_, 
        connection_4__6__31_, connection_4__6__30_, connection_4__6__29_, 
        connection_4__6__28_, connection_4__6__27_, connection_4__6__26_, 
        connection_4__6__25_, connection_4__6__24_, connection_4__6__23_, 
        connection_4__6__22_, connection_4__6__21_, connection_4__6__20_, 
        connection_4__6__19_, connection_4__6__18_, connection_4__6__17_, 
        connection_4__6__16_, connection_4__6__15_, connection_4__6__14_, 
        connection_4__6__13_, connection_4__6__12_, connection_4__6__11_, 
        connection_4__6__10_, connection_4__6__9_, connection_4__6__8_, 
        connection_4__6__7_, connection_4__6__6_, connection_4__6__5_, 
        connection_4__6__4_, connection_4__6__3_, connection_4__6__2_, 
        connection_4__6__1_, connection_4__6__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[153:152]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_76 first_half_stages_3__group_first_half_2__switch_first_half_0__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__10_, 
        connection_valid_3__8_}), .i_data_bus({connection_3__10__31_, 
        connection_3__10__30_, connection_3__10__29_, connection_3__10__28_, 
        connection_3__10__27_, connection_3__10__26_, connection_3__10__25_, 
        connection_3__10__24_, connection_3__10__23_, connection_3__10__22_, 
        connection_3__10__21_, connection_3__10__20_, connection_3__10__19_, 
        connection_3__10__18_, connection_3__10__17_, connection_3__10__16_, 
        connection_3__10__15_, connection_3__10__14_, connection_3__10__13_, 
        connection_3__10__12_, connection_3__10__11_, connection_3__10__10_, 
        connection_3__10__9_, connection_3__10__8_, connection_3__10__7_, 
        connection_3__10__6_, connection_3__10__5_, connection_3__10__4_, 
        connection_3__10__3_, connection_3__10__2_, connection_3__10__1_, 
        connection_3__10__0_, connection_3__8__31_, connection_3__8__30_, 
        connection_3__8__29_, connection_3__8__28_, connection_3__8__27_, 
        connection_3__8__26_, connection_3__8__25_, connection_3__8__24_, 
        connection_3__8__23_, connection_3__8__22_, connection_3__8__21_, 
        connection_3__8__20_, connection_3__8__19_, connection_3__8__18_, 
        connection_3__8__17_, connection_3__8__16_, connection_3__8__15_, 
        connection_3__8__14_, connection_3__8__13_, connection_3__8__12_, 
        connection_3__8__11_, connection_3__8__10_, connection_3__8__9_, 
        connection_3__8__8_, connection_3__8__7_, connection_3__8__6_, 
        connection_3__8__5_, connection_3__8__4_, connection_3__8__3_, 
        connection_3__8__2_, connection_3__8__1_, connection_3__8__0_}), 
        .o_valid({connection_valid_4__9_, connection_valid_4__8_}), 
        .o_data_bus({connection_4__9__31_, connection_4__9__30_, 
        connection_4__9__29_, connection_4__9__28_, connection_4__9__27_, 
        connection_4__9__26_, connection_4__9__25_, connection_4__9__24_, 
        connection_4__9__23_, connection_4__9__22_, connection_4__9__21_, 
        connection_4__9__20_, connection_4__9__19_, connection_4__9__18_, 
        connection_4__9__17_, connection_4__9__16_, connection_4__9__15_, 
        connection_4__9__14_, connection_4__9__13_, connection_4__9__12_, 
        connection_4__9__11_, connection_4__9__10_, connection_4__9__9_, 
        connection_4__9__8_, connection_4__9__7_, connection_4__9__6_, 
        connection_4__9__5_, connection_4__9__4_, connection_4__9__3_, 
        connection_4__9__2_, connection_4__9__1_, connection_4__9__0_, 
        connection_4__8__31_, connection_4__8__30_, connection_4__8__29_, 
        connection_4__8__28_, connection_4__8__27_, connection_4__8__26_, 
        connection_4__8__25_, connection_4__8__24_, connection_4__8__23_, 
        connection_4__8__22_, connection_4__8__21_, connection_4__8__20_, 
        connection_4__8__19_, connection_4__8__18_, connection_4__8__17_, 
        connection_4__8__16_, connection_4__8__15_, connection_4__8__14_, 
        connection_4__8__13_, connection_4__8__12_, connection_4__8__11_, 
        connection_4__8__10_, connection_4__8__9_, connection_4__8__8_, 
        connection_4__8__7_, connection_4__8__6_, connection_4__8__5_, 
        connection_4__8__4_, connection_4__8__3_, connection_4__8__2_, 
        connection_4__8__1_, connection_4__8__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[151:150]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_75 first_half_stages_3__group_first_half_2__switch_first_half_1__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__11_, 
        connection_valid_3__9_}), .i_data_bus({connection_3__11__31_, 
        connection_3__11__30_, connection_3__11__29_, connection_3__11__28_, 
        connection_3__11__27_, connection_3__11__26_, connection_3__11__25_, 
        connection_3__11__24_, connection_3__11__23_, connection_3__11__22_, 
        connection_3__11__21_, connection_3__11__20_, connection_3__11__19_, 
        connection_3__11__18_, connection_3__11__17_, connection_3__11__16_, 
        connection_3__11__15_, connection_3__11__14_, connection_3__11__13_, 
        connection_3__11__12_, connection_3__11__11_, connection_3__11__10_, 
        connection_3__11__9_, connection_3__11__8_, connection_3__11__7_, 
        connection_3__11__6_, connection_3__11__5_, connection_3__11__4_, 
        connection_3__11__3_, connection_3__11__2_, connection_3__11__1_, 
        connection_3__11__0_, connection_3__9__31_, connection_3__9__30_, 
        connection_3__9__29_, connection_3__9__28_, connection_3__9__27_, 
        connection_3__9__26_, connection_3__9__25_, connection_3__9__24_, 
        connection_3__9__23_, connection_3__9__22_, connection_3__9__21_, 
        connection_3__9__20_, connection_3__9__19_, connection_3__9__18_, 
        connection_3__9__17_, connection_3__9__16_, connection_3__9__15_, 
        connection_3__9__14_, connection_3__9__13_, connection_3__9__12_, 
        connection_3__9__11_, connection_3__9__10_, connection_3__9__9_, 
        connection_3__9__8_, connection_3__9__7_, connection_3__9__6_, 
        connection_3__9__5_, connection_3__9__4_, connection_3__9__3_, 
        connection_3__9__2_, connection_3__9__1_, connection_3__9__0_}), 
        .o_valid({connection_valid_4__11_, connection_valid_4__10_}), 
        .o_data_bus({connection_4__11__31_, connection_4__11__30_, 
        connection_4__11__29_, connection_4__11__28_, connection_4__11__27_, 
        connection_4__11__26_, connection_4__11__25_, connection_4__11__24_, 
        connection_4__11__23_, connection_4__11__22_, connection_4__11__21_, 
        connection_4__11__20_, connection_4__11__19_, connection_4__11__18_, 
        connection_4__11__17_, connection_4__11__16_, connection_4__11__15_, 
        connection_4__11__14_, connection_4__11__13_, connection_4__11__12_, 
        connection_4__11__11_, connection_4__11__10_, connection_4__11__9_, 
        connection_4__11__8_, connection_4__11__7_, connection_4__11__6_, 
        connection_4__11__5_, connection_4__11__4_, connection_4__11__3_, 
        connection_4__11__2_, connection_4__11__1_, connection_4__11__0_, 
        connection_4__10__31_, connection_4__10__30_, connection_4__10__29_, 
        connection_4__10__28_, connection_4__10__27_, connection_4__10__26_, 
        connection_4__10__25_, connection_4__10__24_, connection_4__10__23_, 
        connection_4__10__22_, connection_4__10__21_, connection_4__10__20_, 
        connection_4__10__19_, connection_4__10__18_, connection_4__10__17_, 
        connection_4__10__16_, connection_4__10__15_, connection_4__10__14_, 
        connection_4__10__13_, connection_4__10__12_, connection_4__10__11_, 
        connection_4__10__10_, connection_4__10__9_, connection_4__10__8_, 
        connection_4__10__7_, connection_4__10__6_, connection_4__10__5_, 
        connection_4__10__4_, connection_4__10__3_, connection_4__10__2_, 
        connection_4__10__1_, connection_4__10__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[149:148]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_74 first_half_stages_3__group_first_half_3__switch_first_half_0__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__14_, 
        connection_valid_3__12_}), .i_data_bus({connection_3__14__31_, 
        connection_3__14__30_, connection_3__14__29_, connection_3__14__28_, 
        connection_3__14__27_, connection_3__14__26_, connection_3__14__25_, 
        connection_3__14__24_, connection_3__14__23_, connection_3__14__22_, 
        connection_3__14__21_, connection_3__14__20_, connection_3__14__19_, 
        connection_3__14__18_, connection_3__14__17_, connection_3__14__16_, 
        connection_3__14__15_, connection_3__14__14_, connection_3__14__13_, 
        connection_3__14__12_, connection_3__14__11_, connection_3__14__10_, 
        connection_3__14__9_, connection_3__14__8_, connection_3__14__7_, 
        connection_3__14__6_, connection_3__14__5_, connection_3__14__4_, 
        connection_3__14__3_, connection_3__14__2_, connection_3__14__1_, 
        connection_3__14__0_, connection_3__12__31_, connection_3__12__30_, 
        connection_3__12__29_, connection_3__12__28_, connection_3__12__27_, 
        connection_3__12__26_, connection_3__12__25_, connection_3__12__24_, 
        connection_3__12__23_, connection_3__12__22_, connection_3__12__21_, 
        connection_3__12__20_, connection_3__12__19_, connection_3__12__18_, 
        connection_3__12__17_, connection_3__12__16_, connection_3__12__15_, 
        connection_3__12__14_, connection_3__12__13_, connection_3__12__12_, 
        connection_3__12__11_, connection_3__12__10_, connection_3__12__9_, 
        connection_3__12__8_, connection_3__12__7_, connection_3__12__6_, 
        connection_3__12__5_, connection_3__12__4_, connection_3__12__3_, 
        connection_3__12__2_, connection_3__12__1_, connection_3__12__0_}), 
        .o_valid({connection_valid_4__13_, connection_valid_4__12_}), 
        .o_data_bus({connection_4__13__31_, connection_4__13__30_, 
        connection_4__13__29_, connection_4__13__28_, connection_4__13__27_, 
        connection_4__13__26_, connection_4__13__25_, connection_4__13__24_, 
        connection_4__13__23_, connection_4__13__22_, connection_4__13__21_, 
        connection_4__13__20_, connection_4__13__19_, connection_4__13__18_, 
        connection_4__13__17_, connection_4__13__16_, connection_4__13__15_, 
        connection_4__13__14_, connection_4__13__13_, connection_4__13__12_, 
        connection_4__13__11_, connection_4__13__10_, connection_4__13__9_, 
        connection_4__13__8_, connection_4__13__7_, connection_4__13__6_, 
        connection_4__13__5_, connection_4__13__4_, connection_4__13__3_, 
        connection_4__13__2_, connection_4__13__1_, connection_4__13__0_, 
        connection_4__12__31_, connection_4__12__30_, connection_4__12__29_, 
        connection_4__12__28_, connection_4__12__27_, connection_4__12__26_, 
        connection_4__12__25_, connection_4__12__24_, connection_4__12__23_, 
        connection_4__12__22_, connection_4__12__21_, connection_4__12__20_, 
        connection_4__12__19_, connection_4__12__18_, connection_4__12__17_, 
        connection_4__12__16_, connection_4__12__15_, connection_4__12__14_, 
        connection_4__12__13_, connection_4__12__12_, connection_4__12__11_, 
        connection_4__12__10_, connection_4__12__9_, connection_4__12__8_, 
        connection_4__12__7_, connection_4__12__6_, connection_4__12__5_, 
        connection_4__12__4_, connection_4__12__3_, connection_4__12__2_, 
        connection_4__12__1_, connection_4__12__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[147:146]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_73 first_half_stages_3__group_first_half_3__switch_first_half_1__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__15_, 
        connection_valid_3__13_}), .i_data_bus({connection_3__15__31_, 
        connection_3__15__30_, connection_3__15__29_, connection_3__15__28_, 
        connection_3__15__27_, connection_3__15__26_, connection_3__15__25_, 
        connection_3__15__24_, connection_3__15__23_, connection_3__15__22_, 
        connection_3__15__21_, connection_3__15__20_, connection_3__15__19_, 
        connection_3__15__18_, connection_3__15__17_, connection_3__15__16_, 
        connection_3__15__15_, connection_3__15__14_, connection_3__15__13_, 
        connection_3__15__12_, connection_3__15__11_, connection_3__15__10_, 
        connection_3__15__9_, connection_3__15__8_, connection_3__15__7_, 
        connection_3__15__6_, connection_3__15__5_, connection_3__15__4_, 
        connection_3__15__3_, connection_3__15__2_, connection_3__15__1_, 
        connection_3__15__0_, connection_3__13__31_, connection_3__13__30_, 
        connection_3__13__29_, connection_3__13__28_, connection_3__13__27_, 
        connection_3__13__26_, connection_3__13__25_, connection_3__13__24_, 
        connection_3__13__23_, connection_3__13__22_, connection_3__13__21_, 
        connection_3__13__20_, connection_3__13__19_, connection_3__13__18_, 
        connection_3__13__17_, connection_3__13__16_, connection_3__13__15_, 
        connection_3__13__14_, connection_3__13__13_, connection_3__13__12_, 
        connection_3__13__11_, connection_3__13__10_, connection_3__13__9_, 
        connection_3__13__8_, connection_3__13__7_, connection_3__13__6_, 
        connection_3__13__5_, connection_3__13__4_, connection_3__13__3_, 
        connection_3__13__2_, connection_3__13__1_, connection_3__13__0_}), 
        .o_valid({connection_valid_4__15_, connection_valid_4__14_}), 
        .o_data_bus({connection_4__15__31_, connection_4__15__30_, 
        connection_4__15__29_, connection_4__15__28_, connection_4__15__27_, 
        connection_4__15__26_, connection_4__15__25_, connection_4__15__24_, 
        connection_4__15__23_, connection_4__15__22_, connection_4__15__21_, 
        connection_4__15__20_, connection_4__15__19_, connection_4__15__18_, 
        connection_4__15__17_, connection_4__15__16_, connection_4__15__15_, 
        connection_4__15__14_, connection_4__15__13_, connection_4__15__12_, 
        connection_4__15__11_, connection_4__15__10_, connection_4__15__9_, 
        connection_4__15__8_, connection_4__15__7_, connection_4__15__6_, 
        connection_4__15__5_, connection_4__15__4_, connection_4__15__3_, 
        connection_4__15__2_, connection_4__15__1_, connection_4__15__0_, 
        connection_4__14__31_, connection_4__14__30_, connection_4__14__29_, 
        connection_4__14__28_, connection_4__14__27_, connection_4__14__26_, 
        connection_4__14__25_, connection_4__14__24_, connection_4__14__23_, 
        connection_4__14__22_, connection_4__14__21_, connection_4__14__20_, 
        connection_4__14__19_, connection_4__14__18_, connection_4__14__17_, 
        connection_4__14__16_, connection_4__14__15_, connection_4__14__14_, 
        connection_4__14__13_, connection_4__14__12_, connection_4__14__11_, 
        connection_4__14__10_, connection_4__14__9_, connection_4__14__8_, 
        connection_4__14__7_, connection_4__14__6_, connection_4__14__5_, 
        connection_4__14__4_, connection_4__14__3_, connection_4__14__2_, 
        connection_4__14__1_, connection_4__14__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[145:144]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_72 first_half_stages_3__group_first_half_4__switch_first_half_0__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__18_, 
        connection_valid_3__16_}), .i_data_bus({connection_3__18__31_, 
        connection_3__18__30_, connection_3__18__29_, connection_3__18__28_, 
        connection_3__18__27_, connection_3__18__26_, connection_3__18__25_, 
        connection_3__18__24_, connection_3__18__23_, connection_3__18__22_, 
        connection_3__18__21_, connection_3__18__20_, connection_3__18__19_, 
        connection_3__18__18_, connection_3__18__17_, connection_3__18__16_, 
        connection_3__18__15_, connection_3__18__14_, connection_3__18__13_, 
        connection_3__18__12_, connection_3__18__11_, connection_3__18__10_, 
        connection_3__18__9_, connection_3__18__8_, connection_3__18__7_, 
        connection_3__18__6_, connection_3__18__5_, connection_3__18__4_, 
        connection_3__18__3_, connection_3__18__2_, connection_3__18__1_, 
        connection_3__18__0_, connection_3__16__31_, connection_3__16__30_, 
        connection_3__16__29_, connection_3__16__28_, connection_3__16__27_, 
        connection_3__16__26_, connection_3__16__25_, connection_3__16__24_, 
        connection_3__16__23_, connection_3__16__22_, connection_3__16__21_, 
        connection_3__16__20_, connection_3__16__19_, connection_3__16__18_, 
        connection_3__16__17_, connection_3__16__16_, connection_3__16__15_, 
        connection_3__16__14_, connection_3__16__13_, connection_3__16__12_, 
        connection_3__16__11_, connection_3__16__10_, connection_3__16__9_, 
        connection_3__16__8_, connection_3__16__7_, connection_3__16__6_, 
        connection_3__16__5_, connection_3__16__4_, connection_3__16__3_, 
        connection_3__16__2_, connection_3__16__1_, connection_3__16__0_}), 
        .o_valid({connection_valid_4__17_, connection_valid_4__16_}), 
        .o_data_bus({connection_4__17__31_, connection_4__17__30_, 
        connection_4__17__29_, connection_4__17__28_, connection_4__17__27_, 
        connection_4__17__26_, connection_4__17__25_, connection_4__17__24_, 
        connection_4__17__23_, connection_4__17__22_, connection_4__17__21_, 
        connection_4__17__20_, connection_4__17__19_, connection_4__17__18_, 
        connection_4__17__17_, connection_4__17__16_, connection_4__17__15_, 
        connection_4__17__14_, connection_4__17__13_, connection_4__17__12_, 
        connection_4__17__11_, connection_4__17__10_, connection_4__17__9_, 
        connection_4__17__8_, connection_4__17__7_, connection_4__17__6_, 
        connection_4__17__5_, connection_4__17__4_, connection_4__17__3_, 
        connection_4__17__2_, connection_4__17__1_, connection_4__17__0_, 
        connection_4__16__31_, connection_4__16__30_, connection_4__16__29_, 
        connection_4__16__28_, connection_4__16__27_, connection_4__16__26_, 
        connection_4__16__25_, connection_4__16__24_, connection_4__16__23_, 
        connection_4__16__22_, connection_4__16__21_, connection_4__16__20_, 
        connection_4__16__19_, connection_4__16__18_, connection_4__16__17_, 
        connection_4__16__16_, connection_4__16__15_, connection_4__16__14_, 
        connection_4__16__13_, connection_4__16__12_, connection_4__16__11_, 
        connection_4__16__10_, connection_4__16__9_, connection_4__16__8_, 
        connection_4__16__7_, connection_4__16__6_, connection_4__16__5_, 
        connection_4__16__4_, connection_4__16__3_, connection_4__16__2_, 
        connection_4__16__1_, connection_4__16__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[143:142]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_71 first_half_stages_3__group_first_half_4__switch_first_half_1__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__19_, 
        connection_valid_3__17_}), .i_data_bus({connection_3__19__31_, 
        connection_3__19__30_, connection_3__19__29_, connection_3__19__28_, 
        connection_3__19__27_, connection_3__19__26_, connection_3__19__25_, 
        connection_3__19__24_, connection_3__19__23_, connection_3__19__22_, 
        connection_3__19__21_, connection_3__19__20_, connection_3__19__19_, 
        connection_3__19__18_, connection_3__19__17_, connection_3__19__16_, 
        connection_3__19__15_, connection_3__19__14_, connection_3__19__13_, 
        connection_3__19__12_, connection_3__19__11_, connection_3__19__10_, 
        connection_3__19__9_, connection_3__19__8_, connection_3__19__7_, 
        connection_3__19__6_, connection_3__19__5_, connection_3__19__4_, 
        connection_3__19__3_, connection_3__19__2_, connection_3__19__1_, 
        connection_3__19__0_, connection_3__17__31_, connection_3__17__30_, 
        connection_3__17__29_, connection_3__17__28_, connection_3__17__27_, 
        connection_3__17__26_, connection_3__17__25_, connection_3__17__24_, 
        connection_3__17__23_, connection_3__17__22_, connection_3__17__21_, 
        connection_3__17__20_, connection_3__17__19_, connection_3__17__18_, 
        connection_3__17__17_, connection_3__17__16_, connection_3__17__15_, 
        connection_3__17__14_, connection_3__17__13_, connection_3__17__12_, 
        connection_3__17__11_, connection_3__17__10_, connection_3__17__9_, 
        connection_3__17__8_, connection_3__17__7_, connection_3__17__6_, 
        connection_3__17__5_, connection_3__17__4_, connection_3__17__3_, 
        connection_3__17__2_, connection_3__17__1_, connection_3__17__0_}), 
        .o_valid({connection_valid_4__19_, connection_valid_4__18_}), 
        .o_data_bus({connection_4__19__31_, connection_4__19__30_, 
        connection_4__19__29_, connection_4__19__28_, connection_4__19__27_, 
        connection_4__19__26_, connection_4__19__25_, connection_4__19__24_, 
        connection_4__19__23_, connection_4__19__22_, connection_4__19__21_, 
        connection_4__19__20_, connection_4__19__19_, connection_4__19__18_, 
        connection_4__19__17_, connection_4__19__16_, connection_4__19__15_, 
        connection_4__19__14_, connection_4__19__13_, connection_4__19__12_, 
        connection_4__19__11_, connection_4__19__10_, connection_4__19__9_, 
        connection_4__19__8_, connection_4__19__7_, connection_4__19__6_, 
        connection_4__19__5_, connection_4__19__4_, connection_4__19__3_, 
        connection_4__19__2_, connection_4__19__1_, connection_4__19__0_, 
        connection_4__18__31_, connection_4__18__30_, connection_4__18__29_, 
        connection_4__18__28_, connection_4__18__27_, connection_4__18__26_, 
        connection_4__18__25_, connection_4__18__24_, connection_4__18__23_, 
        connection_4__18__22_, connection_4__18__21_, connection_4__18__20_, 
        connection_4__18__19_, connection_4__18__18_, connection_4__18__17_, 
        connection_4__18__16_, connection_4__18__15_, connection_4__18__14_, 
        connection_4__18__13_, connection_4__18__12_, connection_4__18__11_, 
        connection_4__18__10_, connection_4__18__9_, connection_4__18__8_, 
        connection_4__18__7_, connection_4__18__6_, connection_4__18__5_, 
        connection_4__18__4_, connection_4__18__3_, connection_4__18__2_, 
        connection_4__18__1_, connection_4__18__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[141:140]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_70 first_half_stages_3__group_first_half_5__switch_first_half_0__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__22_, 
        connection_valid_3__20_}), .i_data_bus({connection_3__22__31_, 
        connection_3__22__30_, connection_3__22__29_, connection_3__22__28_, 
        connection_3__22__27_, connection_3__22__26_, connection_3__22__25_, 
        connection_3__22__24_, connection_3__22__23_, connection_3__22__22_, 
        connection_3__22__21_, connection_3__22__20_, connection_3__22__19_, 
        connection_3__22__18_, connection_3__22__17_, connection_3__22__16_, 
        connection_3__22__15_, connection_3__22__14_, connection_3__22__13_, 
        connection_3__22__12_, connection_3__22__11_, connection_3__22__10_, 
        connection_3__22__9_, connection_3__22__8_, connection_3__22__7_, 
        connection_3__22__6_, connection_3__22__5_, connection_3__22__4_, 
        connection_3__22__3_, connection_3__22__2_, connection_3__22__1_, 
        connection_3__22__0_, connection_3__20__31_, connection_3__20__30_, 
        connection_3__20__29_, connection_3__20__28_, connection_3__20__27_, 
        connection_3__20__26_, connection_3__20__25_, connection_3__20__24_, 
        connection_3__20__23_, connection_3__20__22_, connection_3__20__21_, 
        connection_3__20__20_, connection_3__20__19_, connection_3__20__18_, 
        connection_3__20__17_, connection_3__20__16_, connection_3__20__15_, 
        connection_3__20__14_, connection_3__20__13_, connection_3__20__12_, 
        connection_3__20__11_, connection_3__20__10_, connection_3__20__9_, 
        connection_3__20__8_, connection_3__20__7_, connection_3__20__6_, 
        connection_3__20__5_, connection_3__20__4_, connection_3__20__3_, 
        connection_3__20__2_, connection_3__20__1_, connection_3__20__0_}), 
        .o_valid({connection_valid_4__21_, connection_valid_4__20_}), 
        .o_data_bus({connection_4__21__31_, connection_4__21__30_, 
        connection_4__21__29_, connection_4__21__28_, connection_4__21__27_, 
        connection_4__21__26_, connection_4__21__25_, connection_4__21__24_, 
        connection_4__21__23_, connection_4__21__22_, connection_4__21__21_, 
        connection_4__21__20_, connection_4__21__19_, connection_4__21__18_, 
        connection_4__21__17_, connection_4__21__16_, connection_4__21__15_, 
        connection_4__21__14_, connection_4__21__13_, connection_4__21__12_, 
        connection_4__21__11_, connection_4__21__10_, connection_4__21__9_, 
        connection_4__21__8_, connection_4__21__7_, connection_4__21__6_, 
        connection_4__21__5_, connection_4__21__4_, connection_4__21__3_, 
        connection_4__21__2_, connection_4__21__1_, connection_4__21__0_, 
        connection_4__20__31_, connection_4__20__30_, connection_4__20__29_, 
        connection_4__20__28_, connection_4__20__27_, connection_4__20__26_, 
        connection_4__20__25_, connection_4__20__24_, connection_4__20__23_, 
        connection_4__20__22_, connection_4__20__21_, connection_4__20__20_, 
        connection_4__20__19_, connection_4__20__18_, connection_4__20__17_, 
        connection_4__20__16_, connection_4__20__15_, connection_4__20__14_, 
        connection_4__20__13_, connection_4__20__12_, connection_4__20__11_, 
        connection_4__20__10_, connection_4__20__9_, connection_4__20__8_, 
        connection_4__20__7_, connection_4__20__6_, connection_4__20__5_, 
        connection_4__20__4_, connection_4__20__3_, connection_4__20__2_, 
        connection_4__20__1_, connection_4__20__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[139:138]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_69 first_half_stages_3__group_first_half_5__switch_first_half_1__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__23_, 
        connection_valid_3__21_}), .i_data_bus({connection_3__23__31_, 
        connection_3__23__30_, connection_3__23__29_, connection_3__23__28_, 
        connection_3__23__27_, connection_3__23__26_, connection_3__23__25_, 
        connection_3__23__24_, connection_3__23__23_, connection_3__23__22_, 
        connection_3__23__21_, connection_3__23__20_, connection_3__23__19_, 
        connection_3__23__18_, connection_3__23__17_, connection_3__23__16_, 
        connection_3__23__15_, connection_3__23__14_, connection_3__23__13_, 
        connection_3__23__12_, connection_3__23__11_, connection_3__23__10_, 
        connection_3__23__9_, connection_3__23__8_, connection_3__23__7_, 
        connection_3__23__6_, connection_3__23__5_, connection_3__23__4_, 
        connection_3__23__3_, connection_3__23__2_, connection_3__23__1_, 
        connection_3__23__0_, connection_3__21__31_, connection_3__21__30_, 
        connection_3__21__29_, connection_3__21__28_, connection_3__21__27_, 
        connection_3__21__26_, connection_3__21__25_, connection_3__21__24_, 
        connection_3__21__23_, connection_3__21__22_, connection_3__21__21_, 
        connection_3__21__20_, connection_3__21__19_, connection_3__21__18_, 
        connection_3__21__17_, connection_3__21__16_, connection_3__21__15_, 
        connection_3__21__14_, connection_3__21__13_, connection_3__21__12_, 
        connection_3__21__11_, connection_3__21__10_, connection_3__21__9_, 
        connection_3__21__8_, connection_3__21__7_, connection_3__21__6_, 
        connection_3__21__5_, connection_3__21__4_, connection_3__21__3_, 
        connection_3__21__2_, connection_3__21__1_, connection_3__21__0_}), 
        .o_valid({connection_valid_4__23_, connection_valid_4__22_}), 
        .o_data_bus({connection_4__23__31_, connection_4__23__30_, 
        connection_4__23__29_, connection_4__23__28_, connection_4__23__27_, 
        connection_4__23__26_, connection_4__23__25_, connection_4__23__24_, 
        connection_4__23__23_, connection_4__23__22_, connection_4__23__21_, 
        connection_4__23__20_, connection_4__23__19_, connection_4__23__18_, 
        connection_4__23__17_, connection_4__23__16_, connection_4__23__15_, 
        connection_4__23__14_, connection_4__23__13_, connection_4__23__12_, 
        connection_4__23__11_, connection_4__23__10_, connection_4__23__9_, 
        connection_4__23__8_, connection_4__23__7_, connection_4__23__6_, 
        connection_4__23__5_, connection_4__23__4_, connection_4__23__3_, 
        connection_4__23__2_, connection_4__23__1_, connection_4__23__0_, 
        connection_4__22__31_, connection_4__22__30_, connection_4__22__29_, 
        connection_4__22__28_, connection_4__22__27_, connection_4__22__26_, 
        connection_4__22__25_, connection_4__22__24_, connection_4__22__23_, 
        connection_4__22__22_, connection_4__22__21_, connection_4__22__20_, 
        connection_4__22__19_, connection_4__22__18_, connection_4__22__17_, 
        connection_4__22__16_, connection_4__22__15_, connection_4__22__14_, 
        connection_4__22__13_, connection_4__22__12_, connection_4__22__11_, 
        connection_4__22__10_, connection_4__22__9_, connection_4__22__8_, 
        connection_4__22__7_, connection_4__22__6_, connection_4__22__5_, 
        connection_4__22__4_, connection_4__22__3_, connection_4__22__2_, 
        connection_4__22__1_, connection_4__22__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[137:136]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_68 first_half_stages_3__group_first_half_6__switch_first_half_0__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__26_, 
        connection_valid_3__24_}), .i_data_bus({connection_3__26__31_, 
        connection_3__26__30_, connection_3__26__29_, connection_3__26__28_, 
        connection_3__26__27_, connection_3__26__26_, connection_3__26__25_, 
        connection_3__26__24_, connection_3__26__23_, connection_3__26__22_, 
        connection_3__26__21_, connection_3__26__20_, connection_3__26__19_, 
        connection_3__26__18_, connection_3__26__17_, connection_3__26__16_, 
        connection_3__26__15_, connection_3__26__14_, connection_3__26__13_, 
        connection_3__26__12_, connection_3__26__11_, connection_3__26__10_, 
        connection_3__26__9_, connection_3__26__8_, connection_3__26__7_, 
        connection_3__26__6_, connection_3__26__5_, connection_3__26__4_, 
        connection_3__26__3_, connection_3__26__2_, connection_3__26__1_, 
        connection_3__26__0_, connection_3__24__31_, connection_3__24__30_, 
        connection_3__24__29_, connection_3__24__28_, connection_3__24__27_, 
        connection_3__24__26_, connection_3__24__25_, connection_3__24__24_, 
        connection_3__24__23_, connection_3__24__22_, connection_3__24__21_, 
        connection_3__24__20_, connection_3__24__19_, connection_3__24__18_, 
        connection_3__24__17_, connection_3__24__16_, connection_3__24__15_, 
        connection_3__24__14_, connection_3__24__13_, connection_3__24__12_, 
        connection_3__24__11_, connection_3__24__10_, connection_3__24__9_, 
        connection_3__24__8_, connection_3__24__7_, connection_3__24__6_, 
        connection_3__24__5_, connection_3__24__4_, connection_3__24__3_, 
        connection_3__24__2_, connection_3__24__1_, connection_3__24__0_}), 
        .o_valid({connection_valid_4__25_, connection_valid_4__24_}), 
        .o_data_bus({connection_4__25__31_, connection_4__25__30_, 
        connection_4__25__29_, connection_4__25__28_, connection_4__25__27_, 
        connection_4__25__26_, connection_4__25__25_, connection_4__25__24_, 
        connection_4__25__23_, connection_4__25__22_, connection_4__25__21_, 
        connection_4__25__20_, connection_4__25__19_, connection_4__25__18_, 
        connection_4__25__17_, connection_4__25__16_, connection_4__25__15_, 
        connection_4__25__14_, connection_4__25__13_, connection_4__25__12_, 
        connection_4__25__11_, connection_4__25__10_, connection_4__25__9_, 
        connection_4__25__8_, connection_4__25__7_, connection_4__25__6_, 
        connection_4__25__5_, connection_4__25__4_, connection_4__25__3_, 
        connection_4__25__2_, connection_4__25__1_, connection_4__25__0_, 
        connection_4__24__31_, connection_4__24__30_, connection_4__24__29_, 
        connection_4__24__28_, connection_4__24__27_, connection_4__24__26_, 
        connection_4__24__25_, connection_4__24__24_, connection_4__24__23_, 
        connection_4__24__22_, connection_4__24__21_, connection_4__24__20_, 
        connection_4__24__19_, connection_4__24__18_, connection_4__24__17_, 
        connection_4__24__16_, connection_4__24__15_, connection_4__24__14_, 
        connection_4__24__13_, connection_4__24__12_, connection_4__24__11_, 
        connection_4__24__10_, connection_4__24__9_, connection_4__24__8_, 
        connection_4__24__7_, connection_4__24__6_, connection_4__24__5_, 
        connection_4__24__4_, connection_4__24__3_, connection_4__24__2_, 
        connection_4__24__1_, connection_4__24__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[135:134]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_67 first_half_stages_3__group_first_half_6__switch_first_half_1__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__27_, 
        connection_valid_3__25_}), .i_data_bus({connection_3__27__31_, 
        connection_3__27__30_, connection_3__27__29_, connection_3__27__28_, 
        connection_3__27__27_, connection_3__27__26_, connection_3__27__25_, 
        connection_3__27__24_, connection_3__27__23_, connection_3__27__22_, 
        connection_3__27__21_, connection_3__27__20_, connection_3__27__19_, 
        connection_3__27__18_, connection_3__27__17_, connection_3__27__16_, 
        connection_3__27__15_, connection_3__27__14_, connection_3__27__13_, 
        connection_3__27__12_, connection_3__27__11_, connection_3__27__10_, 
        connection_3__27__9_, connection_3__27__8_, connection_3__27__7_, 
        connection_3__27__6_, connection_3__27__5_, connection_3__27__4_, 
        connection_3__27__3_, connection_3__27__2_, connection_3__27__1_, 
        connection_3__27__0_, connection_3__25__31_, connection_3__25__30_, 
        connection_3__25__29_, connection_3__25__28_, connection_3__25__27_, 
        connection_3__25__26_, connection_3__25__25_, connection_3__25__24_, 
        connection_3__25__23_, connection_3__25__22_, connection_3__25__21_, 
        connection_3__25__20_, connection_3__25__19_, connection_3__25__18_, 
        connection_3__25__17_, connection_3__25__16_, connection_3__25__15_, 
        connection_3__25__14_, connection_3__25__13_, connection_3__25__12_, 
        connection_3__25__11_, connection_3__25__10_, connection_3__25__9_, 
        connection_3__25__8_, connection_3__25__7_, connection_3__25__6_, 
        connection_3__25__5_, connection_3__25__4_, connection_3__25__3_, 
        connection_3__25__2_, connection_3__25__1_, connection_3__25__0_}), 
        .o_valid({connection_valid_4__27_, connection_valid_4__26_}), 
        .o_data_bus({connection_4__27__31_, connection_4__27__30_, 
        connection_4__27__29_, connection_4__27__28_, connection_4__27__27_, 
        connection_4__27__26_, connection_4__27__25_, connection_4__27__24_, 
        connection_4__27__23_, connection_4__27__22_, connection_4__27__21_, 
        connection_4__27__20_, connection_4__27__19_, connection_4__27__18_, 
        connection_4__27__17_, connection_4__27__16_, connection_4__27__15_, 
        connection_4__27__14_, connection_4__27__13_, connection_4__27__12_, 
        connection_4__27__11_, connection_4__27__10_, connection_4__27__9_, 
        connection_4__27__8_, connection_4__27__7_, connection_4__27__6_, 
        connection_4__27__5_, connection_4__27__4_, connection_4__27__3_, 
        connection_4__27__2_, connection_4__27__1_, connection_4__27__0_, 
        connection_4__26__31_, connection_4__26__30_, connection_4__26__29_, 
        connection_4__26__28_, connection_4__26__27_, connection_4__26__26_, 
        connection_4__26__25_, connection_4__26__24_, connection_4__26__23_, 
        connection_4__26__22_, connection_4__26__21_, connection_4__26__20_, 
        connection_4__26__19_, connection_4__26__18_, connection_4__26__17_, 
        connection_4__26__16_, connection_4__26__15_, connection_4__26__14_, 
        connection_4__26__13_, connection_4__26__12_, connection_4__26__11_, 
        connection_4__26__10_, connection_4__26__9_, connection_4__26__8_, 
        connection_4__26__7_, connection_4__26__6_, connection_4__26__5_, 
        connection_4__26__4_, connection_4__26__3_, connection_4__26__2_, 
        connection_4__26__1_, connection_4__26__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[133:132]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_66 first_half_stages_3__group_first_half_7__switch_first_half_0__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__30_, 
        connection_valid_3__28_}), .i_data_bus({connection_3__30__31_, 
        connection_3__30__30_, connection_3__30__29_, connection_3__30__28_, 
        connection_3__30__27_, connection_3__30__26_, connection_3__30__25_, 
        connection_3__30__24_, connection_3__30__23_, connection_3__30__22_, 
        connection_3__30__21_, connection_3__30__20_, connection_3__30__19_, 
        connection_3__30__18_, connection_3__30__17_, connection_3__30__16_, 
        connection_3__30__15_, connection_3__30__14_, connection_3__30__13_, 
        connection_3__30__12_, connection_3__30__11_, connection_3__30__10_, 
        connection_3__30__9_, connection_3__30__8_, connection_3__30__7_, 
        connection_3__30__6_, connection_3__30__5_, connection_3__30__4_, 
        connection_3__30__3_, connection_3__30__2_, connection_3__30__1_, 
        connection_3__30__0_, connection_3__28__31_, connection_3__28__30_, 
        connection_3__28__29_, connection_3__28__28_, connection_3__28__27_, 
        connection_3__28__26_, connection_3__28__25_, connection_3__28__24_, 
        connection_3__28__23_, connection_3__28__22_, connection_3__28__21_, 
        connection_3__28__20_, connection_3__28__19_, connection_3__28__18_, 
        connection_3__28__17_, connection_3__28__16_, connection_3__28__15_, 
        connection_3__28__14_, connection_3__28__13_, connection_3__28__12_, 
        connection_3__28__11_, connection_3__28__10_, connection_3__28__9_, 
        connection_3__28__8_, connection_3__28__7_, connection_3__28__6_, 
        connection_3__28__5_, connection_3__28__4_, connection_3__28__3_, 
        connection_3__28__2_, connection_3__28__1_, connection_3__28__0_}), 
        .o_valid({connection_valid_4__29_, connection_valid_4__28_}), 
        .o_data_bus({connection_4__29__31_, connection_4__29__30_, 
        connection_4__29__29_, connection_4__29__28_, connection_4__29__27_, 
        connection_4__29__26_, connection_4__29__25_, connection_4__29__24_, 
        connection_4__29__23_, connection_4__29__22_, connection_4__29__21_, 
        connection_4__29__20_, connection_4__29__19_, connection_4__29__18_, 
        connection_4__29__17_, connection_4__29__16_, connection_4__29__15_, 
        connection_4__29__14_, connection_4__29__13_, connection_4__29__12_, 
        connection_4__29__11_, connection_4__29__10_, connection_4__29__9_, 
        connection_4__29__8_, connection_4__29__7_, connection_4__29__6_, 
        connection_4__29__5_, connection_4__29__4_, connection_4__29__3_, 
        connection_4__29__2_, connection_4__29__1_, connection_4__29__0_, 
        connection_4__28__31_, connection_4__28__30_, connection_4__28__29_, 
        connection_4__28__28_, connection_4__28__27_, connection_4__28__26_, 
        connection_4__28__25_, connection_4__28__24_, connection_4__28__23_, 
        connection_4__28__22_, connection_4__28__21_, connection_4__28__20_, 
        connection_4__28__19_, connection_4__28__18_, connection_4__28__17_, 
        connection_4__28__16_, connection_4__28__15_, connection_4__28__14_, 
        connection_4__28__13_, connection_4__28__12_, connection_4__28__11_, 
        connection_4__28__10_, connection_4__28__9_, connection_4__28__8_, 
        connection_4__28__7_, connection_4__28__6_, connection_4__28__5_, 
        connection_4__28__4_, connection_4__28__3_, connection_4__28__2_, 
        connection_4__28__1_, connection_4__28__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[131:130]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_65 first_half_stages_3__group_first_half_7__switch_first_half_1__second_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__31_, 
        connection_valid_3__29_}), .i_data_bus({connection_3__31__31_, 
        connection_3__31__30_, connection_3__31__29_, connection_3__31__28_, 
        connection_3__31__27_, connection_3__31__26_, connection_3__31__25_, 
        connection_3__31__24_, connection_3__31__23_, connection_3__31__22_, 
        connection_3__31__21_, connection_3__31__20_, connection_3__31__19_, 
        connection_3__31__18_, connection_3__31__17_, connection_3__31__16_, 
        connection_3__31__15_, connection_3__31__14_, connection_3__31__13_, 
        connection_3__31__12_, connection_3__31__11_, connection_3__31__10_, 
        connection_3__31__9_, connection_3__31__8_, connection_3__31__7_, 
        connection_3__31__6_, connection_3__31__5_, connection_3__31__4_, 
        connection_3__31__3_, connection_3__31__2_, connection_3__31__1_, 
        connection_3__31__0_, connection_3__29__31_, connection_3__29__30_, 
        connection_3__29__29_, connection_3__29__28_, connection_3__29__27_, 
        connection_3__29__26_, connection_3__29__25_, connection_3__29__24_, 
        connection_3__29__23_, connection_3__29__22_, connection_3__29__21_, 
        connection_3__29__20_, connection_3__29__19_, connection_3__29__18_, 
        connection_3__29__17_, connection_3__29__16_, connection_3__29__15_, 
        connection_3__29__14_, connection_3__29__13_, connection_3__29__12_, 
        connection_3__29__11_, connection_3__29__10_, connection_3__29__9_, 
        connection_3__29__8_, connection_3__29__7_, connection_3__29__6_, 
        connection_3__29__5_, connection_3__29__4_, connection_3__29__3_, 
        connection_3__29__2_, connection_3__29__1_, connection_3__29__0_}), 
        .o_valid({connection_valid_4__31_, connection_valid_4__30_}), 
        .o_data_bus({connection_4__31__31_, connection_4__31__30_, 
        connection_4__31__29_, connection_4__31__28_, connection_4__31__27_, 
        connection_4__31__26_, connection_4__31__25_, connection_4__31__24_, 
        connection_4__31__23_, connection_4__31__22_, connection_4__31__21_, 
        connection_4__31__20_, connection_4__31__19_, connection_4__31__18_, 
        connection_4__31__17_, connection_4__31__16_, connection_4__31__15_, 
        connection_4__31__14_, connection_4__31__13_, connection_4__31__12_, 
        connection_4__31__11_, connection_4__31__10_, connection_4__31__9_, 
        connection_4__31__8_, connection_4__31__7_, connection_4__31__6_, 
        connection_4__31__5_, connection_4__31__4_, connection_4__31__3_, 
        connection_4__31__2_, connection_4__31__1_, connection_4__31__0_, 
        connection_4__30__31_, connection_4__30__30_, connection_4__30__29_, 
        connection_4__30__28_, connection_4__30__27_, connection_4__30__26_, 
        connection_4__30__25_, connection_4__30__24_, connection_4__30__23_, 
        connection_4__30__22_, connection_4__30__21_, connection_4__30__20_, 
        connection_4__30__19_, connection_4__30__18_, connection_4__30__17_, 
        connection_4__30__16_, connection_4__30__15_, connection_4__30__14_, 
        connection_4__30__13_, connection_4__30__12_, connection_4__30__11_, 
        connection_4__30__10_, connection_4__30__9_, connection_4__30__8_, 
        connection_4__30__7_, connection_4__30__6_, connection_4__30__5_, 
        connection_4__30__4_, connection_4__30__3_, connection_4__30__2_, 
        connection_4__30__1_, connection_4__30__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[129:128]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_64 second_half_stages_4__group_sec_half_0__switch_sec_half_0__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__2_, 
        connection_valid_4__0_}), .i_data_bus({connection_4__2__31_, 
        connection_4__2__30_, connection_4__2__29_, connection_4__2__28_, 
        connection_4__2__27_, connection_4__2__26_, connection_4__2__25_, 
        connection_4__2__24_, connection_4__2__23_, connection_4__2__22_, 
        connection_4__2__21_, connection_4__2__20_, connection_4__2__19_, 
        connection_4__2__18_, connection_4__2__17_, connection_4__2__16_, 
        connection_4__2__15_, connection_4__2__14_, connection_4__2__13_, 
        connection_4__2__12_, connection_4__2__11_, connection_4__2__10_, 
        connection_4__2__9_, connection_4__2__8_, connection_4__2__7_, 
        connection_4__2__6_, connection_4__2__5_, connection_4__2__4_, 
        connection_4__2__3_, connection_4__2__2_, connection_4__2__1_, 
        connection_4__2__0_, connection_4__0__31_, connection_4__0__30_, 
        connection_4__0__29_, connection_4__0__28_, connection_4__0__27_, 
        connection_4__0__26_, connection_4__0__25_, connection_4__0__24_, 
        connection_4__0__23_, connection_4__0__22_, connection_4__0__21_, 
        connection_4__0__20_, connection_4__0__19_, connection_4__0__18_, 
        connection_4__0__17_, connection_4__0__16_, connection_4__0__15_, 
        connection_4__0__14_, connection_4__0__13_, connection_4__0__12_, 
        connection_4__0__11_, connection_4__0__10_, connection_4__0__9_, 
        connection_4__0__8_, connection_4__0__7_, connection_4__0__6_, 
        connection_4__0__5_, connection_4__0__4_, connection_4__0__3_, 
        connection_4__0__2_, connection_4__0__1_, connection_4__0__0_}), 
        .o_valid({connection_valid_5__1_, connection_valid_5__0_}), 
        .o_data_bus({connection_5__1__31_, connection_5__1__30_, 
        connection_5__1__29_, connection_5__1__28_, connection_5__1__27_, 
        connection_5__1__26_, connection_5__1__25_, connection_5__1__24_, 
        connection_5__1__23_, connection_5__1__22_, connection_5__1__21_, 
        connection_5__1__20_, connection_5__1__19_, connection_5__1__18_, 
        connection_5__1__17_, connection_5__1__16_, connection_5__1__15_, 
        connection_5__1__14_, connection_5__1__13_, connection_5__1__12_, 
        connection_5__1__11_, connection_5__1__10_, connection_5__1__9_, 
        connection_5__1__8_, connection_5__1__7_, connection_5__1__6_, 
        connection_5__1__5_, connection_5__1__4_, connection_5__1__3_, 
        connection_5__1__2_, connection_5__1__1_, connection_5__1__0_, 
        connection_5__0__31_, connection_5__0__30_, connection_5__0__29_, 
        connection_5__0__28_, connection_5__0__27_, connection_5__0__26_, 
        connection_5__0__25_, connection_5__0__24_, connection_5__0__23_, 
        connection_5__0__22_, connection_5__0__21_, connection_5__0__20_, 
        connection_5__0__19_, connection_5__0__18_, connection_5__0__17_, 
        connection_5__0__16_, connection_5__0__15_, connection_5__0__14_, 
        connection_5__0__13_, connection_5__0__12_, connection_5__0__11_, 
        connection_5__0__10_, connection_5__0__9_, connection_5__0__8_, 
        connection_5__0__7_, connection_5__0__6_, connection_5__0__5_, 
        connection_5__0__4_, connection_5__0__3_, connection_5__0__2_, 
        connection_5__0__1_, connection_5__0__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[127:126]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_63 second_half_stages_4__group_sec_half_0__switch_sec_half_1__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__3_, 
        connection_valid_4__1_}), .i_data_bus({connection_4__3__31_, 
        connection_4__3__30_, connection_4__3__29_, connection_4__3__28_, 
        connection_4__3__27_, connection_4__3__26_, connection_4__3__25_, 
        connection_4__3__24_, connection_4__3__23_, connection_4__3__22_, 
        connection_4__3__21_, connection_4__3__20_, connection_4__3__19_, 
        connection_4__3__18_, connection_4__3__17_, connection_4__3__16_, 
        connection_4__3__15_, connection_4__3__14_, connection_4__3__13_, 
        connection_4__3__12_, connection_4__3__11_, connection_4__3__10_, 
        connection_4__3__9_, connection_4__3__8_, connection_4__3__7_, 
        connection_4__3__6_, connection_4__3__5_, connection_4__3__4_, 
        connection_4__3__3_, connection_4__3__2_, connection_4__3__1_, 
        connection_4__3__0_, connection_4__1__31_, connection_4__1__30_, 
        connection_4__1__29_, connection_4__1__28_, connection_4__1__27_, 
        connection_4__1__26_, connection_4__1__25_, connection_4__1__24_, 
        connection_4__1__23_, connection_4__1__22_, connection_4__1__21_, 
        connection_4__1__20_, connection_4__1__19_, connection_4__1__18_, 
        connection_4__1__17_, connection_4__1__16_, connection_4__1__15_, 
        connection_4__1__14_, connection_4__1__13_, connection_4__1__12_, 
        connection_4__1__11_, connection_4__1__10_, connection_4__1__9_, 
        connection_4__1__8_, connection_4__1__7_, connection_4__1__6_, 
        connection_4__1__5_, connection_4__1__4_, connection_4__1__3_, 
        connection_4__1__2_, connection_4__1__1_, connection_4__1__0_}), 
        .o_valid({connection_valid_5__3_, connection_valid_5__2_}), 
        .o_data_bus({connection_5__3__31_, connection_5__3__30_, 
        connection_5__3__29_, connection_5__3__28_, connection_5__3__27_, 
        connection_5__3__26_, connection_5__3__25_, connection_5__3__24_, 
        connection_5__3__23_, connection_5__3__22_, connection_5__3__21_, 
        connection_5__3__20_, connection_5__3__19_, connection_5__3__18_, 
        connection_5__3__17_, connection_5__3__16_, connection_5__3__15_, 
        connection_5__3__14_, connection_5__3__13_, connection_5__3__12_, 
        connection_5__3__11_, connection_5__3__10_, connection_5__3__9_, 
        connection_5__3__8_, connection_5__3__7_, connection_5__3__6_, 
        connection_5__3__5_, connection_5__3__4_, connection_5__3__3_, 
        connection_5__3__2_, connection_5__3__1_, connection_5__3__0_, 
        connection_5__2__31_, connection_5__2__30_, connection_5__2__29_, 
        connection_5__2__28_, connection_5__2__27_, connection_5__2__26_, 
        connection_5__2__25_, connection_5__2__24_, connection_5__2__23_, 
        connection_5__2__22_, connection_5__2__21_, connection_5__2__20_, 
        connection_5__2__19_, connection_5__2__18_, connection_5__2__17_, 
        connection_5__2__16_, connection_5__2__15_, connection_5__2__14_, 
        connection_5__2__13_, connection_5__2__12_, connection_5__2__11_, 
        connection_5__2__10_, connection_5__2__9_, connection_5__2__8_, 
        connection_5__2__7_, connection_5__2__6_, connection_5__2__5_, 
        connection_5__2__4_, connection_5__2__3_, connection_5__2__2_, 
        connection_5__2__1_, connection_5__2__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[125:124]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_62 second_half_stages_4__group_sec_half_1__switch_sec_half_0__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__6_, 
        connection_valid_4__4_}), .i_data_bus({connection_4__6__31_, 
        connection_4__6__30_, connection_4__6__29_, connection_4__6__28_, 
        connection_4__6__27_, connection_4__6__26_, connection_4__6__25_, 
        connection_4__6__24_, connection_4__6__23_, connection_4__6__22_, 
        connection_4__6__21_, connection_4__6__20_, connection_4__6__19_, 
        connection_4__6__18_, connection_4__6__17_, connection_4__6__16_, 
        connection_4__6__15_, connection_4__6__14_, connection_4__6__13_, 
        connection_4__6__12_, connection_4__6__11_, connection_4__6__10_, 
        connection_4__6__9_, connection_4__6__8_, connection_4__6__7_, 
        connection_4__6__6_, connection_4__6__5_, connection_4__6__4_, 
        connection_4__6__3_, connection_4__6__2_, connection_4__6__1_, 
        connection_4__6__0_, connection_4__4__31_, connection_4__4__30_, 
        connection_4__4__29_, connection_4__4__28_, connection_4__4__27_, 
        connection_4__4__26_, connection_4__4__25_, connection_4__4__24_, 
        connection_4__4__23_, connection_4__4__22_, connection_4__4__21_, 
        connection_4__4__20_, connection_4__4__19_, connection_4__4__18_, 
        connection_4__4__17_, connection_4__4__16_, connection_4__4__15_, 
        connection_4__4__14_, connection_4__4__13_, connection_4__4__12_, 
        connection_4__4__11_, connection_4__4__10_, connection_4__4__9_, 
        connection_4__4__8_, connection_4__4__7_, connection_4__4__6_, 
        connection_4__4__5_, connection_4__4__4_, connection_4__4__3_, 
        connection_4__4__2_, connection_4__4__1_, connection_4__4__0_}), 
        .o_valid({connection_valid_5__5_, connection_valid_5__4_}), 
        .o_data_bus({connection_5__5__31_, connection_5__5__30_, 
        connection_5__5__29_, connection_5__5__28_, connection_5__5__27_, 
        connection_5__5__26_, connection_5__5__25_, connection_5__5__24_, 
        connection_5__5__23_, connection_5__5__22_, connection_5__5__21_, 
        connection_5__5__20_, connection_5__5__19_, connection_5__5__18_, 
        connection_5__5__17_, connection_5__5__16_, connection_5__5__15_, 
        connection_5__5__14_, connection_5__5__13_, connection_5__5__12_, 
        connection_5__5__11_, connection_5__5__10_, connection_5__5__9_, 
        connection_5__5__8_, connection_5__5__7_, connection_5__5__6_, 
        connection_5__5__5_, connection_5__5__4_, connection_5__5__3_, 
        connection_5__5__2_, connection_5__5__1_, connection_5__5__0_, 
        connection_5__4__31_, connection_5__4__30_, connection_5__4__29_, 
        connection_5__4__28_, connection_5__4__27_, connection_5__4__26_, 
        connection_5__4__25_, connection_5__4__24_, connection_5__4__23_, 
        connection_5__4__22_, connection_5__4__21_, connection_5__4__20_, 
        connection_5__4__19_, connection_5__4__18_, connection_5__4__17_, 
        connection_5__4__16_, connection_5__4__15_, connection_5__4__14_, 
        connection_5__4__13_, connection_5__4__12_, connection_5__4__11_, 
        connection_5__4__10_, connection_5__4__9_, connection_5__4__8_, 
        connection_5__4__7_, connection_5__4__6_, connection_5__4__5_, 
        connection_5__4__4_, connection_5__4__3_, connection_5__4__2_, 
        connection_5__4__1_, connection_5__4__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[123:122]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_61 second_half_stages_4__group_sec_half_1__switch_sec_half_1__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__7_, 
        connection_valid_4__5_}), .i_data_bus({connection_4__7__31_, 
        connection_4__7__30_, connection_4__7__29_, connection_4__7__28_, 
        connection_4__7__27_, connection_4__7__26_, connection_4__7__25_, 
        connection_4__7__24_, connection_4__7__23_, connection_4__7__22_, 
        connection_4__7__21_, connection_4__7__20_, connection_4__7__19_, 
        connection_4__7__18_, connection_4__7__17_, connection_4__7__16_, 
        connection_4__7__15_, connection_4__7__14_, connection_4__7__13_, 
        connection_4__7__12_, connection_4__7__11_, connection_4__7__10_, 
        connection_4__7__9_, connection_4__7__8_, connection_4__7__7_, 
        connection_4__7__6_, connection_4__7__5_, connection_4__7__4_, 
        connection_4__7__3_, connection_4__7__2_, connection_4__7__1_, 
        connection_4__7__0_, connection_4__5__31_, connection_4__5__30_, 
        connection_4__5__29_, connection_4__5__28_, connection_4__5__27_, 
        connection_4__5__26_, connection_4__5__25_, connection_4__5__24_, 
        connection_4__5__23_, connection_4__5__22_, connection_4__5__21_, 
        connection_4__5__20_, connection_4__5__19_, connection_4__5__18_, 
        connection_4__5__17_, connection_4__5__16_, connection_4__5__15_, 
        connection_4__5__14_, connection_4__5__13_, connection_4__5__12_, 
        connection_4__5__11_, connection_4__5__10_, connection_4__5__9_, 
        connection_4__5__8_, connection_4__5__7_, connection_4__5__6_, 
        connection_4__5__5_, connection_4__5__4_, connection_4__5__3_, 
        connection_4__5__2_, connection_4__5__1_, connection_4__5__0_}), 
        .o_valid({connection_valid_5__7_, connection_valid_5__6_}), 
        .o_data_bus({connection_5__7__31_, connection_5__7__30_, 
        connection_5__7__29_, connection_5__7__28_, connection_5__7__27_, 
        connection_5__7__26_, connection_5__7__25_, connection_5__7__24_, 
        connection_5__7__23_, connection_5__7__22_, connection_5__7__21_, 
        connection_5__7__20_, connection_5__7__19_, connection_5__7__18_, 
        connection_5__7__17_, connection_5__7__16_, connection_5__7__15_, 
        connection_5__7__14_, connection_5__7__13_, connection_5__7__12_, 
        connection_5__7__11_, connection_5__7__10_, connection_5__7__9_, 
        connection_5__7__8_, connection_5__7__7_, connection_5__7__6_, 
        connection_5__7__5_, connection_5__7__4_, connection_5__7__3_, 
        connection_5__7__2_, connection_5__7__1_, connection_5__7__0_, 
        connection_5__6__31_, connection_5__6__30_, connection_5__6__29_, 
        connection_5__6__28_, connection_5__6__27_, connection_5__6__26_, 
        connection_5__6__25_, connection_5__6__24_, connection_5__6__23_, 
        connection_5__6__22_, connection_5__6__21_, connection_5__6__20_, 
        connection_5__6__19_, connection_5__6__18_, connection_5__6__17_, 
        connection_5__6__16_, connection_5__6__15_, connection_5__6__14_, 
        connection_5__6__13_, connection_5__6__12_, connection_5__6__11_, 
        connection_5__6__10_, connection_5__6__9_, connection_5__6__8_, 
        connection_5__6__7_, connection_5__6__6_, connection_5__6__5_, 
        connection_5__6__4_, connection_5__6__3_, connection_5__6__2_, 
        connection_5__6__1_, connection_5__6__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[121:120]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_60 second_half_stages_4__group_sec_half_2__switch_sec_half_0__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__10_, 
        connection_valid_4__8_}), .i_data_bus({connection_4__10__31_, 
        connection_4__10__30_, connection_4__10__29_, connection_4__10__28_, 
        connection_4__10__27_, connection_4__10__26_, connection_4__10__25_, 
        connection_4__10__24_, connection_4__10__23_, connection_4__10__22_, 
        connection_4__10__21_, connection_4__10__20_, connection_4__10__19_, 
        connection_4__10__18_, connection_4__10__17_, connection_4__10__16_, 
        connection_4__10__15_, connection_4__10__14_, connection_4__10__13_, 
        connection_4__10__12_, connection_4__10__11_, connection_4__10__10_, 
        connection_4__10__9_, connection_4__10__8_, connection_4__10__7_, 
        connection_4__10__6_, connection_4__10__5_, connection_4__10__4_, 
        connection_4__10__3_, connection_4__10__2_, connection_4__10__1_, 
        connection_4__10__0_, connection_4__8__31_, connection_4__8__30_, 
        connection_4__8__29_, connection_4__8__28_, connection_4__8__27_, 
        connection_4__8__26_, connection_4__8__25_, connection_4__8__24_, 
        connection_4__8__23_, connection_4__8__22_, connection_4__8__21_, 
        connection_4__8__20_, connection_4__8__19_, connection_4__8__18_, 
        connection_4__8__17_, connection_4__8__16_, connection_4__8__15_, 
        connection_4__8__14_, connection_4__8__13_, connection_4__8__12_, 
        connection_4__8__11_, connection_4__8__10_, connection_4__8__9_, 
        connection_4__8__8_, connection_4__8__7_, connection_4__8__6_, 
        connection_4__8__5_, connection_4__8__4_, connection_4__8__3_, 
        connection_4__8__2_, connection_4__8__1_, connection_4__8__0_}), 
        .o_valid({connection_valid_5__9_, connection_valid_5__8_}), 
        .o_data_bus({connection_5__9__31_, connection_5__9__30_, 
        connection_5__9__29_, connection_5__9__28_, connection_5__9__27_, 
        connection_5__9__26_, connection_5__9__25_, connection_5__9__24_, 
        connection_5__9__23_, connection_5__9__22_, connection_5__9__21_, 
        connection_5__9__20_, connection_5__9__19_, connection_5__9__18_, 
        connection_5__9__17_, connection_5__9__16_, connection_5__9__15_, 
        connection_5__9__14_, connection_5__9__13_, connection_5__9__12_, 
        connection_5__9__11_, connection_5__9__10_, connection_5__9__9_, 
        connection_5__9__8_, connection_5__9__7_, connection_5__9__6_, 
        connection_5__9__5_, connection_5__9__4_, connection_5__9__3_, 
        connection_5__9__2_, connection_5__9__1_, connection_5__9__0_, 
        connection_5__8__31_, connection_5__8__30_, connection_5__8__29_, 
        connection_5__8__28_, connection_5__8__27_, connection_5__8__26_, 
        connection_5__8__25_, connection_5__8__24_, connection_5__8__23_, 
        connection_5__8__22_, connection_5__8__21_, connection_5__8__20_, 
        connection_5__8__19_, connection_5__8__18_, connection_5__8__17_, 
        connection_5__8__16_, connection_5__8__15_, connection_5__8__14_, 
        connection_5__8__13_, connection_5__8__12_, connection_5__8__11_, 
        connection_5__8__10_, connection_5__8__9_, connection_5__8__8_, 
        connection_5__8__7_, connection_5__8__6_, connection_5__8__5_, 
        connection_5__8__4_, connection_5__8__3_, connection_5__8__2_, 
        connection_5__8__1_, connection_5__8__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[119:118]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_59 second_half_stages_4__group_sec_half_2__switch_sec_half_1__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__11_, 
        connection_valid_4__9_}), .i_data_bus({connection_4__11__31_, 
        connection_4__11__30_, connection_4__11__29_, connection_4__11__28_, 
        connection_4__11__27_, connection_4__11__26_, connection_4__11__25_, 
        connection_4__11__24_, connection_4__11__23_, connection_4__11__22_, 
        connection_4__11__21_, connection_4__11__20_, connection_4__11__19_, 
        connection_4__11__18_, connection_4__11__17_, connection_4__11__16_, 
        connection_4__11__15_, connection_4__11__14_, connection_4__11__13_, 
        connection_4__11__12_, connection_4__11__11_, connection_4__11__10_, 
        connection_4__11__9_, connection_4__11__8_, connection_4__11__7_, 
        connection_4__11__6_, connection_4__11__5_, connection_4__11__4_, 
        connection_4__11__3_, connection_4__11__2_, connection_4__11__1_, 
        connection_4__11__0_, connection_4__9__31_, connection_4__9__30_, 
        connection_4__9__29_, connection_4__9__28_, connection_4__9__27_, 
        connection_4__9__26_, connection_4__9__25_, connection_4__9__24_, 
        connection_4__9__23_, connection_4__9__22_, connection_4__9__21_, 
        connection_4__9__20_, connection_4__9__19_, connection_4__9__18_, 
        connection_4__9__17_, connection_4__9__16_, connection_4__9__15_, 
        connection_4__9__14_, connection_4__9__13_, connection_4__9__12_, 
        connection_4__9__11_, connection_4__9__10_, connection_4__9__9_, 
        connection_4__9__8_, connection_4__9__7_, connection_4__9__6_, 
        connection_4__9__5_, connection_4__9__4_, connection_4__9__3_, 
        connection_4__9__2_, connection_4__9__1_, connection_4__9__0_}), 
        .o_valid({connection_valid_5__11_, connection_valid_5__10_}), 
        .o_data_bus({connection_5__11__31_, connection_5__11__30_, 
        connection_5__11__29_, connection_5__11__28_, connection_5__11__27_, 
        connection_5__11__26_, connection_5__11__25_, connection_5__11__24_, 
        connection_5__11__23_, connection_5__11__22_, connection_5__11__21_, 
        connection_5__11__20_, connection_5__11__19_, connection_5__11__18_, 
        connection_5__11__17_, connection_5__11__16_, connection_5__11__15_, 
        connection_5__11__14_, connection_5__11__13_, connection_5__11__12_, 
        connection_5__11__11_, connection_5__11__10_, connection_5__11__9_, 
        connection_5__11__8_, connection_5__11__7_, connection_5__11__6_, 
        connection_5__11__5_, connection_5__11__4_, connection_5__11__3_, 
        connection_5__11__2_, connection_5__11__1_, connection_5__11__0_, 
        connection_5__10__31_, connection_5__10__30_, connection_5__10__29_, 
        connection_5__10__28_, connection_5__10__27_, connection_5__10__26_, 
        connection_5__10__25_, connection_5__10__24_, connection_5__10__23_, 
        connection_5__10__22_, connection_5__10__21_, connection_5__10__20_, 
        connection_5__10__19_, connection_5__10__18_, connection_5__10__17_, 
        connection_5__10__16_, connection_5__10__15_, connection_5__10__14_, 
        connection_5__10__13_, connection_5__10__12_, connection_5__10__11_, 
        connection_5__10__10_, connection_5__10__9_, connection_5__10__8_, 
        connection_5__10__7_, connection_5__10__6_, connection_5__10__5_, 
        connection_5__10__4_, connection_5__10__3_, connection_5__10__2_, 
        connection_5__10__1_, connection_5__10__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[117:116]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_58 second_half_stages_4__group_sec_half_3__switch_sec_half_0__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__14_, 
        connection_valid_4__12_}), .i_data_bus({connection_4__14__31_, 
        connection_4__14__30_, connection_4__14__29_, connection_4__14__28_, 
        connection_4__14__27_, connection_4__14__26_, connection_4__14__25_, 
        connection_4__14__24_, connection_4__14__23_, connection_4__14__22_, 
        connection_4__14__21_, connection_4__14__20_, connection_4__14__19_, 
        connection_4__14__18_, connection_4__14__17_, connection_4__14__16_, 
        connection_4__14__15_, connection_4__14__14_, connection_4__14__13_, 
        connection_4__14__12_, connection_4__14__11_, connection_4__14__10_, 
        connection_4__14__9_, connection_4__14__8_, connection_4__14__7_, 
        connection_4__14__6_, connection_4__14__5_, connection_4__14__4_, 
        connection_4__14__3_, connection_4__14__2_, connection_4__14__1_, 
        connection_4__14__0_, connection_4__12__31_, connection_4__12__30_, 
        connection_4__12__29_, connection_4__12__28_, connection_4__12__27_, 
        connection_4__12__26_, connection_4__12__25_, connection_4__12__24_, 
        connection_4__12__23_, connection_4__12__22_, connection_4__12__21_, 
        connection_4__12__20_, connection_4__12__19_, connection_4__12__18_, 
        connection_4__12__17_, connection_4__12__16_, connection_4__12__15_, 
        connection_4__12__14_, connection_4__12__13_, connection_4__12__12_, 
        connection_4__12__11_, connection_4__12__10_, connection_4__12__9_, 
        connection_4__12__8_, connection_4__12__7_, connection_4__12__6_, 
        connection_4__12__5_, connection_4__12__4_, connection_4__12__3_, 
        connection_4__12__2_, connection_4__12__1_, connection_4__12__0_}), 
        .o_valid({connection_valid_5__13_, connection_valid_5__12_}), 
        .o_data_bus({connection_5__13__31_, connection_5__13__30_, 
        connection_5__13__29_, connection_5__13__28_, connection_5__13__27_, 
        connection_5__13__26_, connection_5__13__25_, connection_5__13__24_, 
        connection_5__13__23_, connection_5__13__22_, connection_5__13__21_, 
        connection_5__13__20_, connection_5__13__19_, connection_5__13__18_, 
        connection_5__13__17_, connection_5__13__16_, connection_5__13__15_, 
        connection_5__13__14_, connection_5__13__13_, connection_5__13__12_, 
        connection_5__13__11_, connection_5__13__10_, connection_5__13__9_, 
        connection_5__13__8_, connection_5__13__7_, connection_5__13__6_, 
        connection_5__13__5_, connection_5__13__4_, connection_5__13__3_, 
        connection_5__13__2_, connection_5__13__1_, connection_5__13__0_, 
        connection_5__12__31_, connection_5__12__30_, connection_5__12__29_, 
        connection_5__12__28_, connection_5__12__27_, connection_5__12__26_, 
        connection_5__12__25_, connection_5__12__24_, connection_5__12__23_, 
        connection_5__12__22_, connection_5__12__21_, connection_5__12__20_, 
        connection_5__12__19_, connection_5__12__18_, connection_5__12__17_, 
        connection_5__12__16_, connection_5__12__15_, connection_5__12__14_, 
        connection_5__12__13_, connection_5__12__12_, connection_5__12__11_, 
        connection_5__12__10_, connection_5__12__9_, connection_5__12__8_, 
        connection_5__12__7_, connection_5__12__6_, connection_5__12__5_, 
        connection_5__12__4_, connection_5__12__3_, connection_5__12__2_, 
        connection_5__12__1_, connection_5__12__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[115:114]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_57 second_half_stages_4__group_sec_half_3__switch_sec_half_1__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__15_, 
        connection_valid_4__13_}), .i_data_bus({connection_4__15__31_, 
        connection_4__15__30_, connection_4__15__29_, connection_4__15__28_, 
        connection_4__15__27_, connection_4__15__26_, connection_4__15__25_, 
        connection_4__15__24_, connection_4__15__23_, connection_4__15__22_, 
        connection_4__15__21_, connection_4__15__20_, connection_4__15__19_, 
        connection_4__15__18_, connection_4__15__17_, connection_4__15__16_, 
        connection_4__15__15_, connection_4__15__14_, connection_4__15__13_, 
        connection_4__15__12_, connection_4__15__11_, connection_4__15__10_, 
        connection_4__15__9_, connection_4__15__8_, connection_4__15__7_, 
        connection_4__15__6_, connection_4__15__5_, connection_4__15__4_, 
        connection_4__15__3_, connection_4__15__2_, connection_4__15__1_, 
        connection_4__15__0_, connection_4__13__31_, connection_4__13__30_, 
        connection_4__13__29_, connection_4__13__28_, connection_4__13__27_, 
        connection_4__13__26_, connection_4__13__25_, connection_4__13__24_, 
        connection_4__13__23_, connection_4__13__22_, connection_4__13__21_, 
        connection_4__13__20_, connection_4__13__19_, connection_4__13__18_, 
        connection_4__13__17_, connection_4__13__16_, connection_4__13__15_, 
        connection_4__13__14_, connection_4__13__13_, connection_4__13__12_, 
        connection_4__13__11_, connection_4__13__10_, connection_4__13__9_, 
        connection_4__13__8_, connection_4__13__7_, connection_4__13__6_, 
        connection_4__13__5_, connection_4__13__4_, connection_4__13__3_, 
        connection_4__13__2_, connection_4__13__1_, connection_4__13__0_}), 
        .o_valid({connection_valid_5__15_, connection_valid_5__14_}), 
        .o_data_bus({connection_5__15__31_, connection_5__15__30_, 
        connection_5__15__29_, connection_5__15__28_, connection_5__15__27_, 
        connection_5__15__26_, connection_5__15__25_, connection_5__15__24_, 
        connection_5__15__23_, connection_5__15__22_, connection_5__15__21_, 
        connection_5__15__20_, connection_5__15__19_, connection_5__15__18_, 
        connection_5__15__17_, connection_5__15__16_, connection_5__15__15_, 
        connection_5__15__14_, connection_5__15__13_, connection_5__15__12_, 
        connection_5__15__11_, connection_5__15__10_, connection_5__15__9_, 
        connection_5__15__8_, connection_5__15__7_, connection_5__15__6_, 
        connection_5__15__5_, connection_5__15__4_, connection_5__15__3_, 
        connection_5__15__2_, connection_5__15__1_, connection_5__15__0_, 
        connection_5__14__31_, connection_5__14__30_, connection_5__14__29_, 
        connection_5__14__28_, connection_5__14__27_, connection_5__14__26_, 
        connection_5__14__25_, connection_5__14__24_, connection_5__14__23_, 
        connection_5__14__22_, connection_5__14__21_, connection_5__14__20_, 
        connection_5__14__19_, connection_5__14__18_, connection_5__14__17_, 
        connection_5__14__16_, connection_5__14__15_, connection_5__14__14_, 
        connection_5__14__13_, connection_5__14__12_, connection_5__14__11_, 
        connection_5__14__10_, connection_5__14__9_, connection_5__14__8_, 
        connection_5__14__7_, connection_5__14__6_, connection_5__14__5_, 
        connection_5__14__4_, connection_5__14__3_, connection_5__14__2_, 
        connection_5__14__1_, connection_5__14__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[113:112]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_56 second_half_stages_4__group_sec_half_4__switch_sec_half_0__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__18_, 
        connection_valid_4__16_}), .i_data_bus({connection_4__18__31_, 
        connection_4__18__30_, connection_4__18__29_, connection_4__18__28_, 
        connection_4__18__27_, connection_4__18__26_, connection_4__18__25_, 
        connection_4__18__24_, connection_4__18__23_, connection_4__18__22_, 
        connection_4__18__21_, connection_4__18__20_, connection_4__18__19_, 
        connection_4__18__18_, connection_4__18__17_, connection_4__18__16_, 
        connection_4__18__15_, connection_4__18__14_, connection_4__18__13_, 
        connection_4__18__12_, connection_4__18__11_, connection_4__18__10_, 
        connection_4__18__9_, connection_4__18__8_, connection_4__18__7_, 
        connection_4__18__6_, connection_4__18__5_, connection_4__18__4_, 
        connection_4__18__3_, connection_4__18__2_, connection_4__18__1_, 
        connection_4__18__0_, connection_4__16__31_, connection_4__16__30_, 
        connection_4__16__29_, connection_4__16__28_, connection_4__16__27_, 
        connection_4__16__26_, connection_4__16__25_, connection_4__16__24_, 
        connection_4__16__23_, connection_4__16__22_, connection_4__16__21_, 
        connection_4__16__20_, connection_4__16__19_, connection_4__16__18_, 
        connection_4__16__17_, connection_4__16__16_, connection_4__16__15_, 
        connection_4__16__14_, connection_4__16__13_, connection_4__16__12_, 
        connection_4__16__11_, connection_4__16__10_, connection_4__16__9_, 
        connection_4__16__8_, connection_4__16__7_, connection_4__16__6_, 
        connection_4__16__5_, connection_4__16__4_, connection_4__16__3_, 
        connection_4__16__2_, connection_4__16__1_, connection_4__16__0_}), 
        .o_valid({connection_valid_5__17_, connection_valid_5__16_}), 
        .o_data_bus({connection_5__17__31_, connection_5__17__30_, 
        connection_5__17__29_, connection_5__17__28_, connection_5__17__27_, 
        connection_5__17__26_, connection_5__17__25_, connection_5__17__24_, 
        connection_5__17__23_, connection_5__17__22_, connection_5__17__21_, 
        connection_5__17__20_, connection_5__17__19_, connection_5__17__18_, 
        connection_5__17__17_, connection_5__17__16_, connection_5__17__15_, 
        connection_5__17__14_, connection_5__17__13_, connection_5__17__12_, 
        connection_5__17__11_, connection_5__17__10_, connection_5__17__9_, 
        connection_5__17__8_, connection_5__17__7_, connection_5__17__6_, 
        connection_5__17__5_, connection_5__17__4_, connection_5__17__3_, 
        connection_5__17__2_, connection_5__17__1_, connection_5__17__0_, 
        connection_5__16__31_, connection_5__16__30_, connection_5__16__29_, 
        connection_5__16__28_, connection_5__16__27_, connection_5__16__26_, 
        connection_5__16__25_, connection_5__16__24_, connection_5__16__23_, 
        connection_5__16__22_, connection_5__16__21_, connection_5__16__20_, 
        connection_5__16__19_, connection_5__16__18_, connection_5__16__17_, 
        connection_5__16__16_, connection_5__16__15_, connection_5__16__14_, 
        connection_5__16__13_, connection_5__16__12_, connection_5__16__11_, 
        connection_5__16__10_, connection_5__16__9_, connection_5__16__8_, 
        connection_5__16__7_, connection_5__16__6_, connection_5__16__5_, 
        connection_5__16__4_, connection_5__16__3_, connection_5__16__2_, 
        connection_5__16__1_, connection_5__16__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[111:110]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_55 second_half_stages_4__group_sec_half_4__switch_sec_half_1__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__19_, 
        connection_valid_4__17_}), .i_data_bus({connection_4__19__31_, 
        connection_4__19__30_, connection_4__19__29_, connection_4__19__28_, 
        connection_4__19__27_, connection_4__19__26_, connection_4__19__25_, 
        connection_4__19__24_, connection_4__19__23_, connection_4__19__22_, 
        connection_4__19__21_, connection_4__19__20_, connection_4__19__19_, 
        connection_4__19__18_, connection_4__19__17_, connection_4__19__16_, 
        connection_4__19__15_, connection_4__19__14_, connection_4__19__13_, 
        connection_4__19__12_, connection_4__19__11_, connection_4__19__10_, 
        connection_4__19__9_, connection_4__19__8_, connection_4__19__7_, 
        connection_4__19__6_, connection_4__19__5_, connection_4__19__4_, 
        connection_4__19__3_, connection_4__19__2_, connection_4__19__1_, 
        connection_4__19__0_, connection_4__17__31_, connection_4__17__30_, 
        connection_4__17__29_, connection_4__17__28_, connection_4__17__27_, 
        connection_4__17__26_, connection_4__17__25_, connection_4__17__24_, 
        connection_4__17__23_, connection_4__17__22_, connection_4__17__21_, 
        connection_4__17__20_, connection_4__17__19_, connection_4__17__18_, 
        connection_4__17__17_, connection_4__17__16_, connection_4__17__15_, 
        connection_4__17__14_, connection_4__17__13_, connection_4__17__12_, 
        connection_4__17__11_, connection_4__17__10_, connection_4__17__9_, 
        connection_4__17__8_, connection_4__17__7_, connection_4__17__6_, 
        connection_4__17__5_, connection_4__17__4_, connection_4__17__3_, 
        connection_4__17__2_, connection_4__17__1_, connection_4__17__0_}), 
        .o_valid({connection_valid_5__19_, connection_valid_5__18_}), 
        .o_data_bus({connection_5__19__31_, connection_5__19__30_, 
        connection_5__19__29_, connection_5__19__28_, connection_5__19__27_, 
        connection_5__19__26_, connection_5__19__25_, connection_5__19__24_, 
        connection_5__19__23_, connection_5__19__22_, connection_5__19__21_, 
        connection_5__19__20_, connection_5__19__19_, connection_5__19__18_, 
        connection_5__19__17_, connection_5__19__16_, connection_5__19__15_, 
        connection_5__19__14_, connection_5__19__13_, connection_5__19__12_, 
        connection_5__19__11_, connection_5__19__10_, connection_5__19__9_, 
        connection_5__19__8_, connection_5__19__7_, connection_5__19__6_, 
        connection_5__19__5_, connection_5__19__4_, connection_5__19__3_, 
        connection_5__19__2_, connection_5__19__1_, connection_5__19__0_, 
        connection_5__18__31_, connection_5__18__30_, connection_5__18__29_, 
        connection_5__18__28_, connection_5__18__27_, connection_5__18__26_, 
        connection_5__18__25_, connection_5__18__24_, connection_5__18__23_, 
        connection_5__18__22_, connection_5__18__21_, connection_5__18__20_, 
        connection_5__18__19_, connection_5__18__18_, connection_5__18__17_, 
        connection_5__18__16_, connection_5__18__15_, connection_5__18__14_, 
        connection_5__18__13_, connection_5__18__12_, connection_5__18__11_, 
        connection_5__18__10_, connection_5__18__9_, connection_5__18__8_, 
        connection_5__18__7_, connection_5__18__6_, connection_5__18__5_, 
        connection_5__18__4_, connection_5__18__3_, connection_5__18__2_, 
        connection_5__18__1_, connection_5__18__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[109:108]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_54 second_half_stages_4__group_sec_half_5__switch_sec_half_0__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__22_, 
        connection_valid_4__20_}), .i_data_bus({connection_4__22__31_, 
        connection_4__22__30_, connection_4__22__29_, connection_4__22__28_, 
        connection_4__22__27_, connection_4__22__26_, connection_4__22__25_, 
        connection_4__22__24_, connection_4__22__23_, connection_4__22__22_, 
        connection_4__22__21_, connection_4__22__20_, connection_4__22__19_, 
        connection_4__22__18_, connection_4__22__17_, connection_4__22__16_, 
        connection_4__22__15_, connection_4__22__14_, connection_4__22__13_, 
        connection_4__22__12_, connection_4__22__11_, connection_4__22__10_, 
        connection_4__22__9_, connection_4__22__8_, connection_4__22__7_, 
        connection_4__22__6_, connection_4__22__5_, connection_4__22__4_, 
        connection_4__22__3_, connection_4__22__2_, connection_4__22__1_, 
        connection_4__22__0_, connection_4__20__31_, connection_4__20__30_, 
        connection_4__20__29_, connection_4__20__28_, connection_4__20__27_, 
        connection_4__20__26_, connection_4__20__25_, connection_4__20__24_, 
        connection_4__20__23_, connection_4__20__22_, connection_4__20__21_, 
        connection_4__20__20_, connection_4__20__19_, connection_4__20__18_, 
        connection_4__20__17_, connection_4__20__16_, connection_4__20__15_, 
        connection_4__20__14_, connection_4__20__13_, connection_4__20__12_, 
        connection_4__20__11_, connection_4__20__10_, connection_4__20__9_, 
        connection_4__20__8_, connection_4__20__7_, connection_4__20__6_, 
        connection_4__20__5_, connection_4__20__4_, connection_4__20__3_, 
        connection_4__20__2_, connection_4__20__1_, connection_4__20__0_}), 
        .o_valid({connection_valid_5__21_, connection_valid_5__20_}), 
        .o_data_bus({connection_5__21__31_, connection_5__21__30_, 
        connection_5__21__29_, connection_5__21__28_, connection_5__21__27_, 
        connection_5__21__26_, connection_5__21__25_, connection_5__21__24_, 
        connection_5__21__23_, connection_5__21__22_, connection_5__21__21_, 
        connection_5__21__20_, connection_5__21__19_, connection_5__21__18_, 
        connection_5__21__17_, connection_5__21__16_, connection_5__21__15_, 
        connection_5__21__14_, connection_5__21__13_, connection_5__21__12_, 
        connection_5__21__11_, connection_5__21__10_, connection_5__21__9_, 
        connection_5__21__8_, connection_5__21__7_, connection_5__21__6_, 
        connection_5__21__5_, connection_5__21__4_, connection_5__21__3_, 
        connection_5__21__2_, connection_5__21__1_, connection_5__21__0_, 
        connection_5__20__31_, connection_5__20__30_, connection_5__20__29_, 
        connection_5__20__28_, connection_5__20__27_, connection_5__20__26_, 
        connection_5__20__25_, connection_5__20__24_, connection_5__20__23_, 
        connection_5__20__22_, connection_5__20__21_, connection_5__20__20_, 
        connection_5__20__19_, connection_5__20__18_, connection_5__20__17_, 
        connection_5__20__16_, connection_5__20__15_, connection_5__20__14_, 
        connection_5__20__13_, connection_5__20__12_, connection_5__20__11_, 
        connection_5__20__10_, connection_5__20__9_, connection_5__20__8_, 
        connection_5__20__7_, connection_5__20__6_, connection_5__20__5_, 
        connection_5__20__4_, connection_5__20__3_, connection_5__20__2_, 
        connection_5__20__1_, connection_5__20__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[107:106]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_53 second_half_stages_4__group_sec_half_5__switch_sec_half_1__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__23_, 
        connection_valid_4__21_}), .i_data_bus({connection_4__23__31_, 
        connection_4__23__30_, connection_4__23__29_, connection_4__23__28_, 
        connection_4__23__27_, connection_4__23__26_, connection_4__23__25_, 
        connection_4__23__24_, connection_4__23__23_, connection_4__23__22_, 
        connection_4__23__21_, connection_4__23__20_, connection_4__23__19_, 
        connection_4__23__18_, connection_4__23__17_, connection_4__23__16_, 
        connection_4__23__15_, connection_4__23__14_, connection_4__23__13_, 
        connection_4__23__12_, connection_4__23__11_, connection_4__23__10_, 
        connection_4__23__9_, connection_4__23__8_, connection_4__23__7_, 
        connection_4__23__6_, connection_4__23__5_, connection_4__23__4_, 
        connection_4__23__3_, connection_4__23__2_, connection_4__23__1_, 
        connection_4__23__0_, connection_4__21__31_, connection_4__21__30_, 
        connection_4__21__29_, connection_4__21__28_, connection_4__21__27_, 
        connection_4__21__26_, connection_4__21__25_, connection_4__21__24_, 
        connection_4__21__23_, connection_4__21__22_, connection_4__21__21_, 
        connection_4__21__20_, connection_4__21__19_, connection_4__21__18_, 
        connection_4__21__17_, connection_4__21__16_, connection_4__21__15_, 
        connection_4__21__14_, connection_4__21__13_, connection_4__21__12_, 
        connection_4__21__11_, connection_4__21__10_, connection_4__21__9_, 
        connection_4__21__8_, connection_4__21__7_, connection_4__21__6_, 
        connection_4__21__5_, connection_4__21__4_, connection_4__21__3_, 
        connection_4__21__2_, connection_4__21__1_, connection_4__21__0_}), 
        .o_valid({connection_valid_5__23_, connection_valid_5__22_}), 
        .o_data_bus({connection_5__23__31_, connection_5__23__30_, 
        connection_5__23__29_, connection_5__23__28_, connection_5__23__27_, 
        connection_5__23__26_, connection_5__23__25_, connection_5__23__24_, 
        connection_5__23__23_, connection_5__23__22_, connection_5__23__21_, 
        connection_5__23__20_, connection_5__23__19_, connection_5__23__18_, 
        connection_5__23__17_, connection_5__23__16_, connection_5__23__15_, 
        connection_5__23__14_, connection_5__23__13_, connection_5__23__12_, 
        connection_5__23__11_, connection_5__23__10_, connection_5__23__9_, 
        connection_5__23__8_, connection_5__23__7_, connection_5__23__6_, 
        connection_5__23__5_, connection_5__23__4_, connection_5__23__3_, 
        connection_5__23__2_, connection_5__23__1_, connection_5__23__0_, 
        connection_5__22__31_, connection_5__22__30_, connection_5__22__29_, 
        connection_5__22__28_, connection_5__22__27_, connection_5__22__26_, 
        connection_5__22__25_, connection_5__22__24_, connection_5__22__23_, 
        connection_5__22__22_, connection_5__22__21_, connection_5__22__20_, 
        connection_5__22__19_, connection_5__22__18_, connection_5__22__17_, 
        connection_5__22__16_, connection_5__22__15_, connection_5__22__14_, 
        connection_5__22__13_, connection_5__22__12_, connection_5__22__11_, 
        connection_5__22__10_, connection_5__22__9_, connection_5__22__8_, 
        connection_5__22__7_, connection_5__22__6_, connection_5__22__5_, 
        connection_5__22__4_, connection_5__22__3_, connection_5__22__2_, 
        connection_5__22__1_, connection_5__22__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[105:104]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_52 second_half_stages_4__group_sec_half_6__switch_sec_half_0__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__26_, 
        connection_valid_4__24_}), .i_data_bus({connection_4__26__31_, 
        connection_4__26__30_, connection_4__26__29_, connection_4__26__28_, 
        connection_4__26__27_, connection_4__26__26_, connection_4__26__25_, 
        connection_4__26__24_, connection_4__26__23_, connection_4__26__22_, 
        connection_4__26__21_, connection_4__26__20_, connection_4__26__19_, 
        connection_4__26__18_, connection_4__26__17_, connection_4__26__16_, 
        connection_4__26__15_, connection_4__26__14_, connection_4__26__13_, 
        connection_4__26__12_, connection_4__26__11_, connection_4__26__10_, 
        connection_4__26__9_, connection_4__26__8_, connection_4__26__7_, 
        connection_4__26__6_, connection_4__26__5_, connection_4__26__4_, 
        connection_4__26__3_, connection_4__26__2_, connection_4__26__1_, 
        connection_4__26__0_, connection_4__24__31_, connection_4__24__30_, 
        connection_4__24__29_, connection_4__24__28_, connection_4__24__27_, 
        connection_4__24__26_, connection_4__24__25_, connection_4__24__24_, 
        connection_4__24__23_, connection_4__24__22_, connection_4__24__21_, 
        connection_4__24__20_, connection_4__24__19_, connection_4__24__18_, 
        connection_4__24__17_, connection_4__24__16_, connection_4__24__15_, 
        connection_4__24__14_, connection_4__24__13_, connection_4__24__12_, 
        connection_4__24__11_, connection_4__24__10_, connection_4__24__9_, 
        connection_4__24__8_, connection_4__24__7_, connection_4__24__6_, 
        connection_4__24__5_, connection_4__24__4_, connection_4__24__3_, 
        connection_4__24__2_, connection_4__24__1_, connection_4__24__0_}), 
        .o_valid({connection_valid_5__25_, connection_valid_5__24_}), 
        .o_data_bus({connection_5__25__31_, connection_5__25__30_, 
        connection_5__25__29_, connection_5__25__28_, connection_5__25__27_, 
        connection_5__25__26_, connection_5__25__25_, connection_5__25__24_, 
        connection_5__25__23_, connection_5__25__22_, connection_5__25__21_, 
        connection_5__25__20_, connection_5__25__19_, connection_5__25__18_, 
        connection_5__25__17_, connection_5__25__16_, connection_5__25__15_, 
        connection_5__25__14_, connection_5__25__13_, connection_5__25__12_, 
        connection_5__25__11_, connection_5__25__10_, connection_5__25__9_, 
        connection_5__25__8_, connection_5__25__7_, connection_5__25__6_, 
        connection_5__25__5_, connection_5__25__4_, connection_5__25__3_, 
        connection_5__25__2_, connection_5__25__1_, connection_5__25__0_, 
        connection_5__24__31_, connection_5__24__30_, connection_5__24__29_, 
        connection_5__24__28_, connection_5__24__27_, connection_5__24__26_, 
        connection_5__24__25_, connection_5__24__24_, connection_5__24__23_, 
        connection_5__24__22_, connection_5__24__21_, connection_5__24__20_, 
        connection_5__24__19_, connection_5__24__18_, connection_5__24__17_, 
        connection_5__24__16_, connection_5__24__15_, connection_5__24__14_, 
        connection_5__24__13_, connection_5__24__12_, connection_5__24__11_, 
        connection_5__24__10_, connection_5__24__9_, connection_5__24__8_, 
        connection_5__24__7_, connection_5__24__6_, connection_5__24__5_, 
        connection_5__24__4_, connection_5__24__3_, connection_5__24__2_, 
        connection_5__24__1_, connection_5__24__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[103:102]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_51 second_half_stages_4__group_sec_half_6__switch_sec_half_1__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__27_, 
        connection_valid_4__25_}), .i_data_bus({connection_4__27__31_, 
        connection_4__27__30_, connection_4__27__29_, connection_4__27__28_, 
        connection_4__27__27_, connection_4__27__26_, connection_4__27__25_, 
        connection_4__27__24_, connection_4__27__23_, connection_4__27__22_, 
        connection_4__27__21_, connection_4__27__20_, connection_4__27__19_, 
        connection_4__27__18_, connection_4__27__17_, connection_4__27__16_, 
        connection_4__27__15_, connection_4__27__14_, connection_4__27__13_, 
        connection_4__27__12_, connection_4__27__11_, connection_4__27__10_, 
        connection_4__27__9_, connection_4__27__8_, connection_4__27__7_, 
        connection_4__27__6_, connection_4__27__5_, connection_4__27__4_, 
        connection_4__27__3_, connection_4__27__2_, connection_4__27__1_, 
        connection_4__27__0_, connection_4__25__31_, connection_4__25__30_, 
        connection_4__25__29_, connection_4__25__28_, connection_4__25__27_, 
        connection_4__25__26_, connection_4__25__25_, connection_4__25__24_, 
        connection_4__25__23_, connection_4__25__22_, connection_4__25__21_, 
        connection_4__25__20_, connection_4__25__19_, connection_4__25__18_, 
        connection_4__25__17_, connection_4__25__16_, connection_4__25__15_, 
        connection_4__25__14_, connection_4__25__13_, connection_4__25__12_, 
        connection_4__25__11_, connection_4__25__10_, connection_4__25__9_, 
        connection_4__25__8_, connection_4__25__7_, connection_4__25__6_, 
        connection_4__25__5_, connection_4__25__4_, connection_4__25__3_, 
        connection_4__25__2_, connection_4__25__1_, connection_4__25__0_}), 
        .o_valid({connection_valid_5__27_, connection_valid_5__26_}), 
        .o_data_bus({connection_5__27__31_, connection_5__27__30_, 
        connection_5__27__29_, connection_5__27__28_, connection_5__27__27_, 
        connection_5__27__26_, connection_5__27__25_, connection_5__27__24_, 
        connection_5__27__23_, connection_5__27__22_, connection_5__27__21_, 
        connection_5__27__20_, connection_5__27__19_, connection_5__27__18_, 
        connection_5__27__17_, connection_5__27__16_, connection_5__27__15_, 
        connection_5__27__14_, connection_5__27__13_, connection_5__27__12_, 
        connection_5__27__11_, connection_5__27__10_, connection_5__27__9_, 
        connection_5__27__8_, connection_5__27__7_, connection_5__27__6_, 
        connection_5__27__5_, connection_5__27__4_, connection_5__27__3_, 
        connection_5__27__2_, connection_5__27__1_, connection_5__27__0_, 
        connection_5__26__31_, connection_5__26__30_, connection_5__26__29_, 
        connection_5__26__28_, connection_5__26__27_, connection_5__26__26_, 
        connection_5__26__25_, connection_5__26__24_, connection_5__26__23_, 
        connection_5__26__22_, connection_5__26__21_, connection_5__26__20_, 
        connection_5__26__19_, connection_5__26__18_, connection_5__26__17_, 
        connection_5__26__16_, connection_5__26__15_, connection_5__26__14_, 
        connection_5__26__13_, connection_5__26__12_, connection_5__26__11_, 
        connection_5__26__10_, connection_5__26__9_, connection_5__26__8_, 
        connection_5__26__7_, connection_5__26__6_, connection_5__26__5_, 
        connection_5__26__4_, connection_5__26__3_, connection_5__26__2_, 
        connection_5__26__1_, connection_5__26__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[101:100]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_50 second_half_stages_4__group_sec_half_7__switch_sec_half_0__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__30_, 
        connection_valid_4__28_}), .i_data_bus({connection_4__30__31_, 
        connection_4__30__30_, connection_4__30__29_, connection_4__30__28_, 
        connection_4__30__27_, connection_4__30__26_, connection_4__30__25_, 
        connection_4__30__24_, connection_4__30__23_, connection_4__30__22_, 
        connection_4__30__21_, connection_4__30__20_, connection_4__30__19_, 
        connection_4__30__18_, connection_4__30__17_, connection_4__30__16_, 
        connection_4__30__15_, connection_4__30__14_, connection_4__30__13_, 
        connection_4__30__12_, connection_4__30__11_, connection_4__30__10_, 
        connection_4__30__9_, connection_4__30__8_, connection_4__30__7_, 
        connection_4__30__6_, connection_4__30__5_, connection_4__30__4_, 
        connection_4__30__3_, connection_4__30__2_, connection_4__30__1_, 
        connection_4__30__0_, connection_4__28__31_, connection_4__28__30_, 
        connection_4__28__29_, connection_4__28__28_, connection_4__28__27_, 
        connection_4__28__26_, connection_4__28__25_, connection_4__28__24_, 
        connection_4__28__23_, connection_4__28__22_, connection_4__28__21_, 
        connection_4__28__20_, connection_4__28__19_, connection_4__28__18_, 
        connection_4__28__17_, connection_4__28__16_, connection_4__28__15_, 
        connection_4__28__14_, connection_4__28__13_, connection_4__28__12_, 
        connection_4__28__11_, connection_4__28__10_, connection_4__28__9_, 
        connection_4__28__8_, connection_4__28__7_, connection_4__28__6_, 
        connection_4__28__5_, connection_4__28__4_, connection_4__28__3_, 
        connection_4__28__2_, connection_4__28__1_, connection_4__28__0_}), 
        .o_valid({connection_valid_5__29_, connection_valid_5__28_}), 
        .o_data_bus({connection_5__29__31_, connection_5__29__30_, 
        connection_5__29__29_, connection_5__29__28_, connection_5__29__27_, 
        connection_5__29__26_, connection_5__29__25_, connection_5__29__24_, 
        connection_5__29__23_, connection_5__29__22_, connection_5__29__21_, 
        connection_5__29__20_, connection_5__29__19_, connection_5__29__18_, 
        connection_5__29__17_, connection_5__29__16_, connection_5__29__15_, 
        connection_5__29__14_, connection_5__29__13_, connection_5__29__12_, 
        connection_5__29__11_, connection_5__29__10_, connection_5__29__9_, 
        connection_5__29__8_, connection_5__29__7_, connection_5__29__6_, 
        connection_5__29__5_, connection_5__29__4_, connection_5__29__3_, 
        connection_5__29__2_, connection_5__29__1_, connection_5__29__0_, 
        connection_5__28__31_, connection_5__28__30_, connection_5__28__29_, 
        connection_5__28__28_, connection_5__28__27_, connection_5__28__26_, 
        connection_5__28__25_, connection_5__28__24_, connection_5__28__23_, 
        connection_5__28__22_, connection_5__28__21_, connection_5__28__20_, 
        connection_5__28__19_, connection_5__28__18_, connection_5__28__17_, 
        connection_5__28__16_, connection_5__28__15_, connection_5__28__14_, 
        connection_5__28__13_, connection_5__28__12_, connection_5__28__11_, 
        connection_5__28__10_, connection_5__28__9_, connection_5__28__8_, 
        connection_5__28__7_, connection_5__28__6_, connection_5__28__5_, 
        connection_5__28__4_, connection_5__28__3_, connection_5__28__2_, 
        connection_5__28__1_, connection_5__28__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[99:98]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_49 second_half_stages_4__group_sec_half_7__switch_sec_half_1__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__31_, 
        connection_valid_4__29_}), .i_data_bus({connection_4__31__31_, 
        connection_4__31__30_, connection_4__31__29_, connection_4__31__28_, 
        connection_4__31__27_, connection_4__31__26_, connection_4__31__25_, 
        connection_4__31__24_, connection_4__31__23_, connection_4__31__22_, 
        connection_4__31__21_, connection_4__31__20_, connection_4__31__19_, 
        connection_4__31__18_, connection_4__31__17_, connection_4__31__16_, 
        connection_4__31__15_, connection_4__31__14_, connection_4__31__13_, 
        connection_4__31__12_, connection_4__31__11_, connection_4__31__10_, 
        connection_4__31__9_, connection_4__31__8_, connection_4__31__7_, 
        connection_4__31__6_, connection_4__31__5_, connection_4__31__4_, 
        connection_4__31__3_, connection_4__31__2_, connection_4__31__1_, 
        connection_4__31__0_, connection_4__29__31_, connection_4__29__30_, 
        connection_4__29__29_, connection_4__29__28_, connection_4__29__27_, 
        connection_4__29__26_, connection_4__29__25_, connection_4__29__24_, 
        connection_4__29__23_, connection_4__29__22_, connection_4__29__21_, 
        connection_4__29__20_, connection_4__29__19_, connection_4__29__18_, 
        connection_4__29__17_, connection_4__29__16_, connection_4__29__15_, 
        connection_4__29__14_, connection_4__29__13_, connection_4__29__12_, 
        connection_4__29__11_, connection_4__29__10_, connection_4__29__9_, 
        connection_4__29__8_, connection_4__29__7_, connection_4__29__6_, 
        connection_4__29__5_, connection_4__29__4_, connection_4__29__3_, 
        connection_4__29__2_, connection_4__29__1_, connection_4__29__0_}), 
        .o_valid({connection_valid_5__31_, connection_valid_5__30_}), 
        .o_data_bus({connection_5__31__31_, connection_5__31__30_, 
        connection_5__31__29_, connection_5__31__28_, connection_5__31__27_, 
        connection_5__31__26_, connection_5__31__25_, connection_5__31__24_, 
        connection_5__31__23_, connection_5__31__22_, connection_5__31__21_, 
        connection_5__31__20_, connection_5__31__19_, connection_5__31__18_, 
        connection_5__31__17_, connection_5__31__16_, connection_5__31__15_, 
        connection_5__31__14_, connection_5__31__13_, connection_5__31__12_, 
        connection_5__31__11_, connection_5__31__10_, connection_5__31__9_, 
        connection_5__31__8_, connection_5__31__7_, connection_5__31__6_, 
        connection_5__31__5_, connection_5__31__4_, connection_5__31__3_, 
        connection_5__31__2_, connection_5__31__1_, connection_5__31__0_, 
        connection_5__30__31_, connection_5__30__30_, connection_5__30__29_, 
        connection_5__30__28_, connection_5__30__27_, connection_5__30__26_, 
        connection_5__30__25_, connection_5__30__24_, connection_5__30__23_, 
        connection_5__30__22_, connection_5__30__21_, connection_5__30__20_, 
        connection_5__30__19_, connection_5__30__18_, connection_5__30__17_, 
        connection_5__30__16_, connection_5__30__15_, connection_5__30__14_, 
        connection_5__30__13_, connection_5__30__12_, connection_5__30__11_, 
        connection_5__30__10_, connection_5__30__9_, connection_5__30__8_, 
        connection_5__30__7_, connection_5__30__6_, connection_5__30__5_, 
        connection_5__30__4_, connection_5__30__3_, connection_5__30__2_, 
        connection_5__30__1_, connection_5__30__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[97:96]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_48 second_half_stages_5__group_sec_half_0__switch_sec_half_0__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__4_, 
        connection_valid_5__0_}), .i_data_bus({connection_5__4__31_, 
        connection_5__4__30_, connection_5__4__29_, connection_5__4__28_, 
        connection_5__4__27_, connection_5__4__26_, connection_5__4__25_, 
        connection_5__4__24_, connection_5__4__23_, connection_5__4__22_, 
        connection_5__4__21_, connection_5__4__20_, connection_5__4__19_, 
        connection_5__4__18_, connection_5__4__17_, connection_5__4__16_, 
        connection_5__4__15_, connection_5__4__14_, connection_5__4__13_, 
        connection_5__4__12_, connection_5__4__11_, connection_5__4__10_, 
        connection_5__4__9_, connection_5__4__8_, connection_5__4__7_, 
        connection_5__4__6_, connection_5__4__5_, connection_5__4__4_, 
        connection_5__4__3_, connection_5__4__2_, connection_5__4__1_, 
        connection_5__4__0_, connection_5__0__31_, connection_5__0__30_, 
        connection_5__0__29_, connection_5__0__28_, connection_5__0__27_, 
        connection_5__0__26_, connection_5__0__25_, connection_5__0__24_, 
        connection_5__0__23_, connection_5__0__22_, connection_5__0__21_, 
        connection_5__0__20_, connection_5__0__19_, connection_5__0__18_, 
        connection_5__0__17_, connection_5__0__16_, connection_5__0__15_, 
        connection_5__0__14_, connection_5__0__13_, connection_5__0__12_, 
        connection_5__0__11_, connection_5__0__10_, connection_5__0__9_, 
        connection_5__0__8_, connection_5__0__7_, connection_5__0__6_, 
        connection_5__0__5_, connection_5__0__4_, connection_5__0__3_, 
        connection_5__0__2_, connection_5__0__1_, connection_5__0__0_}), 
        .o_valid({connection_valid_6__1_, connection_valid_6__0_}), 
        .o_data_bus({connection_6__1__31_, connection_6__1__30_, 
        connection_6__1__29_, connection_6__1__28_, connection_6__1__27_, 
        connection_6__1__26_, connection_6__1__25_, connection_6__1__24_, 
        connection_6__1__23_, connection_6__1__22_, connection_6__1__21_, 
        connection_6__1__20_, connection_6__1__19_, connection_6__1__18_, 
        connection_6__1__17_, connection_6__1__16_, connection_6__1__15_, 
        connection_6__1__14_, connection_6__1__13_, connection_6__1__12_, 
        connection_6__1__11_, connection_6__1__10_, connection_6__1__9_, 
        connection_6__1__8_, connection_6__1__7_, connection_6__1__6_, 
        connection_6__1__5_, connection_6__1__4_, connection_6__1__3_, 
        connection_6__1__2_, connection_6__1__1_, connection_6__1__0_, 
        connection_6__0__31_, connection_6__0__30_, connection_6__0__29_, 
        connection_6__0__28_, connection_6__0__27_, connection_6__0__26_, 
        connection_6__0__25_, connection_6__0__24_, connection_6__0__23_, 
        connection_6__0__22_, connection_6__0__21_, connection_6__0__20_, 
        connection_6__0__19_, connection_6__0__18_, connection_6__0__17_, 
        connection_6__0__16_, connection_6__0__15_, connection_6__0__14_, 
        connection_6__0__13_, connection_6__0__12_, connection_6__0__11_, 
        connection_6__0__10_, connection_6__0__9_, connection_6__0__8_, 
        connection_6__0__7_, connection_6__0__6_, connection_6__0__5_, 
        connection_6__0__4_, connection_6__0__3_, connection_6__0__2_, 
        connection_6__0__1_, connection_6__0__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[95:94]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_47 second_half_stages_5__group_sec_half_0__switch_sec_half_1__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__5_, 
        connection_valid_5__1_}), .i_data_bus({connection_5__5__31_, 
        connection_5__5__30_, connection_5__5__29_, connection_5__5__28_, 
        connection_5__5__27_, connection_5__5__26_, connection_5__5__25_, 
        connection_5__5__24_, connection_5__5__23_, connection_5__5__22_, 
        connection_5__5__21_, connection_5__5__20_, connection_5__5__19_, 
        connection_5__5__18_, connection_5__5__17_, connection_5__5__16_, 
        connection_5__5__15_, connection_5__5__14_, connection_5__5__13_, 
        connection_5__5__12_, connection_5__5__11_, connection_5__5__10_, 
        connection_5__5__9_, connection_5__5__8_, connection_5__5__7_, 
        connection_5__5__6_, connection_5__5__5_, connection_5__5__4_, 
        connection_5__5__3_, connection_5__5__2_, connection_5__5__1_, 
        connection_5__5__0_, connection_5__1__31_, connection_5__1__30_, 
        connection_5__1__29_, connection_5__1__28_, connection_5__1__27_, 
        connection_5__1__26_, connection_5__1__25_, connection_5__1__24_, 
        connection_5__1__23_, connection_5__1__22_, connection_5__1__21_, 
        connection_5__1__20_, connection_5__1__19_, connection_5__1__18_, 
        connection_5__1__17_, connection_5__1__16_, connection_5__1__15_, 
        connection_5__1__14_, connection_5__1__13_, connection_5__1__12_, 
        connection_5__1__11_, connection_5__1__10_, connection_5__1__9_, 
        connection_5__1__8_, connection_5__1__7_, connection_5__1__6_, 
        connection_5__1__5_, connection_5__1__4_, connection_5__1__3_, 
        connection_5__1__2_, connection_5__1__1_, connection_5__1__0_}), 
        .o_valid({connection_valid_6__3_, connection_valid_6__2_}), 
        .o_data_bus({connection_6__3__31_, connection_6__3__30_, 
        connection_6__3__29_, connection_6__3__28_, connection_6__3__27_, 
        connection_6__3__26_, connection_6__3__25_, connection_6__3__24_, 
        connection_6__3__23_, connection_6__3__22_, connection_6__3__21_, 
        connection_6__3__20_, connection_6__3__19_, connection_6__3__18_, 
        connection_6__3__17_, connection_6__3__16_, connection_6__3__15_, 
        connection_6__3__14_, connection_6__3__13_, connection_6__3__12_, 
        connection_6__3__11_, connection_6__3__10_, connection_6__3__9_, 
        connection_6__3__8_, connection_6__3__7_, connection_6__3__6_, 
        connection_6__3__5_, connection_6__3__4_, connection_6__3__3_, 
        connection_6__3__2_, connection_6__3__1_, connection_6__3__0_, 
        connection_6__2__31_, connection_6__2__30_, connection_6__2__29_, 
        connection_6__2__28_, connection_6__2__27_, connection_6__2__26_, 
        connection_6__2__25_, connection_6__2__24_, connection_6__2__23_, 
        connection_6__2__22_, connection_6__2__21_, connection_6__2__20_, 
        connection_6__2__19_, connection_6__2__18_, connection_6__2__17_, 
        connection_6__2__16_, connection_6__2__15_, connection_6__2__14_, 
        connection_6__2__13_, connection_6__2__12_, connection_6__2__11_, 
        connection_6__2__10_, connection_6__2__9_, connection_6__2__8_, 
        connection_6__2__7_, connection_6__2__6_, connection_6__2__5_, 
        connection_6__2__4_, connection_6__2__3_, connection_6__2__2_, 
        connection_6__2__1_, connection_6__2__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[93:92]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_46 second_half_stages_5__group_sec_half_0__switch_sec_half_2__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__6_, 
        connection_valid_5__2_}), .i_data_bus({connection_5__6__31_, 
        connection_5__6__30_, connection_5__6__29_, connection_5__6__28_, 
        connection_5__6__27_, connection_5__6__26_, connection_5__6__25_, 
        connection_5__6__24_, connection_5__6__23_, connection_5__6__22_, 
        connection_5__6__21_, connection_5__6__20_, connection_5__6__19_, 
        connection_5__6__18_, connection_5__6__17_, connection_5__6__16_, 
        connection_5__6__15_, connection_5__6__14_, connection_5__6__13_, 
        connection_5__6__12_, connection_5__6__11_, connection_5__6__10_, 
        connection_5__6__9_, connection_5__6__8_, connection_5__6__7_, 
        connection_5__6__6_, connection_5__6__5_, connection_5__6__4_, 
        connection_5__6__3_, connection_5__6__2_, connection_5__6__1_, 
        connection_5__6__0_, connection_5__2__31_, connection_5__2__30_, 
        connection_5__2__29_, connection_5__2__28_, connection_5__2__27_, 
        connection_5__2__26_, connection_5__2__25_, connection_5__2__24_, 
        connection_5__2__23_, connection_5__2__22_, connection_5__2__21_, 
        connection_5__2__20_, connection_5__2__19_, connection_5__2__18_, 
        connection_5__2__17_, connection_5__2__16_, connection_5__2__15_, 
        connection_5__2__14_, connection_5__2__13_, connection_5__2__12_, 
        connection_5__2__11_, connection_5__2__10_, connection_5__2__9_, 
        connection_5__2__8_, connection_5__2__7_, connection_5__2__6_, 
        connection_5__2__5_, connection_5__2__4_, connection_5__2__3_, 
        connection_5__2__2_, connection_5__2__1_, connection_5__2__0_}), 
        .o_valid({connection_valid_6__5_, connection_valid_6__4_}), 
        .o_data_bus({connection_6__5__31_, connection_6__5__30_, 
        connection_6__5__29_, connection_6__5__28_, connection_6__5__27_, 
        connection_6__5__26_, connection_6__5__25_, connection_6__5__24_, 
        connection_6__5__23_, connection_6__5__22_, connection_6__5__21_, 
        connection_6__5__20_, connection_6__5__19_, connection_6__5__18_, 
        connection_6__5__17_, connection_6__5__16_, connection_6__5__15_, 
        connection_6__5__14_, connection_6__5__13_, connection_6__5__12_, 
        connection_6__5__11_, connection_6__5__10_, connection_6__5__9_, 
        connection_6__5__8_, connection_6__5__7_, connection_6__5__6_, 
        connection_6__5__5_, connection_6__5__4_, connection_6__5__3_, 
        connection_6__5__2_, connection_6__5__1_, connection_6__5__0_, 
        connection_6__4__31_, connection_6__4__30_, connection_6__4__29_, 
        connection_6__4__28_, connection_6__4__27_, connection_6__4__26_, 
        connection_6__4__25_, connection_6__4__24_, connection_6__4__23_, 
        connection_6__4__22_, connection_6__4__21_, connection_6__4__20_, 
        connection_6__4__19_, connection_6__4__18_, connection_6__4__17_, 
        connection_6__4__16_, connection_6__4__15_, connection_6__4__14_, 
        connection_6__4__13_, connection_6__4__12_, connection_6__4__11_, 
        connection_6__4__10_, connection_6__4__9_, connection_6__4__8_, 
        connection_6__4__7_, connection_6__4__6_, connection_6__4__5_, 
        connection_6__4__4_, connection_6__4__3_, connection_6__4__2_, 
        connection_6__4__1_, connection_6__4__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[91:90]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_45 second_half_stages_5__group_sec_half_0__switch_sec_half_3__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__7_, 
        connection_valid_5__3_}), .i_data_bus({connection_5__7__31_, 
        connection_5__7__30_, connection_5__7__29_, connection_5__7__28_, 
        connection_5__7__27_, connection_5__7__26_, connection_5__7__25_, 
        connection_5__7__24_, connection_5__7__23_, connection_5__7__22_, 
        connection_5__7__21_, connection_5__7__20_, connection_5__7__19_, 
        connection_5__7__18_, connection_5__7__17_, connection_5__7__16_, 
        connection_5__7__15_, connection_5__7__14_, connection_5__7__13_, 
        connection_5__7__12_, connection_5__7__11_, connection_5__7__10_, 
        connection_5__7__9_, connection_5__7__8_, connection_5__7__7_, 
        connection_5__7__6_, connection_5__7__5_, connection_5__7__4_, 
        connection_5__7__3_, connection_5__7__2_, connection_5__7__1_, 
        connection_5__7__0_, connection_5__3__31_, connection_5__3__30_, 
        connection_5__3__29_, connection_5__3__28_, connection_5__3__27_, 
        connection_5__3__26_, connection_5__3__25_, connection_5__3__24_, 
        connection_5__3__23_, connection_5__3__22_, connection_5__3__21_, 
        connection_5__3__20_, connection_5__3__19_, connection_5__3__18_, 
        connection_5__3__17_, connection_5__3__16_, connection_5__3__15_, 
        connection_5__3__14_, connection_5__3__13_, connection_5__3__12_, 
        connection_5__3__11_, connection_5__3__10_, connection_5__3__9_, 
        connection_5__3__8_, connection_5__3__7_, connection_5__3__6_, 
        connection_5__3__5_, connection_5__3__4_, connection_5__3__3_, 
        connection_5__3__2_, connection_5__3__1_, connection_5__3__0_}), 
        .o_valid({connection_valid_6__7_, connection_valid_6__6_}), 
        .o_data_bus({connection_6__7__31_, connection_6__7__30_, 
        connection_6__7__29_, connection_6__7__28_, connection_6__7__27_, 
        connection_6__7__26_, connection_6__7__25_, connection_6__7__24_, 
        connection_6__7__23_, connection_6__7__22_, connection_6__7__21_, 
        connection_6__7__20_, connection_6__7__19_, connection_6__7__18_, 
        connection_6__7__17_, connection_6__7__16_, connection_6__7__15_, 
        connection_6__7__14_, connection_6__7__13_, connection_6__7__12_, 
        connection_6__7__11_, connection_6__7__10_, connection_6__7__9_, 
        connection_6__7__8_, connection_6__7__7_, connection_6__7__6_, 
        connection_6__7__5_, connection_6__7__4_, connection_6__7__3_, 
        connection_6__7__2_, connection_6__7__1_, connection_6__7__0_, 
        connection_6__6__31_, connection_6__6__30_, connection_6__6__29_, 
        connection_6__6__28_, connection_6__6__27_, connection_6__6__26_, 
        connection_6__6__25_, connection_6__6__24_, connection_6__6__23_, 
        connection_6__6__22_, connection_6__6__21_, connection_6__6__20_, 
        connection_6__6__19_, connection_6__6__18_, connection_6__6__17_, 
        connection_6__6__16_, connection_6__6__15_, connection_6__6__14_, 
        connection_6__6__13_, connection_6__6__12_, connection_6__6__11_, 
        connection_6__6__10_, connection_6__6__9_, connection_6__6__8_, 
        connection_6__6__7_, connection_6__6__6_, connection_6__6__5_, 
        connection_6__6__4_, connection_6__6__3_, connection_6__6__2_, 
        connection_6__6__1_, connection_6__6__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[89:88]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_44 second_half_stages_5__group_sec_half_1__switch_sec_half_0__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__12_, 
        connection_valid_5__8_}), .i_data_bus({connection_5__12__31_, 
        connection_5__12__30_, connection_5__12__29_, connection_5__12__28_, 
        connection_5__12__27_, connection_5__12__26_, connection_5__12__25_, 
        connection_5__12__24_, connection_5__12__23_, connection_5__12__22_, 
        connection_5__12__21_, connection_5__12__20_, connection_5__12__19_, 
        connection_5__12__18_, connection_5__12__17_, connection_5__12__16_, 
        connection_5__12__15_, connection_5__12__14_, connection_5__12__13_, 
        connection_5__12__12_, connection_5__12__11_, connection_5__12__10_, 
        connection_5__12__9_, connection_5__12__8_, connection_5__12__7_, 
        connection_5__12__6_, connection_5__12__5_, connection_5__12__4_, 
        connection_5__12__3_, connection_5__12__2_, connection_5__12__1_, 
        connection_5__12__0_, connection_5__8__31_, connection_5__8__30_, 
        connection_5__8__29_, connection_5__8__28_, connection_5__8__27_, 
        connection_5__8__26_, connection_5__8__25_, connection_5__8__24_, 
        connection_5__8__23_, connection_5__8__22_, connection_5__8__21_, 
        connection_5__8__20_, connection_5__8__19_, connection_5__8__18_, 
        connection_5__8__17_, connection_5__8__16_, connection_5__8__15_, 
        connection_5__8__14_, connection_5__8__13_, connection_5__8__12_, 
        connection_5__8__11_, connection_5__8__10_, connection_5__8__9_, 
        connection_5__8__8_, connection_5__8__7_, connection_5__8__6_, 
        connection_5__8__5_, connection_5__8__4_, connection_5__8__3_, 
        connection_5__8__2_, connection_5__8__1_, connection_5__8__0_}), 
        .o_valid({connection_valid_6__9_, connection_valid_6__8_}), 
        .o_data_bus({connection_6__9__31_, connection_6__9__30_, 
        connection_6__9__29_, connection_6__9__28_, connection_6__9__27_, 
        connection_6__9__26_, connection_6__9__25_, connection_6__9__24_, 
        connection_6__9__23_, connection_6__9__22_, connection_6__9__21_, 
        connection_6__9__20_, connection_6__9__19_, connection_6__9__18_, 
        connection_6__9__17_, connection_6__9__16_, connection_6__9__15_, 
        connection_6__9__14_, connection_6__9__13_, connection_6__9__12_, 
        connection_6__9__11_, connection_6__9__10_, connection_6__9__9_, 
        connection_6__9__8_, connection_6__9__7_, connection_6__9__6_, 
        connection_6__9__5_, connection_6__9__4_, connection_6__9__3_, 
        connection_6__9__2_, connection_6__9__1_, connection_6__9__0_, 
        connection_6__8__31_, connection_6__8__30_, connection_6__8__29_, 
        connection_6__8__28_, connection_6__8__27_, connection_6__8__26_, 
        connection_6__8__25_, connection_6__8__24_, connection_6__8__23_, 
        connection_6__8__22_, connection_6__8__21_, connection_6__8__20_, 
        connection_6__8__19_, connection_6__8__18_, connection_6__8__17_, 
        connection_6__8__16_, connection_6__8__15_, connection_6__8__14_, 
        connection_6__8__13_, connection_6__8__12_, connection_6__8__11_, 
        connection_6__8__10_, connection_6__8__9_, connection_6__8__8_, 
        connection_6__8__7_, connection_6__8__6_, connection_6__8__5_, 
        connection_6__8__4_, connection_6__8__3_, connection_6__8__2_, 
        connection_6__8__1_, connection_6__8__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[87:86]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_43 second_half_stages_5__group_sec_half_1__switch_sec_half_1__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__13_, 
        connection_valid_5__9_}), .i_data_bus({connection_5__13__31_, 
        connection_5__13__30_, connection_5__13__29_, connection_5__13__28_, 
        connection_5__13__27_, connection_5__13__26_, connection_5__13__25_, 
        connection_5__13__24_, connection_5__13__23_, connection_5__13__22_, 
        connection_5__13__21_, connection_5__13__20_, connection_5__13__19_, 
        connection_5__13__18_, connection_5__13__17_, connection_5__13__16_, 
        connection_5__13__15_, connection_5__13__14_, connection_5__13__13_, 
        connection_5__13__12_, connection_5__13__11_, connection_5__13__10_, 
        connection_5__13__9_, connection_5__13__8_, connection_5__13__7_, 
        connection_5__13__6_, connection_5__13__5_, connection_5__13__4_, 
        connection_5__13__3_, connection_5__13__2_, connection_5__13__1_, 
        connection_5__13__0_, connection_5__9__31_, connection_5__9__30_, 
        connection_5__9__29_, connection_5__9__28_, connection_5__9__27_, 
        connection_5__9__26_, connection_5__9__25_, connection_5__9__24_, 
        connection_5__9__23_, connection_5__9__22_, connection_5__9__21_, 
        connection_5__9__20_, connection_5__9__19_, connection_5__9__18_, 
        connection_5__9__17_, connection_5__9__16_, connection_5__9__15_, 
        connection_5__9__14_, connection_5__9__13_, connection_5__9__12_, 
        connection_5__9__11_, connection_5__9__10_, connection_5__9__9_, 
        connection_5__9__8_, connection_5__9__7_, connection_5__9__6_, 
        connection_5__9__5_, connection_5__9__4_, connection_5__9__3_, 
        connection_5__9__2_, connection_5__9__1_, connection_5__9__0_}), 
        .o_valid({connection_valid_6__11_, connection_valid_6__10_}), 
        .o_data_bus({connection_6__11__31_, connection_6__11__30_, 
        connection_6__11__29_, connection_6__11__28_, connection_6__11__27_, 
        connection_6__11__26_, connection_6__11__25_, connection_6__11__24_, 
        connection_6__11__23_, connection_6__11__22_, connection_6__11__21_, 
        connection_6__11__20_, connection_6__11__19_, connection_6__11__18_, 
        connection_6__11__17_, connection_6__11__16_, connection_6__11__15_, 
        connection_6__11__14_, connection_6__11__13_, connection_6__11__12_, 
        connection_6__11__11_, connection_6__11__10_, connection_6__11__9_, 
        connection_6__11__8_, connection_6__11__7_, connection_6__11__6_, 
        connection_6__11__5_, connection_6__11__4_, connection_6__11__3_, 
        connection_6__11__2_, connection_6__11__1_, connection_6__11__0_, 
        connection_6__10__31_, connection_6__10__30_, connection_6__10__29_, 
        connection_6__10__28_, connection_6__10__27_, connection_6__10__26_, 
        connection_6__10__25_, connection_6__10__24_, connection_6__10__23_, 
        connection_6__10__22_, connection_6__10__21_, connection_6__10__20_, 
        connection_6__10__19_, connection_6__10__18_, connection_6__10__17_, 
        connection_6__10__16_, connection_6__10__15_, connection_6__10__14_, 
        connection_6__10__13_, connection_6__10__12_, connection_6__10__11_, 
        connection_6__10__10_, connection_6__10__9_, connection_6__10__8_, 
        connection_6__10__7_, connection_6__10__6_, connection_6__10__5_, 
        connection_6__10__4_, connection_6__10__3_, connection_6__10__2_, 
        connection_6__10__1_, connection_6__10__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[85:84]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_42 second_half_stages_5__group_sec_half_1__switch_sec_half_2__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__14_, 
        connection_valid_5__10_}), .i_data_bus({connection_5__14__31_, 
        connection_5__14__30_, connection_5__14__29_, connection_5__14__28_, 
        connection_5__14__27_, connection_5__14__26_, connection_5__14__25_, 
        connection_5__14__24_, connection_5__14__23_, connection_5__14__22_, 
        connection_5__14__21_, connection_5__14__20_, connection_5__14__19_, 
        connection_5__14__18_, connection_5__14__17_, connection_5__14__16_, 
        connection_5__14__15_, connection_5__14__14_, connection_5__14__13_, 
        connection_5__14__12_, connection_5__14__11_, connection_5__14__10_, 
        connection_5__14__9_, connection_5__14__8_, connection_5__14__7_, 
        connection_5__14__6_, connection_5__14__5_, connection_5__14__4_, 
        connection_5__14__3_, connection_5__14__2_, connection_5__14__1_, 
        connection_5__14__0_, connection_5__10__31_, connection_5__10__30_, 
        connection_5__10__29_, connection_5__10__28_, connection_5__10__27_, 
        connection_5__10__26_, connection_5__10__25_, connection_5__10__24_, 
        connection_5__10__23_, connection_5__10__22_, connection_5__10__21_, 
        connection_5__10__20_, connection_5__10__19_, connection_5__10__18_, 
        connection_5__10__17_, connection_5__10__16_, connection_5__10__15_, 
        connection_5__10__14_, connection_5__10__13_, connection_5__10__12_, 
        connection_5__10__11_, connection_5__10__10_, connection_5__10__9_, 
        connection_5__10__8_, connection_5__10__7_, connection_5__10__6_, 
        connection_5__10__5_, connection_5__10__4_, connection_5__10__3_, 
        connection_5__10__2_, connection_5__10__1_, connection_5__10__0_}), 
        .o_valid({connection_valid_6__13_, connection_valid_6__12_}), 
        .o_data_bus({connection_6__13__31_, connection_6__13__30_, 
        connection_6__13__29_, connection_6__13__28_, connection_6__13__27_, 
        connection_6__13__26_, connection_6__13__25_, connection_6__13__24_, 
        connection_6__13__23_, connection_6__13__22_, connection_6__13__21_, 
        connection_6__13__20_, connection_6__13__19_, connection_6__13__18_, 
        connection_6__13__17_, connection_6__13__16_, connection_6__13__15_, 
        connection_6__13__14_, connection_6__13__13_, connection_6__13__12_, 
        connection_6__13__11_, connection_6__13__10_, connection_6__13__9_, 
        connection_6__13__8_, connection_6__13__7_, connection_6__13__6_, 
        connection_6__13__5_, connection_6__13__4_, connection_6__13__3_, 
        connection_6__13__2_, connection_6__13__1_, connection_6__13__0_, 
        connection_6__12__31_, connection_6__12__30_, connection_6__12__29_, 
        connection_6__12__28_, connection_6__12__27_, connection_6__12__26_, 
        connection_6__12__25_, connection_6__12__24_, connection_6__12__23_, 
        connection_6__12__22_, connection_6__12__21_, connection_6__12__20_, 
        connection_6__12__19_, connection_6__12__18_, connection_6__12__17_, 
        connection_6__12__16_, connection_6__12__15_, connection_6__12__14_, 
        connection_6__12__13_, connection_6__12__12_, connection_6__12__11_, 
        connection_6__12__10_, connection_6__12__9_, connection_6__12__8_, 
        connection_6__12__7_, connection_6__12__6_, connection_6__12__5_, 
        connection_6__12__4_, connection_6__12__3_, connection_6__12__2_, 
        connection_6__12__1_, connection_6__12__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[83:82]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_41 second_half_stages_5__group_sec_half_1__switch_sec_half_3__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__15_, 
        connection_valid_5__11_}), .i_data_bus({connection_5__15__31_, 
        connection_5__15__30_, connection_5__15__29_, connection_5__15__28_, 
        connection_5__15__27_, connection_5__15__26_, connection_5__15__25_, 
        connection_5__15__24_, connection_5__15__23_, connection_5__15__22_, 
        connection_5__15__21_, connection_5__15__20_, connection_5__15__19_, 
        connection_5__15__18_, connection_5__15__17_, connection_5__15__16_, 
        connection_5__15__15_, connection_5__15__14_, connection_5__15__13_, 
        connection_5__15__12_, connection_5__15__11_, connection_5__15__10_, 
        connection_5__15__9_, connection_5__15__8_, connection_5__15__7_, 
        connection_5__15__6_, connection_5__15__5_, connection_5__15__4_, 
        connection_5__15__3_, connection_5__15__2_, connection_5__15__1_, 
        connection_5__15__0_, connection_5__11__31_, connection_5__11__30_, 
        connection_5__11__29_, connection_5__11__28_, connection_5__11__27_, 
        connection_5__11__26_, connection_5__11__25_, connection_5__11__24_, 
        connection_5__11__23_, connection_5__11__22_, connection_5__11__21_, 
        connection_5__11__20_, connection_5__11__19_, connection_5__11__18_, 
        connection_5__11__17_, connection_5__11__16_, connection_5__11__15_, 
        connection_5__11__14_, connection_5__11__13_, connection_5__11__12_, 
        connection_5__11__11_, connection_5__11__10_, connection_5__11__9_, 
        connection_5__11__8_, connection_5__11__7_, connection_5__11__6_, 
        connection_5__11__5_, connection_5__11__4_, connection_5__11__3_, 
        connection_5__11__2_, connection_5__11__1_, connection_5__11__0_}), 
        .o_valid({connection_valid_6__15_, connection_valid_6__14_}), 
        .o_data_bus({connection_6__15__31_, connection_6__15__30_, 
        connection_6__15__29_, connection_6__15__28_, connection_6__15__27_, 
        connection_6__15__26_, connection_6__15__25_, connection_6__15__24_, 
        connection_6__15__23_, connection_6__15__22_, connection_6__15__21_, 
        connection_6__15__20_, connection_6__15__19_, connection_6__15__18_, 
        connection_6__15__17_, connection_6__15__16_, connection_6__15__15_, 
        connection_6__15__14_, connection_6__15__13_, connection_6__15__12_, 
        connection_6__15__11_, connection_6__15__10_, connection_6__15__9_, 
        connection_6__15__8_, connection_6__15__7_, connection_6__15__6_, 
        connection_6__15__5_, connection_6__15__4_, connection_6__15__3_, 
        connection_6__15__2_, connection_6__15__1_, connection_6__15__0_, 
        connection_6__14__31_, connection_6__14__30_, connection_6__14__29_, 
        connection_6__14__28_, connection_6__14__27_, connection_6__14__26_, 
        connection_6__14__25_, connection_6__14__24_, connection_6__14__23_, 
        connection_6__14__22_, connection_6__14__21_, connection_6__14__20_, 
        connection_6__14__19_, connection_6__14__18_, connection_6__14__17_, 
        connection_6__14__16_, connection_6__14__15_, connection_6__14__14_, 
        connection_6__14__13_, connection_6__14__12_, connection_6__14__11_, 
        connection_6__14__10_, connection_6__14__9_, connection_6__14__8_, 
        connection_6__14__7_, connection_6__14__6_, connection_6__14__5_, 
        connection_6__14__4_, connection_6__14__3_, connection_6__14__2_, 
        connection_6__14__1_, connection_6__14__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[81:80]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_40 second_half_stages_5__group_sec_half_2__switch_sec_half_0__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__20_, 
        connection_valid_5__16_}), .i_data_bus({connection_5__20__31_, 
        connection_5__20__30_, connection_5__20__29_, connection_5__20__28_, 
        connection_5__20__27_, connection_5__20__26_, connection_5__20__25_, 
        connection_5__20__24_, connection_5__20__23_, connection_5__20__22_, 
        connection_5__20__21_, connection_5__20__20_, connection_5__20__19_, 
        connection_5__20__18_, connection_5__20__17_, connection_5__20__16_, 
        connection_5__20__15_, connection_5__20__14_, connection_5__20__13_, 
        connection_5__20__12_, connection_5__20__11_, connection_5__20__10_, 
        connection_5__20__9_, connection_5__20__8_, connection_5__20__7_, 
        connection_5__20__6_, connection_5__20__5_, connection_5__20__4_, 
        connection_5__20__3_, connection_5__20__2_, connection_5__20__1_, 
        connection_5__20__0_, connection_5__16__31_, connection_5__16__30_, 
        connection_5__16__29_, connection_5__16__28_, connection_5__16__27_, 
        connection_5__16__26_, connection_5__16__25_, connection_5__16__24_, 
        connection_5__16__23_, connection_5__16__22_, connection_5__16__21_, 
        connection_5__16__20_, connection_5__16__19_, connection_5__16__18_, 
        connection_5__16__17_, connection_5__16__16_, connection_5__16__15_, 
        connection_5__16__14_, connection_5__16__13_, connection_5__16__12_, 
        connection_5__16__11_, connection_5__16__10_, connection_5__16__9_, 
        connection_5__16__8_, connection_5__16__7_, connection_5__16__6_, 
        connection_5__16__5_, connection_5__16__4_, connection_5__16__3_, 
        connection_5__16__2_, connection_5__16__1_, connection_5__16__0_}), 
        .o_valid({connection_valid_6__17_, connection_valid_6__16_}), 
        .o_data_bus({connection_6__17__31_, connection_6__17__30_, 
        connection_6__17__29_, connection_6__17__28_, connection_6__17__27_, 
        connection_6__17__26_, connection_6__17__25_, connection_6__17__24_, 
        connection_6__17__23_, connection_6__17__22_, connection_6__17__21_, 
        connection_6__17__20_, connection_6__17__19_, connection_6__17__18_, 
        connection_6__17__17_, connection_6__17__16_, connection_6__17__15_, 
        connection_6__17__14_, connection_6__17__13_, connection_6__17__12_, 
        connection_6__17__11_, connection_6__17__10_, connection_6__17__9_, 
        connection_6__17__8_, connection_6__17__7_, connection_6__17__6_, 
        connection_6__17__5_, connection_6__17__4_, connection_6__17__3_, 
        connection_6__17__2_, connection_6__17__1_, connection_6__17__0_, 
        connection_6__16__31_, connection_6__16__30_, connection_6__16__29_, 
        connection_6__16__28_, connection_6__16__27_, connection_6__16__26_, 
        connection_6__16__25_, connection_6__16__24_, connection_6__16__23_, 
        connection_6__16__22_, connection_6__16__21_, connection_6__16__20_, 
        connection_6__16__19_, connection_6__16__18_, connection_6__16__17_, 
        connection_6__16__16_, connection_6__16__15_, connection_6__16__14_, 
        connection_6__16__13_, connection_6__16__12_, connection_6__16__11_, 
        connection_6__16__10_, connection_6__16__9_, connection_6__16__8_, 
        connection_6__16__7_, connection_6__16__6_, connection_6__16__5_, 
        connection_6__16__4_, connection_6__16__3_, connection_6__16__2_, 
        connection_6__16__1_, connection_6__16__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[79:78]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_39 second_half_stages_5__group_sec_half_2__switch_sec_half_1__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__21_, 
        connection_valid_5__17_}), .i_data_bus({connection_5__21__31_, 
        connection_5__21__30_, connection_5__21__29_, connection_5__21__28_, 
        connection_5__21__27_, connection_5__21__26_, connection_5__21__25_, 
        connection_5__21__24_, connection_5__21__23_, connection_5__21__22_, 
        connection_5__21__21_, connection_5__21__20_, connection_5__21__19_, 
        connection_5__21__18_, connection_5__21__17_, connection_5__21__16_, 
        connection_5__21__15_, connection_5__21__14_, connection_5__21__13_, 
        connection_5__21__12_, connection_5__21__11_, connection_5__21__10_, 
        connection_5__21__9_, connection_5__21__8_, connection_5__21__7_, 
        connection_5__21__6_, connection_5__21__5_, connection_5__21__4_, 
        connection_5__21__3_, connection_5__21__2_, connection_5__21__1_, 
        connection_5__21__0_, connection_5__17__31_, connection_5__17__30_, 
        connection_5__17__29_, connection_5__17__28_, connection_5__17__27_, 
        connection_5__17__26_, connection_5__17__25_, connection_5__17__24_, 
        connection_5__17__23_, connection_5__17__22_, connection_5__17__21_, 
        connection_5__17__20_, connection_5__17__19_, connection_5__17__18_, 
        connection_5__17__17_, connection_5__17__16_, connection_5__17__15_, 
        connection_5__17__14_, connection_5__17__13_, connection_5__17__12_, 
        connection_5__17__11_, connection_5__17__10_, connection_5__17__9_, 
        connection_5__17__8_, connection_5__17__7_, connection_5__17__6_, 
        connection_5__17__5_, connection_5__17__4_, connection_5__17__3_, 
        connection_5__17__2_, connection_5__17__1_, connection_5__17__0_}), 
        .o_valid({connection_valid_6__19_, connection_valid_6__18_}), 
        .o_data_bus({connection_6__19__31_, connection_6__19__30_, 
        connection_6__19__29_, connection_6__19__28_, connection_6__19__27_, 
        connection_6__19__26_, connection_6__19__25_, connection_6__19__24_, 
        connection_6__19__23_, connection_6__19__22_, connection_6__19__21_, 
        connection_6__19__20_, connection_6__19__19_, connection_6__19__18_, 
        connection_6__19__17_, connection_6__19__16_, connection_6__19__15_, 
        connection_6__19__14_, connection_6__19__13_, connection_6__19__12_, 
        connection_6__19__11_, connection_6__19__10_, connection_6__19__9_, 
        connection_6__19__8_, connection_6__19__7_, connection_6__19__6_, 
        connection_6__19__5_, connection_6__19__4_, connection_6__19__3_, 
        connection_6__19__2_, connection_6__19__1_, connection_6__19__0_, 
        connection_6__18__31_, connection_6__18__30_, connection_6__18__29_, 
        connection_6__18__28_, connection_6__18__27_, connection_6__18__26_, 
        connection_6__18__25_, connection_6__18__24_, connection_6__18__23_, 
        connection_6__18__22_, connection_6__18__21_, connection_6__18__20_, 
        connection_6__18__19_, connection_6__18__18_, connection_6__18__17_, 
        connection_6__18__16_, connection_6__18__15_, connection_6__18__14_, 
        connection_6__18__13_, connection_6__18__12_, connection_6__18__11_, 
        connection_6__18__10_, connection_6__18__9_, connection_6__18__8_, 
        connection_6__18__7_, connection_6__18__6_, connection_6__18__5_, 
        connection_6__18__4_, connection_6__18__3_, connection_6__18__2_, 
        connection_6__18__1_, connection_6__18__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[77:76]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_38 second_half_stages_5__group_sec_half_2__switch_sec_half_2__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__22_, 
        connection_valid_5__18_}), .i_data_bus({connection_5__22__31_, 
        connection_5__22__30_, connection_5__22__29_, connection_5__22__28_, 
        connection_5__22__27_, connection_5__22__26_, connection_5__22__25_, 
        connection_5__22__24_, connection_5__22__23_, connection_5__22__22_, 
        connection_5__22__21_, connection_5__22__20_, connection_5__22__19_, 
        connection_5__22__18_, connection_5__22__17_, connection_5__22__16_, 
        connection_5__22__15_, connection_5__22__14_, connection_5__22__13_, 
        connection_5__22__12_, connection_5__22__11_, connection_5__22__10_, 
        connection_5__22__9_, connection_5__22__8_, connection_5__22__7_, 
        connection_5__22__6_, connection_5__22__5_, connection_5__22__4_, 
        connection_5__22__3_, connection_5__22__2_, connection_5__22__1_, 
        connection_5__22__0_, connection_5__18__31_, connection_5__18__30_, 
        connection_5__18__29_, connection_5__18__28_, connection_5__18__27_, 
        connection_5__18__26_, connection_5__18__25_, connection_5__18__24_, 
        connection_5__18__23_, connection_5__18__22_, connection_5__18__21_, 
        connection_5__18__20_, connection_5__18__19_, connection_5__18__18_, 
        connection_5__18__17_, connection_5__18__16_, connection_5__18__15_, 
        connection_5__18__14_, connection_5__18__13_, connection_5__18__12_, 
        connection_5__18__11_, connection_5__18__10_, connection_5__18__9_, 
        connection_5__18__8_, connection_5__18__7_, connection_5__18__6_, 
        connection_5__18__5_, connection_5__18__4_, connection_5__18__3_, 
        connection_5__18__2_, connection_5__18__1_, connection_5__18__0_}), 
        .o_valid({connection_valid_6__21_, connection_valid_6__20_}), 
        .o_data_bus({connection_6__21__31_, connection_6__21__30_, 
        connection_6__21__29_, connection_6__21__28_, connection_6__21__27_, 
        connection_6__21__26_, connection_6__21__25_, connection_6__21__24_, 
        connection_6__21__23_, connection_6__21__22_, connection_6__21__21_, 
        connection_6__21__20_, connection_6__21__19_, connection_6__21__18_, 
        connection_6__21__17_, connection_6__21__16_, connection_6__21__15_, 
        connection_6__21__14_, connection_6__21__13_, connection_6__21__12_, 
        connection_6__21__11_, connection_6__21__10_, connection_6__21__9_, 
        connection_6__21__8_, connection_6__21__7_, connection_6__21__6_, 
        connection_6__21__5_, connection_6__21__4_, connection_6__21__3_, 
        connection_6__21__2_, connection_6__21__1_, connection_6__21__0_, 
        connection_6__20__31_, connection_6__20__30_, connection_6__20__29_, 
        connection_6__20__28_, connection_6__20__27_, connection_6__20__26_, 
        connection_6__20__25_, connection_6__20__24_, connection_6__20__23_, 
        connection_6__20__22_, connection_6__20__21_, connection_6__20__20_, 
        connection_6__20__19_, connection_6__20__18_, connection_6__20__17_, 
        connection_6__20__16_, connection_6__20__15_, connection_6__20__14_, 
        connection_6__20__13_, connection_6__20__12_, connection_6__20__11_, 
        connection_6__20__10_, connection_6__20__9_, connection_6__20__8_, 
        connection_6__20__7_, connection_6__20__6_, connection_6__20__5_, 
        connection_6__20__4_, connection_6__20__3_, connection_6__20__2_, 
        connection_6__20__1_, connection_6__20__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[75:74]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_37 second_half_stages_5__group_sec_half_2__switch_sec_half_3__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__23_, 
        connection_valid_5__19_}), .i_data_bus({connection_5__23__31_, 
        connection_5__23__30_, connection_5__23__29_, connection_5__23__28_, 
        connection_5__23__27_, connection_5__23__26_, connection_5__23__25_, 
        connection_5__23__24_, connection_5__23__23_, connection_5__23__22_, 
        connection_5__23__21_, connection_5__23__20_, connection_5__23__19_, 
        connection_5__23__18_, connection_5__23__17_, connection_5__23__16_, 
        connection_5__23__15_, connection_5__23__14_, connection_5__23__13_, 
        connection_5__23__12_, connection_5__23__11_, connection_5__23__10_, 
        connection_5__23__9_, connection_5__23__8_, connection_5__23__7_, 
        connection_5__23__6_, connection_5__23__5_, connection_5__23__4_, 
        connection_5__23__3_, connection_5__23__2_, connection_5__23__1_, 
        connection_5__23__0_, connection_5__19__31_, connection_5__19__30_, 
        connection_5__19__29_, connection_5__19__28_, connection_5__19__27_, 
        connection_5__19__26_, connection_5__19__25_, connection_5__19__24_, 
        connection_5__19__23_, connection_5__19__22_, connection_5__19__21_, 
        connection_5__19__20_, connection_5__19__19_, connection_5__19__18_, 
        connection_5__19__17_, connection_5__19__16_, connection_5__19__15_, 
        connection_5__19__14_, connection_5__19__13_, connection_5__19__12_, 
        connection_5__19__11_, connection_5__19__10_, connection_5__19__9_, 
        connection_5__19__8_, connection_5__19__7_, connection_5__19__6_, 
        connection_5__19__5_, connection_5__19__4_, connection_5__19__3_, 
        connection_5__19__2_, connection_5__19__1_, connection_5__19__0_}), 
        .o_valid({connection_valid_6__23_, connection_valid_6__22_}), 
        .o_data_bus({connection_6__23__31_, connection_6__23__30_, 
        connection_6__23__29_, connection_6__23__28_, connection_6__23__27_, 
        connection_6__23__26_, connection_6__23__25_, connection_6__23__24_, 
        connection_6__23__23_, connection_6__23__22_, connection_6__23__21_, 
        connection_6__23__20_, connection_6__23__19_, connection_6__23__18_, 
        connection_6__23__17_, connection_6__23__16_, connection_6__23__15_, 
        connection_6__23__14_, connection_6__23__13_, connection_6__23__12_, 
        connection_6__23__11_, connection_6__23__10_, connection_6__23__9_, 
        connection_6__23__8_, connection_6__23__7_, connection_6__23__6_, 
        connection_6__23__5_, connection_6__23__4_, connection_6__23__3_, 
        connection_6__23__2_, connection_6__23__1_, connection_6__23__0_, 
        connection_6__22__31_, connection_6__22__30_, connection_6__22__29_, 
        connection_6__22__28_, connection_6__22__27_, connection_6__22__26_, 
        connection_6__22__25_, connection_6__22__24_, connection_6__22__23_, 
        connection_6__22__22_, connection_6__22__21_, connection_6__22__20_, 
        connection_6__22__19_, connection_6__22__18_, connection_6__22__17_, 
        connection_6__22__16_, connection_6__22__15_, connection_6__22__14_, 
        connection_6__22__13_, connection_6__22__12_, connection_6__22__11_, 
        connection_6__22__10_, connection_6__22__9_, connection_6__22__8_, 
        connection_6__22__7_, connection_6__22__6_, connection_6__22__5_, 
        connection_6__22__4_, connection_6__22__3_, connection_6__22__2_, 
        connection_6__22__1_, connection_6__22__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[73:72]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_36 second_half_stages_5__group_sec_half_3__switch_sec_half_0__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__28_, 
        connection_valid_5__24_}), .i_data_bus({connection_5__28__31_, 
        connection_5__28__30_, connection_5__28__29_, connection_5__28__28_, 
        connection_5__28__27_, connection_5__28__26_, connection_5__28__25_, 
        connection_5__28__24_, connection_5__28__23_, connection_5__28__22_, 
        connection_5__28__21_, connection_5__28__20_, connection_5__28__19_, 
        connection_5__28__18_, connection_5__28__17_, connection_5__28__16_, 
        connection_5__28__15_, connection_5__28__14_, connection_5__28__13_, 
        connection_5__28__12_, connection_5__28__11_, connection_5__28__10_, 
        connection_5__28__9_, connection_5__28__8_, connection_5__28__7_, 
        connection_5__28__6_, connection_5__28__5_, connection_5__28__4_, 
        connection_5__28__3_, connection_5__28__2_, connection_5__28__1_, 
        connection_5__28__0_, connection_5__24__31_, connection_5__24__30_, 
        connection_5__24__29_, connection_5__24__28_, connection_5__24__27_, 
        connection_5__24__26_, connection_5__24__25_, connection_5__24__24_, 
        connection_5__24__23_, connection_5__24__22_, connection_5__24__21_, 
        connection_5__24__20_, connection_5__24__19_, connection_5__24__18_, 
        connection_5__24__17_, connection_5__24__16_, connection_5__24__15_, 
        connection_5__24__14_, connection_5__24__13_, connection_5__24__12_, 
        connection_5__24__11_, connection_5__24__10_, connection_5__24__9_, 
        connection_5__24__8_, connection_5__24__7_, connection_5__24__6_, 
        connection_5__24__5_, connection_5__24__4_, connection_5__24__3_, 
        connection_5__24__2_, connection_5__24__1_, connection_5__24__0_}), 
        .o_valid({connection_valid_6__25_, connection_valid_6__24_}), 
        .o_data_bus({connection_6__25__31_, connection_6__25__30_, 
        connection_6__25__29_, connection_6__25__28_, connection_6__25__27_, 
        connection_6__25__26_, connection_6__25__25_, connection_6__25__24_, 
        connection_6__25__23_, connection_6__25__22_, connection_6__25__21_, 
        connection_6__25__20_, connection_6__25__19_, connection_6__25__18_, 
        connection_6__25__17_, connection_6__25__16_, connection_6__25__15_, 
        connection_6__25__14_, connection_6__25__13_, connection_6__25__12_, 
        connection_6__25__11_, connection_6__25__10_, connection_6__25__9_, 
        connection_6__25__8_, connection_6__25__7_, connection_6__25__6_, 
        connection_6__25__5_, connection_6__25__4_, connection_6__25__3_, 
        connection_6__25__2_, connection_6__25__1_, connection_6__25__0_, 
        connection_6__24__31_, connection_6__24__30_, connection_6__24__29_, 
        connection_6__24__28_, connection_6__24__27_, connection_6__24__26_, 
        connection_6__24__25_, connection_6__24__24_, connection_6__24__23_, 
        connection_6__24__22_, connection_6__24__21_, connection_6__24__20_, 
        connection_6__24__19_, connection_6__24__18_, connection_6__24__17_, 
        connection_6__24__16_, connection_6__24__15_, connection_6__24__14_, 
        connection_6__24__13_, connection_6__24__12_, connection_6__24__11_, 
        connection_6__24__10_, connection_6__24__9_, connection_6__24__8_, 
        connection_6__24__7_, connection_6__24__6_, connection_6__24__5_, 
        connection_6__24__4_, connection_6__24__3_, connection_6__24__2_, 
        connection_6__24__1_, connection_6__24__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[71:70]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_35 second_half_stages_5__group_sec_half_3__switch_sec_half_1__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__29_, 
        connection_valid_5__25_}), .i_data_bus({connection_5__29__31_, 
        connection_5__29__30_, connection_5__29__29_, connection_5__29__28_, 
        connection_5__29__27_, connection_5__29__26_, connection_5__29__25_, 
        connection_5__29__24_, connection_5__29__23_, connection_5__29__22_, 
        connection_5__29__21_, connection_5__29__20_, connection_5__29__19_, 
        connection_5__29__18_, connection_5__29__17_, connection_5__29__16_, 
        connection_5__29__15_, connection_5__29__14_, connection_5__29__13_, 
        connection_5__29__12_, connection_5__29__11_, connection_5__29__10_, 
        connection_5__29__9_, connection_5__29__8_, connection_5__29__7_, 
        connection_5__29__6_, connection_5__29__5_, connection_5__29__4_, 
        connection_5__29__3_, connection_5__29__2_, connection_5__29__1_, 
        connection_5__29__0_, connection_5__25__31_, connection_5__25__30_, 
        connection_5__25__29_, connection_5__25__28_, connection_5__25__27_, 
        connection_5__25__26_, connection_5__25__25_, connection_5__25__24_, 
        connection_5__25__23_, connection_5__25__22_, connection_5__25__21_, 
        connection_5__25__20_, connection_5__25__19_, connection_5__25__18_, 
        connection_5__25__17_, connection_5__25__16_, connection_5__25__15_, 
        connection_5__25__14_, connection_5__25__13_, connection_5__25__12_, 
        connection_5__25__11_, connection_5__25__10_, connection_5__25__9_, 
        connection_5__25__8_, connection_5__25__7_, connection_5__25__6_, 
        connection_5__25__5_, connection_5__25__4_, connection_5__25__3_, 
        connection_5__25__2_, connection_5__25__1_, connection_5__25__0_}), 
        .o_valid({connection_valid_6__27_, connection_valid_6__26_}), 
        .o_data_bus({connection_6__27__31_, connection_6__27__30_, 
        connection_6__27__29_, connection_6__27__28_, connection_6__27__27_, 
        connection_6__27__26_, connection_6__27__25_, connection_6__27__24_, 
        connection_6__27__23_, connection_6__27__22_, connection_6__27__21_, 
        connection_6__27__20_, connection_6__27__19_, connection_6__27__18_, 
        connection_6__27__17_, connection_6__27__16_, connection_6__27__15_, 
        connection_6__27__14_, connection_6__27__13_, connection_6__27__12_, 
        connection_6__27__11_, connection_6__27__10_, connection_6__27__9_, 
        connection_6__27__8_, connection_6__27__7_, connection_6__27__6_, 
        connection_6__27__5_, connection_6__27__4_, connection_6__27__3_, 
        connection_6__27__2_, connection_6__27__1_, connection_6__27__0_, 
        connection_6__26__31_, connection_6__26__30_, connection_6__26__29_, 
        connection_6__26__28_, connection_6__26__27_, connection_6__26__26_, 
        connection_6__26__25_, connection_6__26__24_, connection_6__26__23_, 
        connection_6__26__22_, connection_6__26__21_, connection_6__26__20_, 
        connection_6__26__19_, connection_6__26__18_, connection_6__26__17_, 
        connection_6__26__16_, connection_6__26__15_, connection_6__26__14_, 
        connection_6__26__13_, connection_6__26__12_, connection_6__26__11_, 
        connection_6__26__10_, connection_6__26__9_, connection_6__26__8_, 
        connection_6__26__7_, connection_6__26__6_, connection_6__26__5_, 
        connection_6__26__4_, connection_6__26__3_, connection_6__26__2_, 
        connection_6__26__1_, connection_6__26__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[69:68]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_34 second_half_stages_5__group_sec_half_3__switch_sec_half_2__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__30_, 
        connection_valid_5__26_}), .i_data_bus({connection_5__30__31_, 
        connection_5__30__30_, connection_5__30__29_, connection_5__30__28_, 
        connection_5__30__27_, connection_5__30__26_, connection_5__30__25_, 
        connection_5__30__24_, connection_5__30__23_, connection_5__30__22_, 
        connection_5__30__21_, connection_5__30__20_, connection_5__30__19_, 
        connection_5__30__18_, connection_5__30__17_, connection_5__30__16_, 
        connection_5__30__15_, connection_5__30__14_, connection_5__30__13_, 
        connection_5__30__12_, connection_5__30__11_, connection_5__30__10_, 
        connection_5__30__9_, connection_5__30__8_, connection_5__30__7_, 
        connection_5__30__6_, connection_5__30__5_, connection_5__30__4_, 
        connection_5__30__3_, connection_5__30__2_, connection_5__30__1_, 
        connection_5__30__0_, connection_5__26__31_, connection_5__26__30_, 
        connection_5__26__29_, connection_5__26__28_, connection_5__26__27_, 
        connection_5__26__26_, connection_5__26__25_, connection_5__26__24_, 
        connection_5__26__23_, connection_5__26__22_, connection_5__26__21_, 
        connection_5__26__20_, connection_5__26__19_, connection_5__26__18_, 
        connection_5__26__17_, connection_5__26__16_, connection_5__26__15_, 
        connection_5__26__14_, connection_5__26__13_, connection_5__26__12_, 
        connection_5__26__11_, connection_5__26__10_, connection_5__26__9_, 
        connection_5__26__8_, connection_5__26__7_, connection_5__26__6_, 
        connection_5__26__5_, connection_5__26__4_, connection_5__26__3_, 
        connection_5__26__2_, connection_5__26__1_, connection_5__26__0_}), 
        .o_valid({connection_valid_6__29_, connection_valid_6__28_}), 
        .o_data_bus({connection_6__29__31_, connection_6__29__30_, 
        connection_6__29__29_, connection_6__29__28_, connection_6__29__27_, 
        connection_6__29__26_, connection_6__29__25_, connection_6__29__24_, 
        connection_6__29__23_, connection_6__29__22_, connection_6__29__21_, 
        connection_6__29__20_, connection_6__29__19_, connection_6__29__18_, 
        connection_6__29__17_, connection_6__29__16_, connection_6__29__15_, 
        connection_6__29__14_, connection_6__29__13_, connection_6__29__12_, 
        connection_6__29__11_, connection_6__29__10_, connection_6__29__9_, 
        connection_6__29__8_, connection_6__29__7_, connection_6__29__6_, 
        connection_6__29__5_, connection_6__29__4_, connection_6__29__3_, 
        connection_6__29__2_, connection_6__29__1_, connection_6__29__0_, 
        connection_6__28__31_, connection_6__28__30_, connection_6__28__29_, 
        connection_6__28__28_, connection_6__28__27_, connection_6__28__26_, 
        connection_6__28__25_, connection_6__28__24_, connection_6__28__23_, 
        connection_6__28__22_, connection_6__28__21_, connection_6__28__20_, 
        connection_6__28__19_, connection_6__28__18_, connection_6__28__17_, 
        connection_6__28__16_, connection_6__28__15_, connection_6__28__14_, 
        connection_6__28__13_, connection_6__28__12_, connection_6__28__11_, 
        connection_6__28__10_, connection_6__28__9_, connection_6__28__8_, 
        connection_6__28__7_, connection_6__28__6_, connection_6__28__5_, 
        connection_6__28__4_, connection_6__28__3_, connection_6__28__2_, 
        connection_6__28__1_, connection_6__28__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[67:66]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_33 second_half_stages_5__group_sec_half_3__switch_sec_half_3__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__31_, 
        connection_valid_5__27_}), .i_data_bus({connection_5__31__31_, 
        connection_5__31__30_, connection_5__31__29_, connection_5__31__28_, 
        connection_5__31__27_, connection_5__31__26_, connection_5__31__25_, 
        connection_5__31__24_, connection_5__31__23_, connection_5__31__22_, 
        connection_5__31__21_, connection_5__31__20_, connection_5__31__19_, 
        connection_5__31__18_, connection_5__31__17_, connection_5__31__16_, 
        connection_5__31__15_, connection_5__31__14_, connection_5__31__13_, 
        connection_5__31__12_, connection_5__31__11_, connection_5__31__10_, 
        connection_5__31__9_, connection_5__31__8_, connection_5__31__7_, 
        connection_5__31__6_, connection_5__31__5_, connection_5__31__4_, 
        connection_5__31__3_, connection_5__31__2_, connection_5__31__1_, 
        connection_5__31__0_, connection_5__27__31_, connection_5__27__30_, 
        connection_5__27__29_, connection_5__27__28_, connection_5__27__27_, 
        connection_5__27__26_, connection_5__27__25_, connection_5__27__24_, 
        connection_5__27__23_, connection_5__27__22_, connection_5__27__21_, 
        connection_5__27__20_, connection_5__27__19_, connection_5__27__18_, 
        connection_5__27__17_, connection_5__27__16_, connection_5__27__15_, 
        connection_5__27__14_, connection_5__27__13_, connection_5__27__12_, 
        connection_5__27__11_, connection_5__27__10_, connection_5__27__9_, 
        connection_5__27__8_, connection_5__27__7_, connection_5__27__6_, 
        connection_5__27__5_, connection_5__27__4_, connection_5__27__3_, 
        connection_5__27__2_, connection_5__27__1_, connection_5__27__0_}), 
        .o_valid({connection_valid_6__31_, connection_valid_6__30_}), 
        .o_data_bus({connection_6__31__31_, connection_6__31__30_, 
        connection_6__31__29_, connection_6__31__28_, connection_6__31__27_, 
        connection_6__31__26_, connection_6__31__25_, connection_6__31__24_, 
        connection_6__31__23_, connection_6__31__22_, connection_6__31__21_, 
        connection_6__31__20_, connection_6__31__19_, connection_6__31__18_, 
        connection_6__31__17_, connection_6__31__16_, connection_6__31__15_, 
        connection_6__31__14_, connection_6__31__13_, connection_6__31__12_, 
        connection_6__31__11_, connection_6__31__10_, connection_6__31__9_, 
        connection_6__31__8_, connection_6__31__7_, connection_6__31__6_, 
        connection_6__31__5_, connection_6__31__4_, connection_6__31__3_, 
        connection_6__31__2_, connection_6__31__1_, connection_6__31__0_, 
        connection_6__30__31_, connection_6__30__30_, connection_6__30__29_, 
        connection_6__30__28_, connection_6__30__27_, connection_6__30__26_, 
        connection_6__30__25_, connection_6__30__24_, connection_6__30__23_, 
        connection_6__30__22_, connection_6__30__21_, connection_6__30__20_, 
        connection_6__30__19_, connection_6__30__18_, connection_6__30__17_, 
        connection_6__30__16_, connection_6__30__15_, connection_6__30__14_, 
        connection_6__30__13_, connection_6__30__12_, connection_6__30__11_, 
        connection_6__30__10_, connection_6__30__9_, connection_6__30__8_, 
        connection_6__30__7_, connection_6__30__6_, connection_6__30__5_, 
        connection_6__30__4_, connection_6__30__3_, connection_6__30__2_, 
        connection_6__30__1_, connection_6__30__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[65:64]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_32 second_half_stages_6__group_sec_half_0__switch_sec_half_0__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_6__8_, 
        connection_valid_6__0_}), .i_data_bus({connection_6__8__31_, 
        connection_6__8__30_, connection_6__8__29_, connection_6__8__28_, 
        connection_6__8__27_, connection_6__8__26_, connection_6__8__25_, 
        connection_6__8__24_, connection_6__8__23_, connection_6__8__22_, 
        connection_6__8__21_, connection_6__8__20_, connection_6__8__19_, 
        connection_6__8__18_, connection_6__8__17_, connection_6__8__16_, 
        connection_6__8__15_, connection_6__8__14_, connection_6__8__13_, 
        connection_6__8__12_, connection_6__8__11_, connection_6__8__10_, 
        connection_6__8__9_, connection_6__8__8_, connection_6__8__7_, 
        connection_6__8__6_, connection_6__8__5_, connection_6__8__4_, 
        connection_6__8__3_, connection_6__8__2_, connection_6__8__1_, 
        connection_6__8__0_, connection_6__0__31_, connection_6__0__30_, 
        connection_6__0__29_, connection_6__0__28_, connection_6__0__27_, 
        connection_6__0__26_, connection_6__0__25_, connection_6__0__24_, 
        connection_6__0__23_, connection_6__0__22_, connection_6__0__21_, 
        connection_6__0__20_, connection_6__0__19_, connection_6__0__18_, 
        connection_6__0__17_, connection_6__0__16_, connection_6__0__15_, 
        connection_6__0__14_, connection_6__0__13_, connection_6__0__12_, 
        connection_6__0__11_, connection_6__0__10_, connection_6__0__9_, 
        connection_6__0__8_, connection_6__0__7_, connection_6__0__6_, 
        connection_6__0__5_, connection_6__0__4_, connection_6__0__3_, 
        connection_6__0__2_, connection_6__0__1_, connection_6__0__0_}), 
        .o_valid({connection_valid_7__1_, connection_valid_7__0_}), 
        .o_data_bus({connection_7__1__31_, connection_7__1__30_, 
        connection_7__1__29_, connection_7__1__28_, connection_7__1__27_, 
        connection_7__1__26_, connection_7__1__25_, connection_7__1__24_, 
        connection_7__1__23_, connection_7__1__22_, connection_7__1__21_, 
        connection_7__1__20_, connection_7__1__19_, connection_7__1__18_, 
        connection_7__1__17_, connection_7__1__16_, connection_7__1__15_, 
        connection_7__1__14_, connection_7__1__13_, connection_7__1__12_, 
        connection_7__1__11_, connection_7__1__10_, connection_7__1__9_, 
        connection_7__1__8_, connection_7__1__7_, connection_7__1__6_, 
        connection_7__1__5_, connection_7__1__4_, connection_7__1__3_, 
        connection_7__1__2_, connection_7__1__1_, connection_7__1__0_, 
        connection_7__0__31_, connection_7__0__30_, connection_7__0__29_, 
        connection_7__0__28_, connection_7__0__27_, connection_7__0__26_, 
        connection_7__0__25_, connection_7__0__24_, connection_7__0__23_, 
        connection_7__0__22_, connection_7__0__21_, connection_7__0__20_, 
        connection_7__0__19_, connection_7__0__18_, connection_7__0__17_, 
        connection_7__0__16_, connection_7__0__15_, connection_7__0__14_, 
        connection_7__0__13_, connection_7__0__12_, connection_7__0__11_, 
        connection_7__0__10_, connection_7__0__9_, connection_7__0__8_, 
        connection_7__0__7_, connection_7__0__6_, connection_7__0__5_, 
        connection_7__0__4_, connection_7__0__3_, connection_7__0__2_, 
        connection_7__0__1_, connection_7__0__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[63:62]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_31 second_half_stages_6__group_sec_half_0__switch_sec_half_1__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_6__9_, 
        connection_valid_6__1_}), .i_data_bus({connection_6__9__31_, 
        connection_6__9__30_, connection_6__9__29_, connection_6__9__28_, 
        connection_6__9__27_, connection_6__9__26_, connection_6__9__25_, 
        connection_6__9__24_, connection_6__9__23_, connection_6__9__22_, 
        connection_6__9__21_, connection_6__9__20_, connection_6__9__19_, 
        connection_6__9__18_, connection_6__9__17_, connection_6__9__16_, 
        connection_6__9__15_, connection_6__9__14_, connection_6__9__13_, 
        connection_6__9__12_, connection_6__9__11_, connection_6__9__10_, 
        connection_6__9__9_, connection_6__9__8_, connection_6__9__7_, 
        connection_6__9__6_, connection_6__9__5_, connection_6__9__4_, 
        connection_6__9__3_, connection_6__9__2_, connection_6__9__1_, 
        connection_6__9__0_, connection_6__1__31_, connection_6__1__30_, 
        connection_6__1__29_, connection_6__1__28_, connection_6__1__27_, 
        connection_6__1__26_, connection_6__1__25_, connection_6__1__24_, 
        connection_6__1__23_, connection_6__1__22_, connection_6__1__21_, 
        connection_6__1__20_, connection_6__1__19_, connection_6__1__18_, 
        connection_6__1__17_, connection_6__1__16_, connection_6__1__15_, 
        connection_6__1__14_, connection_6__1__13_, connection_6__1__12_, 
        connection_6__1__11_, connection_6__1__10_, connection_6__1__9_, 
        connection_6__1__8_, connection_6__1__7_, connection_6__1__6_, 
        connection_6__1__5_, connection_6__1__4_, connection_6__1__3_, 
        connection_6__1__2_, connection_6__1__1_, connection_6__1__0_}), 
        .o_valid({connection_valid_7__3_, connection_valid_7__2_}), 
        .o_data_bus({connection_7__3__31_, connection_7__3__30_, 
        connection_7__3__29_, connection_7__3__28_, connection_7__3__27_, 
        connection_7__3__26_, connection_7__3__25_, connection_7__3__24_, 
        connection_7__3__23_, connection_7__3__22_, connection_7__3__21_, 
        connection_7__3__20_, connection_7__3__19_, connection_7__3__18_, 
        connection_7__3__17_, connection_7__3__16_, connection_7__3__15_, 
        connection_7__3__14_, connection_7__3__13_, connection_7__3__12_, 
        connection_7__3__11_, connection_7__3__10_, connection_7__3__9_, 
        connection_7__3__8_, connection_7__3__7_, connection_7__3__6_, 
        connection_7__3__5_, connection_7__3__4_, connection_7__3__3_, 
        connection_7__3__2_, connection_7__3__1_, connection_7__3__0_, 
        connection_7__2__31_, connection_7__2__30_, connection_7__2__29_, 
        connection_7__2__28_, connection_7__2__27_, connection_7__2__26_, 
        connection_7__2__25_, connection_7__2__24_, connection_7__2__23_, 
        connection_7__2__22_, connection_7__2__21_, connection_7__2__20_, 
        connection_7__2__19_, connection_7__2__18_, connection_7__2__17_, 
        connection_7__2__16_, connection_7__2__15_, connection_7__2__14_, 
        connection_7__2__13_, connection_7__2__12_, connection_7__2__11_, 
        connection_7__2__10_, connection_7__2__9_, connection_7__2__8_, 
        connection_7__2__7_, connection_7__2__6_, connection_7__2__5_, 
        connection_7__2__4_, connection_7__2__3_, connection_7__2__2_, 
        connection_7__2__1_, connection_7__2__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[61:60]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_30 second_half_stages_6__group_sec_half_0__switch_sec_half_2__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_6__10_, 
        connection_valid_6__2_}), .i_data_bus({connection_6__10__31_, 
        connection_6__10__30_, connection_6__10__29_, connection_6__10__28_, 
        connection_6__10__27_, connection_6__10__26_, connection_6__10__25_, 
        connection_6__10__24_, connection_6__10__23_, connection_6__10__22_, 
        connection_6__10__21_, connection_6__10__20_, connection_6__10__19_, 
        connection_6__10__18_, connection_6__10__17_, connection_6__10__16_, 
        connection_6__10__15_, connection_6__10__14_, connection_6__10__13_, 
        connection_6__10__12_, connection_6__10__11_, connection_6__10__10_, 
        connection_6__10__9_, connection_6__10__8_, connection_6__10__7_, 
        connection_6__10__6_, connection_6__10__5_, connection_6__10__4_, 
        connection_6__10__3_, connection_6__10__2_, connection_6__10__1_, 
        connection_6__10__0_, connection_6__2__31_, connection_6__2__30_, 
        connection_6__2__29_, connection_6__2__28_, connection_6__2__27_, 
        connection_6__2__26_, connection_6__2__25_, connection_6__2__24_, 
        connection_6__2__23_, connection_6__2__22_, connection_6__2__21_, 
        connection_6__2__20_, connection_6__2__19_, connection_6__2__18_, 
        connection_6__2__17_, connection_6__2__16_, connection_6__2__15_, 
        connection_6__2__14_, connection_6__2__13_, connection_6__2__12_, 
        connection_6__2__11_, connection_6__2__10_, connection_6__2__9_, 
        connection_6__2__8_, connection_6__2__7_, connection_6__2__6_, 
        connection_6__2__5_, connection_6__2__4_, connection_6__2__3_, 
        connection_6__2__2_, connection_6__2__1_, connection_6__2__0_}), 
        .o_valid({connection_valid_7__5_, connection_valid_7__4_}), 
        .o_data_bus({connection_7__5__31_, connection_7__5__30_, 
        connection_7__5__29_, connection_7__5__28_, connection_7__5__27_, 
        connection_7__5__26_, connection_7__5__25_, connection_7__5__24_, 
        connection_7__5__23_, connection_7__5__22_, connection_7__5__21_, 
        connection_7__5__20_, connection_7__5__19_, connection_7__5__18_, 
        connection_7__5__17_, connection_7__5__16_, connection_7__5__15_, 
        connection_7__5__14_, connection_7__5__13_, connection_7__5__12_, 
        connection_7__5__11_, connection_7__5__10_, connection_7__5__9_, 
        connection_7__5__8_, connection_7__5__7_, connection_7__5__6_, 
        connection_7__5__5_, connection_7__5__4_, connection_7__5__3_, 
        connection_7__5__2_, connection_7__5__1_, connection_7__5__0_, 
        connection_7__4__31_, connection_7__4__30_, connection_7__4__29_, 
        connection_7__4__28_, connection_7__4__27_, connection_7__4__26_, 
        connection_7__4__25_, connection_7__4__24_, connection_7__4__23_, 
        connection_7__4__22_, connection_7__4__21_, connection_7__4__20_, 
        connection_7__4__19_, connection_7__4__18_, connection_7__4__17_, 
        connection_7__4__16_, connection_7__4__15_, connection_7__4__14_, 
        connection_7__4__13_, connection_7__4__12_, connection_7__4__11_, 
        connection_7__4__10_, connection_7__4__9_, connection_7__4__8_, 
        connection_7__4__7_, connection_7__4__6_, connection_7__4__5_, 
        connection_7__4__4_, connection_7__4__3_, connection_7__4__2_, 
        connection_7__4__1_, connection_7__4__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[59:58]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_29 second_half_stages_6__group_sec_half_0__switch_sec_half_3__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_6__11_, 
        connection_valid_6__3_}), .i_data_bus({connection_6__11__31_, 
        connection_6__11__30_, connection_6__11__29_, connection_6__11__28_, 
        connection_6__11__27_, connection_6__11__26_, connection_6__11__25_, 
        connection_6__11__24_, connection_6__11__23_, connection_6__11__22_, 
        connection_6__11__21_, connection_6__11__20_, connection_6__11__19_, 
        connection_6__11__18_, connection_6__11__17_, connection_6__11__16_, 
        connection_6__11__15_, connection_6__11__14_, connection_6__11__13_, 
        connection_6__11__12_, connection_6__11__11_, connection_6__11__10_, 
        connection_6__11__9_, connection_6__11__8_, connection_6__11__7_, 
        connection_6__11__6_, connection_6__11__5_, connection_6__11__4_, 
        connection_6__11__3_, connection_6__11__2_, connection_6__11__1_, 
        connection_6__11__0_, connection_6__3__31_, connection_6__3__30_, 
        connection_6__3__29_, connection_6__3__28_, connection_6__3__27_, 
        connection_6__3__26_, connection_6__3__25_, connection_6__3__24_, 
        connection_6__3__23_, connection_6__3__22_, connection_6__3__21_, 
        connection_6__3__20_, connection_6__3__19_, connection_6__3__18_, 
        connection_6__3__17_, connection_6__3__16_, connection_6__3__15_, 
        connection_6__3__14_, connection_6__3__13_, connection_6__3__12_, 
        connection_6__3__11_, connection_6__3__10_, connection_6__3__9_, 
        connection_6__3__8_, connection_6__3__7_, connection_6__3__6_, 
        connection_6__3__5_, connection_6__3__4_, connection_6__3__3_, 
        connection_6__3__2_, connection_6__3__1_, connection_6__3__0_}), 
        .o_valid({connection_valid_7__7_, connection_valid_7__6_}), 
        .o_data_bus({connection_7__7__31_, connection_7__7__30_, 
        connection_7__7__29_, connection_7__7__28_, connection_7__7__27_, 
        connection_7__7__26_, connection_7__7__25_, connection_7__7__24_, 
        connection_7__7__23_, connection_7__7__22_, connection_7__7__21_, 
        connection_7__7__20_, connection_7__7__19_, connection_7__7__18_, 
        connection_7__7__17_, connection_7__7__16_, connection_7__7__15_, 
        connection_7__7__14_, connection_7__7__13_, connection_7__7__12_, 
        connection_7__7__11_, connection_7__7__10_, connection_7__7__9_, 
        connection_7__7__8_, connection_7__7__7_, connection_7__7__6_, 
        connection_7__7__5_, connection_7__7__4_, connection_7__7__3_, 
        connection_7__7__2_, connection_7__7__1_, connection_7__7__0_, 
        connection_7__6__31_, connection_7__6__30_, connection_7__6__29_, 
        connection_7__6__28_, connection_7__6__27_, connection_7__6__26_, 
        connection_7__6__25_, connection_7__6__24_, connection_7__6__23_, 
        connection_7__6__22_, connection_7__6__21_, connection_7__6__20_, 
        connection_7__6__19_, connection_7__6__18_, connection_7__6__17_, 
        connection_7__6__16_, connection_7__6__15_, connection_7__6__14_, 
        connection_7__6__13_, connection_7__6__12_, connection_7__6__11_, 
        connection_7__6__10_, connection_7__6__9_, connection_7__6__8_, 
        connection_7__6__7_, connection_7__6__6_, connection_7__6__5_, 
        connection_7__6__4_, connection_7__6__3_, connection_7__6__2_, 
        connection_7__6__1_, connection_7__6__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[57:56]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_28 second_half_stages_6__group_sec_half_0__switch_sec_half_4__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_6__12_, 
        connection_valid_6__4_}), .i_data_bus({connection_6__12__31_, 
        connection_6__12__30_, connection_6__12__29_, connection_6__12__28_, 
        connection_6__12__27_, connection_6__12__26_, connection_6__12__25_, 
        connection_6__12__24_, connection_6__12__23_, connection_6__12__22_, 
        connection_6__12__21_, connection_6__12__20_, connection_6__12__19_, 
        connection_6__12__18_, connection_6__12__17_, connection_6__12__16_, 
        connection_6__12__15_, connection_6__12__14_, connection_6__12__13_, 
        connection_6__12__12_, connection_6__12__11_, connection_6__12__10_, 
        connection_6__12__9_, connection_6__12__8_, connection_6__12__7_, 
        connection_6__12__6_, connection_6__12__5_, connection_6__12__4_, 
        connection_6__12__3_, connection_6__12__2_, connection_6__12__1_, 
        connection_6__12__0_, connection_6__4__31_, connection_6__4__30_, 
        connection_6__4__29_, connection_6__4__28_, connection_6__4__27_, 
        connection_6__4__26_, connection_6__4__25_, connection_6__4__24_, 
        connection_6__4__23_, connection_6__4__22_, connection_6__4__21_, 
        connection_6__4__20_, connection_6__4__19_, connection_6__4__18_, 
        connection_6__4__17_, connection_6__4__16_, connection_6__4__15_, 
        connection_6__4__14_, connection_6__4__13_, connection_6__4__12_, 
        connection_6__4__11_, connection_6__4__10_, connection_6__4__9_, 
        connection_6__4__8_, connection_6__4__7_, connection_6__4__6_, 
        connection_6__4__5_, connection_6__4__4_, connection_6__4__3_, 
        connection_6__4__2_, connection_6__4__1_, connection_6__4__0_}), 
        .o_valid({connection_valid_7__9_, connection_valid_7__8_}), 
        .o_data_bus({connection_7__9__31_, connection_7__9__30_, 
        connection_7__9__29_, connection_7__9__28_, connection_7__9__27_, 
        connection_7__9__26_, connection_7__9__25_, connection_7__9__24_, 
        connection_7__9__23_, connection_7__9__22_, connection_7__9__21_, 
        connection_7__9__20_, connection_7__9__19_, connection_7__9__18_, 
        connection_7__9__17_, connection_7__9__16_, connection_7__9__15_, 
        connection_7__9__14_, connection_7__9__13_, connection_7__9__12_, 
        connection_7__9__11_, connection_7__9__10_, connection_7__9__9_, 
        connection_7__9__8_, connection_7__9__7_, connection_7__9__6_, 
        connection_7__9__5_, connection_7__9__4_, connection_7__9__3_, 
        connection_7__9__2_, connection_7__9__1_, connection_7__9__0_, 
        connection_7__8__31_, connection_7__8__30_, connection_7__8__29_, 
        connection_7__8__28_, connection_7__8__27_, connection_7__8__26_, 
        connection_7__8__25_, connection_7__8__24_, connection_7__8__23_, 
        connection_7__8__22_, connection_7__8__21_, connection_7__8__20_, 
        connection_7__8__19_, connection_7__8__18_, connection_7__8__17_, 
        connection_7__8__16_, connection_7__8__15_, connection_7__8__14_, 
        connection_7__8__13_, connection_7__8__12_, connection_7__8__11_, 
        connection_7__8__10_, connection_7__8__9_, connection_7__8__8_, 
        connection_7__8__7_, connection_7__8__6_, connection_7__8__5_, 
        connection_7__8__4_, connection_7__8__3_, connection_7__8__2_, 
        connection_7__8__1_, connection_7__8__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[55:54]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_27 second_half_stages_6__group_sec_half_0__switch_sec_half_5__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_6__13_, 
        connection_valid_6__5_}), .i_data_bus({connection_6__13__31_, 
        connection_6__13__30_, connection_6__13__29_, connection_6__13__28_, 
        connection_6__13__27_, connection_6__13__26_, connection_6__13__25_, 
        connection_6__13__24_, connection_6__13__23_, connection_6__13__22_, 
        connection_6__13__21_, connection_6__13__20_, connection_6__13__19_, 
        connection_6__13__18_, connection_6__13__17_, connection_6__13__16_, 
        connection_6__13__15_, connection_6__13__14_, connection_6__13__13_, 
        connection_6__13__12_, connection_6__13__11_, connection_6__13__10_, 
        connection_6__13__9_, connection_6__13__8_, connection_6__13__7_, 
        connection_6__13__6_, connection_6__13__5_, connection_6__13__4_, 
        connection_6__13__3_, connection_6__13__2_, connection_6__13__1_, 
        connection_6__13__0_, connection_6__5__31_, connection_6__5__30_, 
        connection_6__5__29_, connection_6__5__28_, connection_6__5__27_, 
        connection_6__5__26_, connection_6__5__25_, connection_6__5__24_, 
        connection_6__5__23_, connection_6__5__22_, connection_6__5__21_, 
        connection_6__5__20_, connection_6__5__19_, connection_6__5__18_, 
        connection_6__5__17_, connection_6__5__16_, connection_6__5__15_, 
        connection_6__5__14_, connection_6__5__13_, connection_6__5__12_, 
        connection_6__5__11_, connection_6__5__10_, connection_6__5__9_, 
        connection_6__5__8_, connection_6__5__7_, connection_6__5__6_, 
        connection_6__5__5_, connection_6__5__4_, connection_6__5__3_, 
        connection_6__5__2_, connection_6__5__1_, connection_6__5__0_}), 
        .o_valid({connection_valid_7__11_, connection_valid_7__10_}), 
        .o_data_bus({connection_7__11__31_, connection_7__11__30_, 
        connection_7__11__29_, connection_7__11__28_, connection_7__11__27_, 
        connection_7__11__26_, connection_7__11__25_, connection_7__11__24_, 
        connection_7__11__23_, connection_7__11__22_, connection_7__11__21_, 
        connection_7__11__20_, connection_7__11__19_, connection_7__11__18_, 
        connection_7__11__17_, connection_7__11__16_, connection_7__11__15_, 
        connection_7__11__14_, connection_7__11__13_, connection_7__11__12_, 
        connection_7__11__11_, connection_7__11__10_, connection_7__11__9_, 
        connection_7__11__8_, connection_7__11__7_, connection_7__11__6_, 
        connection_7__11__5_, connection_7__11__4_, connection_7__11__3_, 
        connection_7__11__2_, connection_7__11__1_, connection_7__11__0_, 
        connection_7__10__31_, connection_7__10__30_, connection_7__10__29_, 
        connection_7__10__28_, connection_7__10__27_, connection_7__10__26_, 
        connection_7__10__25_, connection_7__10__24_, connection_7__10__23_, 
        connection_7__10__22_, connection_7__10__21_, connection_7__10__20_, 
        connection_7__10__19_, connection_7__10__18_, connection_7__10__17_, 
        connection_7__10__16_, connection_7__10__15_, connection_7__10__14_, 
        connection_7__10__13_, connection_7__10__12_, connection_7__10__11_, 
        connection_7__10__10_, connection_7__10__9_, connection_7__10__8_, 
        connection_7__10__7_, connection_7__10__6_, connection_7__10__5_, 
        connection_7__10__4_, connection_7__10__3_, connection_7__10__2_, 
        connection_7__10__1_, connection_7__10__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[53:52]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_26 second_half_stages_6__group_sec_half_0__switch_sec_half_6__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_6__14_, 
        connection_valid_6__6_}), .i_data_bus({connection_6__14__31_, 
        connection_6__14__30_, connection_6__14__29_, connection_6__14__28_, 
        connection_6__14__27_, connection_6__14__26_, connection_6__14__25_, 
        connection_6__14__24_, connection_6__14__23_, connection_6__14__22_, 
        connection_6__14__21_, connection_6__14__20_, connection_6__14__19_, 
        connection_6__14__18_, connection_6__14__17_, connection_6__14__16_, 
        connection_6__14__15_, connection_6__14__14_, connection_6__14__13_, 
        connection_6__14__12_, connection_6__14__11_, connection_6__14__10_, 
        connection_6__14__9_, connection_6__14__8_, connection_6__14__7_, 
        connection_6__14__6_, connection_6__14__5_, connection_6__14__4_, 
        connection_6__14__3_, connection_6__14__2_, connection_6__14__1_, 
        connection_6__14__0_, connection_6__6__31_, connection_6__6__30_, 
        connection_6__6__29_, connection_6__6__28_, connection_6__6__27_, 
        connection_6__6__26_, connection_6__6__25_, connection_6__6__24_, 
        connection_6__6__23_, connection_6__6__22_, connection_6__6__21_, 
        connection_6__6__20_, connection_6__6__19_, connection_6__6__18_, 
        connection_6__6__17_, connection_6__6__16_, connection_6__6__15_, 
        connection_6__6__14_, connection_6__6__13_, connection_6__6__12_, 
        connection_6__6__11_, connection_6__6__10_, connection_6__6__9_, 
        connection_6__6__8_, connection_6__6__7_, connection_6__6__6_, 
        connection_6__6__5_, connection_6__6__4_, connection_6__6__3_, 
        connection_6__6__2_, connection_6__6__1_, connection_6__6__0_}), 
        .o_valid({connection_valid_7__13_, connection_valid_7__12_}), 
        .o_data_bus({connection_7__13__31_, connection_7__13__30_, 
        connection_7__13__29_, connection_7__13__28_, connection_7__13__27_, 
        connection_7__13__26_, connection_7__13__25_, connection_7__13__24_, 
        connection_7__13__23_, connection_7__13__22_, connection_7__13__21_, 
        connection_7__13__20_, connection_7__13__19_, connection_7__13__18_, 
        connection_7__13__17_, connection_7__13__16_, connection_7__13__15_, 
        connection_7__13__14_, connection_7__13__13_, connection_7__13__12_, 
        connection_7__13__11_, connection_7__13__10_, connection_7__13__9_, 
        connection_7__13__8_, connection_7__13__7_, connection_7__13__6_, 
        connection_7__13__5_, connection_7__13__4_, connection_7__13__3_, 
        connection_7__13__2_, connection_7__13__1_, connection_7__13__0_, 
        connection_7__12__31_, connection_7__12__30_, connection_7__12__29_, 
        connection_7__12__28_, connection_7__12__27_, connection_7__12__26_, 
        connection_7__12__25_, connection_7__12__24_, connection_7__12__23_, 
        connection_7__12__22_, connection_7__12__21_, connection_7__12__20_, 
        connection_7__12__19_, connection_7__12__18_, connection_7__12__17_, 
        connection_7__12__16_, connection_7__12__15_, connection_7__12__14_, 
        connection_7__12__13_, connection_7__12__12_, connection_7__12__11_, 
        connection_7__12__10_, connection_7__12__9_, connection_7__12__8_, 
        connection_7__12__7_, connection_7__12__6_, connection_7__12__5_, 
        connection_7__12__4_, connection_7__12__3_, connection_7__12__2_, 
        connection_7__12__1_, connection_7__12__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[51:50]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_25 second_half_stages_6__group_sec_half_0__switch_sec_half_7__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_6__15_, 
        connection_valid_6__7_}), .i_data_bus({connection_6__15__31_, 
        connection_6__15__30_, connection_6__15__29_, connection_6__15__28_, 
        connection_6__15__27_, connection_6__15__26_, connection_6__15__25_, 
        connection_6__15__24_, connection_6__15__23_, connection_6__15__22_, 
        connection_6__15__21_, connection_6__15__20_, connection_6__15__19_, 
        connection_6__15__18_, connection_6__15__17_, connection_6__15__16_, 
        connection_6__15__15_, connection_6__15__14_, connection_6__15__13_, 
        connection_6__15__12_, connection_6__15__11_, connection_6__15__10_, 
        connection_6__15__9_, connection_6__15__8_, connection_6__15__7_, 
        connection_6__15__6_, connection_6__15__5_, connection_6__15__4_, 
        connection_6__15__3_, connection_6__15__2_, connection_6__15__1_, 
        connection_6__15__0_, connection_6__7__31_, connection_6__7__30_, 
        connection_6__7__29_, connection_6__7__28_, connection_6__7__27_, 
        connection_6__7__26_, connection_6__7__25_, connection_6__7__24_, 
        connection_6__7__23_, connection_6__7__22_, connection_6__7__21_, 
        connection_6__7__20_, connection_6__7__19_, connection_6__7__18_, 
        connection_6__7__17_, connection_6__7__16_, connection_6__7__15_, 
        connection_6__7__14_, connection_6__7__13_, connection_6__7__12_, 
        connection_6__7__11_, connection_6__7__10_, connection_6__7__9_, 
        connection_6__7__8_, connection_6__7__7_, connection_6__7__6_, 
        connection_6__7__5_, connection_6__7__4_, connection_6__7__3_, 
        connection_6__7__2_, connection_6__7__1_, connection_6__7__0_}), 
        .o_valid({connection_valid_7__15_, connection_valid_7__14_}), 
        .o_data_bus({connection_7__15__31_, connection_7__15__30_, 
        connection_7__15__29_, connection_7__15__28_, connection_7__15__27_, 
        connection_7__15__26_, connection_7__15__25_, connection_7__15__24_, 
        connection_7__15__23_, connection_7__15__22_, connection_7__15__21_, 
        connection_7__15__20_, connection_7__15__19_, connection_7__15__18_, 
        connection_7__15__17_, connection_7__15__16_, connection_7__15__15_, 
        connection_7__15__14_, connection_7__15__13_, connection_7__15__12_, 
        connection_7__15__11_, connection_7__15__10_, connection_7__15__9_, 
        connection_7__15__8_, connection_7__15__7_, connection_7__15__6_, 
        connection_7__15__5_, connection_7__15__4_, connection_7__15__3_, 
        connection_7__15__2_, connection_7__15__1_, connection_7__15__0_, 
        connection_7__14__31_, connection_7__14__30_, connection_7__14__29_, 
        connection_7__14__28_, connection_7__14__27_, connection_7__14__26_, 
        connection_7__14__25_, connection_7__14__24_, connection_7__14__23_, 
        connection_7__14__22_, connection_7__14__21_, connection_7__14__20_, 
        connection_7__14__19_, connection_7__14__18_, connection_7__14__17_, 
        connection_7__14__16_, connection_7__14__15_, connection_7__14__14_, 
        connection_7__14__13_, connection_7__14__12_, connection_7__14__11_, 
        connection_7__14__10_, connection_7__14__9_, connection_7__14__8_, 
        connection_7__14__7_, connection_7__14__6_, connection_7__14__5_, 
        connection_7__14__4_, connection_7__14__3_, connection_7__14__2_, 
        connection_7__14__1_, connection_7__14__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[49:48]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_24 second_half_stages_6__group_sec_half_1__switch_sec_half_0__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_6__24_, 
        connection_valid_6__16_}), .i_data_bus({connection_6__24__31_, 
        connection_6__24__30_, connection_6__24__29_, connection_6__24__28_, 
        connection_6__24__27_, connection_6__24__26_, connection_6__24__25_, 
        connection_6__24__24_, connection_6__24__23_, connection_6__24__22_, 
        connection_6__24__21_, connection_6__24__20_, connection_6__24__19_, 
        connection_6__24__18_, connection_6__24__17_, connection_6__24__16_, 
        connection_6__24__15_, connection_6__24__14_, connection_6__24__13_, 
        connection_6__24__12_, connection_6__24__11_, connection_6__24__10_, 
        connection_6__24__9_, connection_6__24__8_, connection_6__24__7_, 
        connection_6__24__6_, connection_6__24__5_, connection_6__24__4_, 
        connection_6__24__3_, connection_6__24__2_, connection_6__24__1_, 
        connection_6__24__0_, connection_6__16__31_, connection_6__16__30_, 
        connection_6__16__29_, connection_6__16__28_, connection_6__16__27_, 
        connection_6__16__26_, connection_6__16__25_, connection_6__16__24_, 
        connection_6__16__23_, connection_6__16__22_, connection_6__16__21_, 
        connection_6__16__20_, connection_6__16__19_, connection_6__16__18_, 
        connection_6__16__17_, connection_6__16__16_, connection_6__16__15_, 
        connection_6__16__14_, connection_6__16__13_, connection_6__16__12_, 
        connection_6__16__11_, connection_6__16__10_, connection_6__16__9_, 
        connection_6__16__8_, connection_6__16__7_, connection_6__16__6_, 
        connection_6__16__5_, connection_6__16__4_, connection_6__16__3_, 
        connection_6__16__2_, connection_6__16__1_, connection_6__16__0_}), 
        .o_valid({connection_valid_7__17_, connection_valid_7__16_}), 
        .o_data_bus({connection_7__17__31_, connection_7__17__30_, 
        connection_7__17__29_, connection_7__17__28_, connection_7__17__27_, 
        connection_7__17__26_, connection_7__17__25_, connection_7__17__24_, 
        connection_7__17__23_, connection_7__17__22_, connection_7__17__21_, 
        connection_7__17__20_, connection_7__17__19_, connection_7__17__18_, 
        connection_7__17__17_, connection_7__17__16_, connection_7__17__15_, 
        connection_7__17__14_, connection_7__17__13_, connection_7__17__12_, 
        connection_7__17__11_, connection_7__17__10_, connection_7__17__9_, 
        connection_7__17__8_, connection_7__17__7_, connection_7__17__6_, 
        connection_7__17__5_, connection_7__17__4_, connection_7__17__3_, 
        connection_7__17__2_, connection_7__17__1_, connection_7__17__0_, 
        connection_7__16__31_, connection_7__16__30_, connection_7__16__29_, 
        connection_7__16__28_, connection_7__16__27_, connection_7__16__26_, 
        connection_7__16__25_, connection_7__16__24_, connection_7__16__23_, 
        connection_7__16__22_, connection_7__16__21_, connection_7__16__20_, 
        connection_7__16__19_, connection_7__16__18_, connection_7__16__17_, 
        connection_7__16__16_, connection_7__16__15_, connection_7__16__14_, 
        connection_7__16__13_, connection_7__16__12_, connection_7__16__11_, 
        connection_7__16__10_, connection_7__16__9_, connection_7__16__8_, 
        connection_7__16__7_, connection_7__16__6_, connection_7__16__5_, 
        connection_7__16__4_, connection_7__16__3_, connection_7__16__2_, 
        connection_7__16__1_, connection_7__16__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[47:46]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_23 second_half_stages_6__group_sec_half_1__switch_sec_half_1__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_6__25_, 
        connection_valid_6__17_}), .i_data_bus({connection_6__25__31_, 
        connection_6__25__30_, connection_6__25__29_, connection_6__25__28_, 
        connection_6__25__27_, connection_6__25__26_, connection_6__25__25_, 
        connection_6__25__24_, connection_6__25__23_, connection_6__25__22_, 
        connection_6__25__21_, connection_6__25__20_, connection_6__25__19_, 
        connection_6__25__18_, connection_6__25__17_, connection_6__25__16_, 
        connection_6__25__15_, connection_6__25__14_, connection_6__25__13_, 
        connection_6__25__12_, connection_6__25__11_, connection_6__25__10_, 
        connection_6__25__9_, connection_6__25__8_, connection_6__25__7_, 
        connection_6__25__6_, connection_6__25__5_, connection_6__25__4_, 
        connection_6__25__3_, connection_6__25__2_, connection_6__25__1_, 
        connection_6__25__0_, connection_6__17__31_, connection_6__17__30_, 
        connection_6__17__29_, connection_6__17__28_, connection_6__17__27_, 
        connection_6__17__26_, connection_6__17__25_, connection_6__17__24_, 
        connection_6__17__23_, connection_6__17__22_, connection_6__17__21_, 
        connection_6__17__20_, connection_6__17__19_, connection_6__17__18_, 
        connection_6__17__17_, connection_6__17__16_, connection_6__17__15_, 
        connection_6__17__14_, connection_6__17__13_, connection_6__17__12_, 
        connection_6__17__11_, connection_6__17__10_, connection_6__17__9_, 
        connection_6__17__8_, connection_6__17__7_, connection_6__17__6_, 
        connection_6__17__5_, connection_6__17__4_, connection_6__17__3_, 
        connection_6__17__2_, connection_6__17__1_, connection_6__17__0_}), 
        .o_valid({connection_valid_7__19_, connection_valid_7__18_}), 
        .o_data_bus({connection_7__19__31_, connection_7__19__30_, 
        connection_7__19__29_, connection_7__19__28_, connection_7__19__27_, 
        connection_7__19__26_, connection_7__19__25_, connection_7__19__24_, 
        connection_7__19__23_, connection_7__19__22_, connection_7__19__21_, 
        connection_7__19__20_, connection_7__19__19_, connection_7__19__18_, 
        connection_7__19__17_, connection_7__19__16_, connection_7__19__15_, 
        connection_7__19__14_, connection_7__19__13_, connection_7__19__12_, 
        connection_7__19__11_, connection_7__19__10_, connection_7__19__9_, 
        connection_7__19__8_, connection_7__19__7_, connection_7__19__6_, 
        connection_7__19__5_, connection_7__19__4_, connection_7__19__3_, 
        connection_7__19__2_, connection_7__19__1_, connection_7__19__0_, 
        connection_7__18__31_, connection_7__18__30_, connection_7__18__29_, 
        connection_7__18__28_, connection_7__18__27_, connection_7__18__26_, 
        connection_7__18__25_, connection_7__18__24_, connection_7__18__23_, 
        connection_7__18__22_, connection_7__18__21_, connection_7__18__20_, 
        connection_7__18__19_, connection_7__18__18_, connection_7__18__17_, 
        connection_7__18__16_, connection_7__18__15_, connection_7__18__14_, 
        connection_7__18__13_, connection_7__18__12_, connection_7__18__11_, 
        connection_7__18__10_, connection_7__18__9_, connection_7__18__8_, 
        connection_7__18__7_, connection_7__18__6_, connection_7__18__5_, 
        connection_7__18__4_, connection_7__18__3_, connection_7__18__2_, 
        connection_7__18__1_, connection_7__18__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[45:44]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_22 second_half_stages_6__group_sec_half_1__switch_sec_half_2__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_6__26_, 
        connection_valid_6__18_}), .i_data_bus({connection_6__26__31_, 
        connection_6__26__30_, connection_6__26__29_, connection_6__26__28_, 
        connection_6__26__27_, connection_6__26__26_, connection_6__26__25_, 
        connection_6__26__24_, connection_6__26__23_, connection_6__26__22_, 
        connection_6__26__21_, connection_6__26__20_, connection_6__26__19_, 
        connection_6__26__18_, connection_6__26__17_, connection_6__26__16_, 
        connection_6__26__15_, connection_6__26__14_, connection_6__26__13_, 
        connection_6__26__12_, connection_6__26__11_, connection_6__26__10_, 
        connection_6__26__9_, connection_6__26__8_, connection_6__26__7_, 
        connection_6__26__6_, connection_6__26__5_, connection_6__26__4_, 
        connection_6__26__3_, connection_6__26__2_, connection_6__26__1_, 
        connection_6__26__0_, connection_6__18__31_, connection_6__18__30_, 
        connection_6__18__29_, connection_6__18__28_, connection_6__18__27_, 
        connection_6__18__26_, connection_6__18__25_, connection_6__18__24_, 
        connection_6__18__23_, connection_6__18__22_, connection_6__18__21_, 
        connection_6__18__20_, connection_6__18__19_, connection_6__18__18_, 
        connection_6__18__17_, connection_6__18__16_, connection_6__18__15_, 
        connection_6__18__14_, connection_6__18__13_, connection_6__18__12_, 
        connection_6__18__11_, connection_6__18__10_, connection_6__18__9_, 
        connection_6__18__8_, connection_6__18__7_, connection_6__18__6_, 
        connection_6__18__5_, connection_6__18__4_, connection_6__18__3_, 
        connection_6__18__2_, connection_6__18__1_, connection_6__18__0_}), 
        .o_valid({connection_valid_7__21_, connection_valid_7__20_}), 
        .o_data_bus({connection_7__21__31_, connection_7__21__30_, 
        connection_7__21__29_, connection_7__21__28_, connection_7__21__27_, 
        connection_7__21__26_, connection_7__21__25_, connection_7__21__24_, 
        connection_7__21__23_, connection_7__21__22_, connection_7__21__21_, 
        connection_7__21__20_, connection_7__21__19_, connection_7__21__18_, 
        connection_7__21__17_, connection_7__21__16_, connection_7__21__15_, 
        connection_7__21__14_, connection_7__21__13_, connection_7__21__12_, 
        connection_7__21__11_, connection_7__21__10_, connection_7__21__9_, 
        connection_7__21__8_, connection_7__21__7_, connection_7__21__6_, 
        connection_7__21__5_, connection_7__21__4_, connection_7__21__3_, 
        connection_7__21__2_, connection_7__21__1_, connection_7__21__0_, 
        connection_7__20__31_, connection_7__20__30_, connection_7__20__29_, 
        connection_7__20__28_, connection_7__20__27_, connection_7__20__26_, 
        connection_7__20__25_, connection_7__20__24_, connection_7__20__23_, 
        connection_7__20__22_, connection_7__20__21_, connection_7__20__20_, 
        connection_7__20__19_, connection_7__20__18_, connection_7__20__17_, 
        connection_7__20__16_, connection_7__20__15_, connection_7__20__14_, 
        connection_7__20__13_, connection_7__20__12_, connection_7__20__11_, 
        connection_7__20__10_, connection_7__20__9_, connection_7__20__8_, 
        connection_7__20__7_, connection_7__20__6_, connection_7__20__5_, 
        connection_7__20__4_, connection_7__20__3_, connection_7__20__2_, 
        connection_7__20__1_, connection_7__20__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[43:42]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_21 second_half_stages_6__group_sec_half_1__switch_sec_half_3__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_6__27_, 
        connection_valid_6__19_}), .i_data_bus({connection_6__27__31_, 
        connection_6__27__30_, connection_6__27__29_, connection_6__27__28_, 
        connection_6__27__27_, connection_6__27__26_, connection_6__27__25_, 
        connection_6__27__24_, connection_6__27__23_, connection_6__27__22_, 
        connection_6__27__21_, connection_6__27__20_, connection_6__27__19_, 
        connection_6__27__18_, connection_6__27__17_, connection_6__27__16_, 
        connection_6__27__15_, connection_6__27__14_, connection_6__27__13_, 
        connection_6__27__12_, connection_6__27__11_, connection_6__27__10_, 
        connection_6__27__9_, connection_6__27__8_, connection_6__27__7_, 
        connection_6__27__6_, connection_6__27__5_, connection_6__27__4_, 
        connection_6__27__3_, connection_6__27__2_, connection_6__27__1_, 
        connection_6__27__0_, connection_6__19__31_, connection_6__19__30_, 
        connection_6__19__29_, connection_6__19__28_, connection_6__19__27_, 
        connection_6__19__26_, connection_6__19__25_, connection_6__19__24_, 
        connection_6__19__23_, connection_6__19__22_, connection_6__19__21_, 
        connection_6__19__20_, connection_6__19__19_, connection_6__19__18_, 
        connection_6__19__17_, connection_6__19__16_, connection_6__19__15_, 
        connection_6__19__14_, connection_6__19__13_, connection_6__19__12_, 
        connection_6__19__11_, connection_6__19__10_, connection_6__19__9_, 
        connection_6__19__8_, connection_6__19__7_, connection_6__19__6_, 
        connection_6__19__5_, connection_6__19__4_, connection_6__19__3_, 
        connection_6__19__2_, connection_6__19__1_, connection_6__19__0_}), 
        .o_valid({connection_valid_7__23_, connection_valid_7__22_}), 
        .o_data_bus({connection_7__23__31_, connection_7__23__30_, 
        connection_7__23__29_, connection_7__23__28_, connection_7__23__27_, 
        connection_7__23__26_, connection_7__23__25_, connection_7__23__24_, 
        connection_7__23__23_, connection_7__23__22_, connection_7__23__21_, 
        connection_7__23__20_, connection_7__23__19_, connection_7__23__18_, 
        connection_7__23__17_, connection_7__23__16_, connection_7__23__15_, 
        connection_7__23__14_, connection_7__23__13_, connection_7__23__12_, 
        connection_7__23__11_, connection_7__23__10_, connection_7__23__9_, 
        connection_7__23__8_, connection_7__23__7_, connection_7__23__6_, 
        connection_7__23__5_, connection_7__23__4_, connection_7__23__3_, 
        connection_7__23__2_, connection_7__23__1_, connection_7__23__0_, 
        connection_7__22__31_, connection_7__22__30_, connection_7__22__29_, 
        connection_7__22__28_, connection_7__22__27_, connection_7__22__26_, 
        connection_7__22__25_, connection_7__22__24_, connection_7__22__23_, 
        connection_7__22__22_, connection_7__22__21_, connection_7__22__20_, 
        connection_7__22__19_, connection_7__22__18_, connection_7__22__17_, 
        connection_7__22__16_, connection_7__22__15_, connection_7__22__14_, 
        connection_7__22__13_, connection_7__22__12_, connection_7__22__11_, 
        connection_7__22__10_, connection_7__22__9_, connection_7__22__8_, 
        connection_7__22__7_, connection_7__22__6_, connection_7__22__5_, 
        connection_7__22__4_, connection_7__22__3_, connection_7__22__2_, 
        connection_7__22__1_, connection_7__22__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[41:40]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_20 second_half_stages_6__group_sec_half_1__switch_sec_half_4__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_6__28_, 
        connection_valid_6__20_}), .i_data_bus({connection_6__28__31_, 
        connection_6__28__30_, connection_6__28__29_, connection_6__28__28_, 
        connection_6__28__27_, connection_6__28__26_, connection_6__28__25_, 
        connection_6__28__24_, connection_6__28__23_, connection_6__28__22_, 
        connection_6__28__21_, connection_6__28__20_, connection_6__28__19_, 
        connection_6__28__18_, connection_6__28__17_, connection_6__28__16_, 
        connection_6__28__15_, connection_6__28__14_, connection_6__28__13_, 
        connection_6__28__12_, connection_6__28__11_, connection_6__28__10_, 
        connection_6__28__9_, connection_6__28__8_, connection_6__28__7_, 
        connection_6__28__6_, connection_6__28__5_, connection_6__28__4_, 
        connection_6__28__3_, connection_6__28__2_, connection_6__28__1_, 
        connection_6__28__0_, connection_6__20__31_, connection_6__20__30_, 
        connection_6__20__29_, connection_6__20__28_, connection_6__20__27_, 
        connection_6__20__26_, connection_6__20__25_, connection_6__20__24_, 
        connection_6__20__23_, connection_6__20__22_, connection_6__20__21_, 
        connection_6__20__20_, connection_6__20__19_, connection_6__20__18_, 
        connection_6__20__17_, connection_6__20__16_, connection_6__20__15_, 
        connection_6__20__14_, connection_6__20__13_, connection_6__20__12_, 
        connection_6__20__11_, connection_6__20__10_, connection_6__20__9_, 
        connection_6__20__8_, connection_6__20__7_, connection_6__20__6_, 
        connection_6__20__5_, connection_6__20__4_, connection_6__20__3_, 
        connection_6__20__2_, connection_6__20__1_, connection_6__20__0_}), 
        .o_valid({connection_valid_7__25_, connection_valid_7__24_}), 
        .o_data_bus({connection_7__25__31_, connection_7__25__30_, 
        connection_7__25__29_, connection_7__25__28_, connection_7__25__27_, 
        connection_7__25__26_, connection_7__25__25_, connection_7__25__24_, 
        connection_7__25__23_, connection_7__25__22_, connection_7__25__21_, 
        connection_7__25__20_, connection_7__25__19_, connection_7__25__18_, 
        connection_7__25__17_, connection_7__25__16_, connection_7__25__15_, 
        connection_7__25__14_, connection_7__25__13_, connection_7__25__12_, 
        connection_7__25__11_, connection_7__25__10_, connection_7__25__9_, 
        connection_7__25__8_, connection_7__25__7_, connection_7__25__6_, 
        connection_7__25__5_, connection_7__25__4_, connection_7__25__3_, 
        connection_7__25__2_, connection_7__25__1_, connection_7__25__0_, 
        connection_7__24__31_, connection_7__24__30_, connection_7__24__29_, 
        connection_7__24__28_, connection_7__24__27_, connection_7__24__26_, 
        connection_7__24__25_, connection_7__24__24_, connection_7__24__23_, 
        connection_7__24__22_, connection_7__24__21_, connection_7__24__20_, 
        connection_7__24__19_, connection_7__24__18_, connection_7__24__17_, 
        connection_7__24__16_, connection_7__24__15_, connection_7__24__14_, 
        connection_7__24__13_, connection_7__24__12_, connection_7__24__11_, 
        connection_7__24__10_, connection_7__24__9_, connection_7__24__8_, 
        connection_7__24__7_, connection_7__24__6_, connection_7__24__5_, 
        connection_7__24__4_, connection_7__24__3_, connection_7__24__2_, 
        connection_7__24__1_, connection_7__24__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[39:38]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_19 second_half_stages_6__group_sec_half_1__switch_sec_half_5__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_6__29_, 
        connection_valid_6__21_}), .i_data_bus({connection_6__29__31_, 
        connection_6__29__30_, connection_6__29__29_, connection_6__29__28_, 
        connection_6__29__27_, connection_6__29__26_, connection_6__29__25_, 
        connection_6__29__24_, connection_6__29__23_, connection_6__29__22_, 
        connection_6__29__21_, connection_6__29__20_, connection_6__29__19_, 
        connection_6__29__18_, connection_6__29__17_, connection_6__29__16_, 
        connection_6__29__15_, connection_6__29__14_, connection_6__29__13_, 
        connection_6__29__12_, connection_6__29__11_, connection_6__29__10_, 
        connection_6__29__9_, connection_6__29__8_, connection_6__29__7_, 
        connection_6__29__6_, connection_6__29__5_, connection_6__29__4_, 
        connection_6__29__3_, connection_6__29__2_, connection_6__29__1_, 
        connection_6__29__0_, connection_6__21__31_, connection_6__21__30_, 
        connection_6__21__29_, connection_6__21__28_, connection_6__21__27_, 
        connection_6__21__26_, connection_6__21__25_, connection_6__21__24_, 
        connection_6__21__23_, connection_6__21__22_, connection_6__21__21_, 
        connection_6__21__20_, connection_6__21__19_, connection_6__21__18_, 
        connection_6__21__17_, connection_6__21__16_, connection_6__21__15_, 
        connection_6__21__14_, connection_6__21__13_, connection_6__21__12_, 
        connection_6__21__11_, connection_6__21__10_, connection_6__21__9_, 
        connection_6__21__8_, connection_6__21__7_, connection_6__21__6_, 
        connection_6__21__5_, connection_6__21__4_, connection_6__21__3_, 
        connection_6__21__2_, connection_6__21__1_, connection_6__21__0_}), 
        .o_valid({connection_valid_7__27_, connection_valid_7__26_}), 
        .o_data_bus({connection_7__27__31_, connection_7__27__30_, 
        connection_7__27__29_, connection_7__27__28_, connection_7__27__27_, 
        connection_7__27__26_, connection_7__27__25_, connection_7__27__24_, 
        connection_7__27__23_, connection_7__27__22_, connection_7__27__21_, 
        connection_7__27__20_, connection_7__27__19_, connection_7__27__18_, 
        connection_7__27__17_, connection_7__27__16_, connection_7__27__15_, 
        connection_7__27__14_, connection_7__27__13_, connection_7__27__12_, 
        connection_7__27__11_, connection_7__27__10_, connection_7__27__9_, 
        connection_7__27__8_, connection_7__27__7_, connection_7__27__6_, 
        connection_7__27__5_, connection_7__27__4_, connection_7__27__3_, 
        connection_7__27__2_, connection_7__27__1_, connection_7__27__0_, 
        connection_7__26__31_, connection_7__26__30_, connection_7__26__29_, 
        connection_7__26__28_, connection_7__26__27_, connection_7__26__26_, 
        connection_7__26__25_, connection_7__26__24_, connection_7__26__23_, 
        connection_7__26__22_, connection_7__26__21_, connection_7__26__20_, 
        connection_7__26__19_, connection_7__26__18_, connection_7__26__17_, 
        connection_7__26__16_, connection_7__26__15_, connection_7__26__14_, 
        connection_7__26__13_, connection_7__26__12_, connection_7__26__11_, 
        connection_7__26__10_, connection_7__26__9_, connection_7__26__8_, 
        connection_7__26__7_, connection_7__26__6_, connection_7__26__5_, 
        connection_7__26__4_, connection_7__26__3_, connection_7__26__2_, 
        connection_7__26__1_, connection_7__26__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[37:36]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_18 second_half_stages_6__group_sec_half_1__switch_sec_half_6__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_6__30_, 
        connection_valid_6__22_}), .i_data_bus({connection_6__30__31_, 
        connection_6__30__30_, connection_6__30__29_, connection_6__30__28_, 
        connection_6__30__27_, connection_6__30__26_, connection_6__30__25_, 
        connection_6__30__24_, connection_6__30__23_, connection_6__30__22_, 
        connection_6__30__21_, connection_6__30__20_, connection_6__30__19_, 
        connection_6__30__18_, connection_6__30__17_, connection_6__30__16_, 
        connection_6__30__15_, connection_6__30__14_, connection_6__30__13_, 
        connection_6__30__12_, connection_6__30__11_, connection_6__30__10_, 
        connection_6__30__9_, connection_6__30__8_, connection_6__30__7_, 
        connection_6__30__6_, connection_6__30__5_, connection_6__30__4_, 
        connection_6__30__3_, connection_6__30__2_, connection_6__30__1_, 
        connection_6__30__0_, connection_6__22__31_, connection_6__22__30_, 
        connection_6__22__29_, connection_6__22__28_, connection_6__22__27_, 
        connection_6__22__26_, connection_6__22__25_, connection_6__22__24_, 
        connection_6__22__23_, connection_6__22__22_, connection_6__22__21_, 
        connection_6__22__20_, connection_6__22__19_, connection_6__22__18_, 
        connection_6__22__17_, connection_6__22__16_, connection_6__22__15_, 
        connection_6__22__14_, connection_6__22__13_, connection_6__22__12_, 
        connection_6__22__11_, connection_6__22__10_, connection_6__22__9_, 
        connection_6__22__8_, connection_6__22__7_, connection_6__22__6_, 
        connection_6__22__5_, connection_6__22__4_, connection_6__22__3_, 
        connection_6__22__2_, connection_6__22__1_, connection_6__22__0_}), 
        .o_valid({connection_valid_7__29_, connection_valid_7__28_}), 
        .o_data_bus({connection_7__29__31_, connection_7__29__30_, 
        connection_7__29__29_, connection_7__29__28_, connection_7__29__27_, 
        connection_7__29__26_, connection_7__29__25_, connection_7__29__24_, 
        connection_7__29__23_, connection_7__29__22_, connection_7__29__21_, 
        connection_7__29__20_, connection_7__29__19_, connection_7__29__18_, 
        connection_7__29__17_, connection_7__29__16_, connection_7__29__15_, 
        connection_7__29__14_, connection_7__29__13_, connection_7__29__12_, 
        connection_7__29__11_, connection_7__29__10_, connection_7__29__9_, 
        connection_7__29__8_, connection_7__29__7_, connection_7__29__6_, 
        connection_7__29__5_, connection_7__29__4_, connection_7__29__3_, 
        connection_7__29__2_, connection_7__29__1_, connection_7__29__0_, 
        connection_7__28__31_, connection_7__28__30_, connection_7__28__29_, 
        connection_7__28__28_, connection_7__28__27_, connection_7__28__26_, 
        connection_7__28__25_, connection_7__28__24_, connection_7__28__23_, 
        connection_7__28__22_, connection_7__28__21_, connection_7__28__20_, 
        connection_7__28__19_, connection_7__28__18_, connection_7__28__17_, 
        connection_7__28__16_, connection_7__28__15_, connection_7__28__14_, 
        connection_7__28__13_, connection_7__28__12_, connection_7__28__11_, 
        connection_7__28__10_, connection_7__28__9_, connection_7__28__8_, 
        connection_7__28__7_, connection_7__28__6_, connection_7__28__5_, 
        connection_7__28__4_, connection_7__28__3_, connection_7__28__2_, 
        connection_7__28__1_, connection_7__28__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[35:34]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_17 second_half_stages_6__group_sec_half_1__switch_sec_half_7__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_6__31_, 
        connection_valid_6__23_}), .i_data_bus({connection_6__31__31_, 
        connection_6__31__30_, connection_6__31__29_, connection_6__31__28_, 
        connection_6__31__27_, connection_6__31__26_, connection_6__31__25_, 
        connection_6__31__24_, connection_6__31__23_, connection_6__31__22_, 
        connection_6__31__21_, connection_6__31__20_, connection_6__31__19_, 
        connection_6__31__18_, connection_6__31__17_, connection_6__31__16_, 
        connection_6__31__15_, connection_6__31__14_, connection_6__31__13_, 
        connection_6__31__12_, connection_6__31__11_, connection_6__31__10_, 
        connection_6__31__9_, connection_6__31__8_, connection_6__31__7_, 
        connection_6__31__6_, connection_6__31__5_, connection_6__31__4_, 
        connection_6__31__3_, connection_6__31__2_, connection_6__31__1_, 
        connection_6__31__0_, connection_6__23__31_, connection_6__23__30_, 
        connection_6__23__29_, connection_6__23__28_, connection_6__23__27_, 
        connection_6__23__26_, connection_6__23__25_, connection_6__23__24_, 
        connection_6__23__23_, connection_6__23__22_, connection_6__23__21_, 
        connection_6__23__20_, connection_6__23__19_, connection_6__23__18_, 
        connection_6__23__17_, connection_6__23__16_, connection_6__23__15_, 
        connection_6__23__14_, connection_6__23__13_, connection_6__23__12_, 
        connection_6__23__11_, connection_6__23__10_, connection_6__23__9_, 
        connection_6__23__8_, connection_6__23__7_, connection_6__23__6_, 
        connection_6__23__5_, connection_6__23__4_, connection_6__23__3_, 
        connection_6__23__2_, connection_6__23__1_, connection_6__23__0_}), 
        .o_valid({connection_valid_7__31_, connection_valid_7__30_}), 
        .o_data_bus({connection_7__31__31_, connection_7__31__30_, 
        connection_7__31__29_, connection_7__31__28_, connection_7__31__27_, 
        connection_7__31__26_, connection_7__31__25_, connection_7__31__24_, 
        connection_7__31__23_, connection_7__31__22_, connection_7__31__21_, 
        connection_7__31__20_, connection_7__31__19_, connection_7__31__18_, 
        connection_7__31__17_, connection_7__31__16_, connection_7__31__15_, 
        connection_7__31__14_, connection_7__31__13_, connection_7__31__12_, 
        connection_7__31__11_, connection_7__31__10_, connection_7__31__9_, 
        connection_7__31__8_, connection_7__31__7_, connection_7__31__6_, 
        connection_7__31__5_, connection_7__31__4_, connection_7__31__3_, 
        connection_7__31__2_, connection_7__31__1_, connection_7__31__0_, 
        connection_7__30__31_, connection_7__30__30_, connection_7__30__29_, 
        connection_7__30__28_, connection_7__30__27_, connection_7__30__26_, 
        connection_7__30__25_, connection_7__30__24_, connection_7__30__23_, 
        connection_7__30__22_, connection_7__30__21_, connection_7__30__20_, 
        connection_7__30__19_, connection_7__30__18_, connection_7__30__17_, 
        connection_7__30__16_, connection_7__30__15_, connection_7__30__14_, 
        connection_7__30__13_, connection_7__30__12_, connection_7__30__11_, 
        connection_7__30__10_, connection_7__30__9_, connection_7__30__8_, 
        connection_7__30__7_, connection_7__30__6_, connection_7__30__5_, 
        connection_7__30__4_, connection_7__30__3_, connection_7__30__2_, 
        connection_7__30__1_, connection_7__30__0_}), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[33:32]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_16 second_half_stages_7__group_sec_half_0__switch_sec_half_0__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_7__16_, 
        connection_valid_7__0_}), .i_data_bus({connection_7__16__31_, 
        connection_7__16__30_, connection_7__16__29_, connection_7__16__28_, 
        connection_7__16__27_, connection_7__16__26_, connection_7__16__25_, 
        connection_7__16__24_, connection_7__16__23_, connection_7__16__22_, 
        connection_7__16__21_, connection_7__16__20_, connection_7__16__19_, 
        connection_7__16__18_, connection_7__16__17_, connection_7__16__16_, 
        connection_7__16__15_, connection_7__16__14_, connection_7__16__13_, 
        connection_7__16__12_, connection_7__16__11_, connection_7__16__10_, 
        connection_7__16__9_, connection_7__16__8_, connection_7__16__7_, 
        connection_7__16__6_, connection_7__16__5_, connection_7__16__4_, 
        connection_7__16__3_, connection_7__16__2_, connection_7__16__1_, 
        connection_7__16__0_, connection_7__0__31_, connection_7__0__30_, 
        connection_7__0__29_, connection_7__0__28_, connection_7__0__27_, 
        connection_7__0__26_, connection_7__0__25_, connection_7__0__24_, 
        connection_7__0__23_, connection_7__0__22_, connection_7__0__21_, 
        connection_7__0__20_, connection_7__0__19_, connection_7__0__18_, 
        connection_7__0__17_, connection_7__0__16_, connection_7__0__15_, 
        connection_7__0__14_, connection_7__0__13_, connection_7__0__12_, 
        connection_7__0__11_, connection_7__0__10_, connection_7__0__9_, 
        connection_7__0__8_, connection_7__0__7_, connection_7__0__6_, 
        connection_7__0__5_, connection_7__0__4_, connection_7__0__3_, 
        connection_7__0__2_, connection_7__0__1_, connection_7__0__0_}), 
        .o_valid({n1615, n1616}), .o_data_bus({n2577, n2578, n2579, n2580, 
        n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, 
        n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, 
        n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, 
        n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, 
        n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, 
        n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640}), 
        .i_en(i_en), .i_cmd(cmd_pipeline_stage_7__pipeline_i_cmd_reg[31:30])
         );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_15 second_half_stages_7__group_sec_half_0__switch_sec_half_1__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_7__17_, 
        connection_valid_7__1_}), .i_data_bus({connection_7__17__31_, 
        connection_7__17__30_, connection_7__17__29_, connection_7__17__28_, 
        connection_7__17__27_, connection_7__17__26_, connection_7__17__25_, 
        connection_7__17__24_, connection_7__17__23_, connection_7__17__22_, 
        connection_7__17__21_, connection_7__17__20_, connection_7__17__19_, 
        connection_7__17__18_, connection_7__17__17_, connection_7__17__16_, 
        connection_7__17__15_, connection_7__17__14_, connection_7__17__13_, 
        connection_7__17__12_, connection_7__17__11_, connection_7__17__10_, 
        connection_7__17__9_, connection_7__17__8_, connection_7__17__7_, 
        connection_7__17__6_, connection_7__17__5_, connection_7__17__4_, 
        connection_7__17__3_, connection_7__17__2_, connection_7__17__1_, 
        connection_7__17__0_, connection_7__1__31_, connection_7__1__30_, 
        connection_7__1__29_, connection_7__1__28_, connection_7__1__27_, 
        connection_7__1__26_, connection_7__1__25_, connection_7__1__24_, 
        connection_7__1__23_, connection_7__1__22_, connection_7__1__21_, 
        connection_7__1__20_, connection_7__1__19_, connection_7__1__18_, 
        connection_7__1__17_, connection_7__1__16_, connection_7__1__15_, 
        connection_7__1__14_, connection_7__1__13_, connection_7__1__12_, 
        connection_7__1__11_, connection_7__1__10_, connection_7__1__9_, 
        connection_7__1__8_, connection_7__1__7_, connection_7__1__6_, 
        connection_7__1__5_, connection_7__1__4_, connection_7__1__3_, 
        connection_7__1__2_, connection_7__1__1_, connection_7__1__0_}), 
        .o_valid({n1613, n1614}), .o_data_bus({n2513, n2514, n2515, n2516, 
        n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, 
        n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, 
        n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, 
        n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, 
        n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, 
        n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576}), 
        .i_en(i_en), .i_cmd(cmd_pipeline_stage_7__pipeline_i_cmd_reg[29:28])
         );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_14 second_half_stages_7__group_sec_half_0__switch_sec_half_2__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_7__18_, 
        connection_valid_7__2_}), .i_data_bus({connection_7__18__31_, 
        connection_7__18__30_, connection_7__18__29_, connection_7__18__28_, 
        connection_7__18__27_, connection_7__18__26_, connection_7__18__25_, 
        connection_7__18__24_, connection_7__18__23_, connection_7__18__22_, 
        connection_7__18__21_, connection_7__18__20_, connection_7__18__19_, 
        connection_7__18__18_, connection_7__18__17_, connection_7__18__16_, 
        connection_7__18__15_, connection_7__18__14_, connection_7__18__13_, 
        connection_7__18__12_, connection_7__18__11_, connection_7__18__10_, 
        connection_7__18__9_, connection_7__18__8_, connection_7__18__7_, 
        connection_7__18__6_, connection_7__18__5_, connection_7__18__4_, 
        connection_7__18__3_, connection_7__18__2_, connection_7__18__1_, 
        connection_7__18__0_, connection_7__2__31_, connection_7__2__30_, 
        connection_7__2__29_, connection_7__2__28_, connection_7__2__27_, 
        connection_7__2__26_, connection_7__2__25_, connection_7__2__24_, 
        connection_7__2__23_, connection_7__2__22_, connection_7__2__21_, 
        connection_7__2__20_, connection_7__2__19_, connection_7__2__18_, 
        connection_7__2__17_, connection_7__2__16_, connection_7__2__15_, 
        connection_7__2__14_, connection_7__2__13_, connection_7__2__12_, 
        connection_7__2__11_, connection_7__2__10_, connection_7__2__9_, 
        connection_7__2__8_, connection_7__2__7_, connection_7__2__6_, 
        connection_7__2__5_, connection_7__2__4_, connection_7__2__3_, 
        connection_7__2__2_, connection_7__2__1_, connection_7__2__0_}), 
        .o_valid({n1611, n1612}), .o_data_bus({n2449, n2450, n2451, n2452, 
        n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, 
        n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, 
        n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, 
        n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, 
        n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, 
        n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512}), 
        .i_en(i_en), .i_cmd(cmd_pipeline_stage_7__pipeline_i_cmd_reg[27:26])
         );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_13 second_half_stages_7__group_sec_half_0__switch_sec_half_3__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_7__19_, 
        connection_valid_7__3_}), .i_data_bus({connection_7__19__31_, 
        connection_7__19__30_, connection_7__19__29_, connection_7__19__28_, 
        connection_7__19__27_, connection_7__19__26_, connection_7__19__25_, 
        connection_7__19__24_, connection_7__19__23_, connection_7__19__22_, 
        connection_7__19__21_, connection_7__19__20_, connection_7__19__19_, 
        connection_7__19__18_, connection_7__19__17_, connection_7__19__16_, 
        connection_7__19__15_, connection_7__19__14_, connection_7__19__13_, 
        connection_7__19__12_, connection_7__19__11_, connection_7__19__10_, 
        connection_7__19__9_, connection_7__19__8_, connection_7__19__7_, 
        connection_7__19__6_, connection_7__19__5_, connection_7__19__4_, 
        connection_7__19__3_, connection_7__19__2_, connection_7__19__1_, 
        connection_7__19__0_, connection_7__3__31_, connection_7__3__30_, 
        connection_7__3__29_, connection_7__3__28_, connection_7__3__27_, 
        connection_7__3__26_, connection_7__3__25_, connection_7__3__24_, 
        connection_7__3__23_, connection_7__3__22_, connection_7__3__21_, 
        connection_7__3__20_, connection_7__3__19_, connection_7__3__18_, 
        connection_7__3__17_, connection_7__3__16_, connection_7__3__15_, 
        connection_7__3__14_, connection_7__3__13_, connection_7__3__12_, 
        connection_7__3__11_, connection_7__3__10_, connection_7__3__9_, 
        connection_7__3__8_, connection_7__3__7_, connection_7__3__6_, 
        connection_7__3__5_, connection_7__3__4_, connection_7__3__3_, 
        connection_7__3__2_, connection_7__3__1_, connection_7__3__0_}), 
        .o_valid({n1609, n1610}), .o_data_bus({n2385, n2386, n2387, n2388, 
        n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, 
        n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, 
        n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, 
        n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, 
        n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, 
        n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448}), 
        .i_en(i_en), .i_cmd(cmd_pipeline_stage_7__pipeline_i_cmd_reg[25:24])
         );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_12 second_half_stages_7__group_sec_half_0__switch_sec_half_4__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_7__20_, 
        connection_valid_7__4_}), .i_data_bus({connection_7__20__31_, 
        connection_7__20__30_, connection_7__20__29_, connection_7__20__28_, 
        connection_7__20__27_, connection_7__20__26_, connection_7__20__25_, 
        connection_7__20__24_, connection_7__20__23_, connection_7__20__22_, 
        connection_7__20__21_, connection_7__20__20_, connection_7__20__19_, 
        connection_7__20__18_, connection_7__20__17_, connection_7__20__16_, 
        connection_7__20__15_, connection_7__20__14_, connection_7__20__13_, 
        connection_7__20__12_, connection_7__20__11_, connection_7__20__10_, 
        connection_7__20__9_, connection_7__20__8_, connection_7__20__7_, 
        connection_7__20__6_, connection_7__20__5_, connection_7__20__4_, 
        connection_7__20__3_, connection_7__20__2_, connection_7__20__1_, 
        connection_7__20__0_, connection_7__4__31_, connection_7__4__30_, 
        connection_7__4__29_, connection_7__4__28_, connection_7__4__27_, 
        connection_7__4__26_, connection_7__4__25_, connection_7__4__24_, 
        connection_7__4__23_, connection_7__4__22_, connection_7__4__21_, 
        connection_7__4__20_, connection_7__4__19_, connection_7__4__18_, 
        connection_7__4__17_, connection_7__4__16_, connection_7__4__15_, 
        connection_7__4__14_, connection_7__4__13_, connection_7__4__12_, 
        connection_7__4__11_, connection_7__4__10_, connection_7__4__9_, 
        connection_7__4__8_, connection_7__4__7_, connection_7__4__6_, 
        connection_7__4__5_, connection_7__4__4_, connection_7__4__3_, 
        connection_7__4__2_, connection_7__4__1_, connection_7__4__0_}), 
        .o_valid({n1607, n1608}), .o_data_bus({n2321, n2322, n2323, n2324, 
        n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, 
        n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, 
        n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, 
        n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, 
        n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, 
        n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384}), 
        .i_en(i_en), .i_cmd(cmd_pipeline_stage_7__pipeline_i_cmd_reg[23:22])
         );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_11 second_half_stages_7__group_sec_half_0__switch_sec_half_5__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_7__21_, 
        connection_valid_7__5_}), .i_data_bus({connection_7__21__31_, 
        connection_7__21__30_, connection_7__21__29_, connection_7__21__28_, 
        connection_7__21__27_, connection_7__21__26_, connection_7__21__25_, 
        connection_7__21__24_, connection_7__21__23_, connection_7__21__22_, 
        connection_7__21__21_, connection_7__21__20_, connection_7__21__19_, 
        connection_7__21__18_, connection_7__21__17_, connection_7__21__16_, 
        connection_7__21__15_, connection_7__21__14_, connection_7__21__13_, 
        connection_7__21__12_, connection_7__21__11_, connection_7__21__10_, 
        connection_7__21__9_, connection_7__21__8_, connection_7__21__7_, 
        connection_7__21__6_, connection_7__21__5_, connection_7__21__4_, 
        connection_7__21__3_, connection_7__21__2_, connection_7__21__1_, 
        connection_7__21__0_, connection_7__5__31_, connection_7__5__30_, 
        connection_7__5__29_, connection_7__5__28_, connection_7__5__27_, 
        connection_7__5__26_, connection_7__5__25_, connection_7__5__24_, 
        connection_7__5__23_, connection_7__5__22_, connection_7__5__21_, 
        connection_7__5__20_, connection_7__5__19_, connection_7__5__18_, 
        connection_7__5__17_, connection_7__5__16_, connection_7__5__15_, 
        connection_7__5__14_, connection_7__5__13_, connection_7__5__12_, 
        connection_7__5__11_, connection_7__5__10_, connection_7__5__9_, 
        connection_7__5__8_, connection_7__5__7_, connection_7__5__6_, 
        connection_7__5__5_, connection_7__5__4_, connection_7__5__3_, 
        connection_7__5__2_, connection_7__5__1_, connection_7__5__0_}), 
        .o_valid({n1605, n1606}), .o_data_bus({n2257, n2258, n2259, n2260, 
        n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, 
        n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, 
        n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, 
        n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, 
        n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, 
        n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320}), 
        .i_en(i_en), .i_cmd(cmd_pipeline_stage_7__pipeline_i_cmd_reg[21:20])
         );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_10 second_half_stages_7__group_sec_half_0__switch_sec_half_6__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_7__22_, 
        connection_valid_7__6_}), .i_data_bus({connection_7__22__31_, 
        connection_7__22__30_, connection_7__22__29_, connection_7__22__28_, 
        connection_7__22__27_, connection_7__22__26_, connection_7__22__25_, 
        connection_7__22__24_, connection_7__22__23_, connection_7__22__22_, 
        connection_7__22__21_, connection_7__22__20_, connection_7__22__19_, 
        connection_7__22__18_, connection_7__22__17_, connection_7__22__16_, 
        connection_7__22__15_, connection_7__22__14_, connection_7__22__13_, 
        connection_7__22__12_, connection_7__22__11_, connection_7__22__10_, 
        connection_7__22__9_, connection_7__22__8_, connection_7__22__7_, 
        connection_7__22__6_, connection_7__22__5_, connection_7__22__4_, 
        connection_7__22__3_, connection_7__22__2_, connection_7__22__1_, 
        connection_7__22__0_, connection_7__6__31_, connection_7__6__30_, 
        connection_7__6__29_, connection_7__6__28_, connection_7__6__27_, 
        connection_7__6__26_, connection_7__6__25_, connection_7__6__24_, 
        connection_7__6__23_, connection_7__6__22_, connection_7__6__21_, 
        connection_7__6__20_, connection_7__6__19_, connection_7__6__18_, 
        connection_7__6__17_, connection_7__6__16_, connection_7__6__15_, 
        connection_7__6__14_, connection_7__6__13_, connection_7__6__12_, 
        connection_7__6__11_, connection_7__6__10_, connection_7__6__9_, 
        connection_7__6__8_, connection_7__6__7_, connection_7__6__6_, 
        connection_7__6__5_, connection_7__6__4_, connection_7__6__3_, 
        connection_7__6__2_, connection_7__6__1_, connection_7__6__0_}), 
        .o_valid({n1603, n1604}), .o_data_bus({n2193, n2194, n2195, n2196, 
        n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, 
        n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, 
        n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, 
        n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, 
        n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, 
        n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256}), 
        .i_en(i_en), .i_cmd(cmd_pipeline_stage_7__pipeline_i_cmd_reg[19:18])
         );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_9 second_half_stages_7__group_sec_half_0__switch_sec_half_7__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_7__23_, 
        connection_valid_7__7_}), .i_data_bus({connection_7__23__31_, 
        connection_7__23__30_, connection_7__23__29_, connection_7__23__28_, 
        connection_7__23__27_, connection_7__23__26_, connection_7__23__25_, 
        connection_7__23__24_, connection_7__23__23_, connection_7__23__22_, 
        connection_7__23__21_, connection_7__23__20_, connection_7__23__19_, 
        connection_7__23__18_, connection_7__23__17_, connection_7__23__16_, 
        connection_7__23__15_, connection_7__23__14_, connection_7__23__13_, 
        connection_7__23__12_, connection_7__23__11_, connection_7__23__10_, 
        connection_7__23__9_, connection_7__23__8_, connection_7__23__7_, 
        connection_7__23__6_, connection_7__23__5_, connection_7__23__4_, 
        connection_7__23__3_, connection_7__23__2_, connection_7__23__1_, 
        connection_7__23__0_, connection_7__7__31_, connection_7__7__30_, 
        connection_7__7__29_, connection_7__7__28_, connection_7__7__27_, 
        connection_7__7__26_, connection_7__7__25_, connection_7__7__24_, 
        connection_7__7__23_, connection_7__7__22_, connection_7__7__21_, 
        connection_7__7__20_, connection_7__7__19_, connection_7__7__18_, 
        connection_7__7__17_, connection_7__7__16_, connection_7__7__15_, 
        connection_7__7__14_, connection_7__7__13_, connection_7__7__12_, 
        connection_7__7__11_, connection_7__7__10_, connection_7__7__9_, 
        connection_7__7__8_, connection_7__7__7_, connection_7__7__6_, 
        connection_7__7__5_, connection_7__7__4_, connection_7__7__3_, 
        connection_7__7__2_, connection_7__7__1_, connection_7__7__0_}), 
        .o_valid({n1601, n1602}), .o_data_bus({n2129, n2130, n2131, n2132, 
        n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, 
        n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, 
        n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, 
        n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, 
        n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, 
        n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192}), 
        .i_en(i_en), .i_cmd(cmd_pipeline_stage_7__pipeline_i_cmd_reg[17:16])
         );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_8 second_half_stages_7__group_sec_half_0__switch_sec_half_8__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_7__24_, 
        connection_valid_7__8_}), .i_data_bus({connection_7__24__31_, 
        connection_7__24__30_, connection_7__24__29_, connection_7__24__28_, 
        connection_7__24__27_, connection_7__24__26_, connection_7__24__25_, 
        connection_7__24__24_, connection_7__24__23_, connection_7__24__22_, 
        connection_7__24__21_, connection_7__24__20_, connection_7__24__19_, 
        connection_7__24__18_, connection_7__24__17_, connection_7__24__16_, 
        connection_7__24__15_, connection_7__24__14_, connection_7__24__13_, 
        connection_7__24__12_, connection_7__24__11_, connection_7__24__10_, 
        connection_7__24__9_, connection_7__24__8_, connection_7__24__7_, 
        connection_7__24__6_, connection_7__24__5_, connection_7__24__4_, 
        connection_7__24__3_, connection_7__24__2_, connection_7__24__1_, 
        connection_7__24__0_, connection_7__8__31_, connection_7__8__30_, 
        connection_7__8__29_, connection_7__8__28_, connection_7__8__27_, 
        connection_7__8__26_, connection_7__8__25_, connection_7__8__24_, 
        connection_7__8__23_, connection_7__8__22_, connection_7__8__21_, 
        connection_7__8__20_, connection_7__8__19_, connection_7__8__18_, 
        connection_7__8__17_, connection_7__8__16_, connection_7__8__15_, 
        connection_7__8__14_, connection_7__8__13_, connection_7__8__12_, 
        connection_7__8__11_, connection_7__8__10_, connection_7__8__9_, 
        connection_7__8__8_, connection_7__8__7_, connection_7__8__6_, 
        connection_7__8__5_, connection_7__8__4_, connection_7__8__3_, 
        connection_7__8__2_, connection_7__8__1_, connection_7__8__0_}), 
        .o_valid({n1599, n1600}), .o_data_bus({n2065, n2066, n2067, n2068, 
        n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, 
        n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, 
        n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, 
        n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, 
        n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, 
        n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128}), 
        .i_en(i_en), .i_cmd(cmd_pipeline_stage_7__pipeline_i_cmd_reg[15:14])
         );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_7 second_half_stages_7__group_sec_half_0__switch_sec_half_9__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_7__25_, 
        connection_valid_7__9_}), .i_data_bus({connection_7__25__31_, 
        connection_7__25__30_, connection_7__25__29_, connection_7__25__28_, 
        connection_7__25__27_, connection_7__25__26_, connection_7__25__25_, 
        connection_7__25__24_, connection_7__25__23_, connection_7__25__22_, 
        connection_7__25__21_, connection_7__25__20_, connection_7__25__19_, 
        connection_7__25__18_, connection_7__25__17_, connection_7__25__16_, 
        connection_7__25__15_, connection_7__25__14_, connection_7__25__13_, 
        connection_7__25__12_, connection_7__25__11_, connection_7__25__10_, 
        connection_7__25__9_, connection_7__25__8_, connection_7__25__7_, 
        connection_7__25__6_, connection_7__25__5_, connection_7__25__4_, 
        connection_7__25__3_, connection_7__25__2_, connection_7__25__1_, 
        connection_7__25__0_, connection_7__9__31_, connection_7__9__30_, 
        connection_7__9__29_, connection_7__9__28_, connection_7__9__27_, 
        connection_7__9__26_, connection_7__9__25_, connection_7__9__24_, 
        connection_7__9__23_, connection_7__9__22_, connection_7__9__21_, 
        connection_7__9__20_, connection_7__9__19_, connection_7__9__18_, 
        connection_7__9__17_, connection_7__9__16_, connection_7__9__15_, 
        connection_7__9__14_, connection_7__9__13_, connection_7__9__12_, 
        connection_7__9__11_, connection_7__9__10_, connection_7__9__9_, 
        connection_7__9__8_, connection_7__9__7_, connection_7__9__6_, 
        connection_7__9__5_, connection_7__9__4_, connection_7__9__3_, 
        connection_7__9__2_, connection_7__9__1_, connection_7__9__0_}), 
        .o_valid({n1597, n1598}), .o_data_bus({n2001, n2002, n2003, n2004, 
        n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, 
        n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, 
        n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, 
        n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, 
        n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, 
        n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064}), 
        .i_en(i_en), .i_cmd(cmd_pipeline_stage_7__pipeline_i_cmd_reg[13:12])
         );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_6 second_half_stages_7__group_sec_half_0__switch_sec_half_10__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_7__26_, 
        connection_valid_7__10_}), .i_data_bus({connection_7__26__31_, 
        connection_7__26__30_, connection_7__26__29_, connection_7__26__28_, 
        connection_7__26__27_, connection_7__26__26_, connection_7__26__25_, 
        connection_7__26__24_, connection_7__26__23_, connection_7__26__22_, 
        connection_7__26__21_, connection_7__26__20_, connection_7__26__19_, 
        connection_7__26__18_, connection_7__26__17_, connection_7__26__16_, 
        connection_7__26__15_, connection_7__26__14_, connection_7__26__13_, 
        connection_7__26__12_, connection_7__26__11_, connection_7__26__10_, 
        connection_7__26__9_, connection_7__26__8_, connection_7__26__7_, 
        connection_7__26__6_, connection_7__26__5_, connection_7__26__4_, 
        connection_7__26__3_, connection_7__26__2_, connection_7__26__1_, 
        connection_7__26__0_, connection_7__10__31_, connection_7__10__30_, 
        connection_7__10__29_, connection_7__10__28_, connection_7__10__27_, 
        connection_7__10__26_, connection_7__10__25_, connection_7__10__24_, 
        connection_7__10__23_, connection_7__10__22_, connection_7__10__21_, 
        connection_7__10__20_, connection_7__10__19_, connection_7__10__18_, 
        connection_7__10__17_, connection_7__10__16_, connection_7__10__15_, 
        connection_7__10__14_, connection_7__10__13_, connection_7__10__12_, 
        connection_7__10__11_, connection_7__10__10_, connection_7__10__9_, 
        connection_7__10__8_, connection_7__10__7_, connection_7__10__6_, 
        connection_7__10__5_, connection_7__10__4_, connection_7__10__3_, 
        connection_7__10__2_, connection_7__10__1_, connection_7__10__0_}), 
        .o_valid({n1595, n1596}), .o_data_bus({n1937, n1938, n1939, n1940, 
        n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, 
        n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, 
        n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, 
        n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, 
        n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, 
        n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000}), 
        .i_en(i_en), .i_cmd(cmd_pipeline_stage_7__pipeline_i_cmd_reg[11:10])
         );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_5 second_half_stages_7__group_sec_half_0__switch_sec_half_11__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_7__27_, 
        connection_valid_7__11_}), .i_data_bus({connection_7__27__31_, 
        connection_7__27__30_, connection_7__27__29_, connection_7__27__28_, 
        connection_7__27__27_, connection_7__27__26_, connection_7__27__25_, 
        connection_7__27__24_, connection_7__27__23_, connection_7__27__22_, 
        connection_7__27__21_, connection_7__27__20_, connection_7__27__19_, 
        connection_7__27__18_, connection_7__27__17_, connection_7__27__16_, 
        connection_7__27__15_, connection_7__27__14_, connection_7__27__13_, 
        connection_7__27__12_, connection_7__27__11_, connection_7__27__10_, 
        connection_7__27__9_, connection_7__27__8_, connection_7__27__7_, 
        connection_7__27__6_, connection_7__27__5_, connection_7__27__4_, 
        connection_7__27__3_, connection_7__27__2_, connection_7__27__1_, 
        connection_7__27__0_, connection_7__11__31_, connection_7__11__30_, 
        connection_7__11__29_, connection_7__11__28_, connection_7__11__27_, 
        connection_7__11__26_, connection_7__11__25_, connection_7__11__24_, 
        connection_7__11__23_, connection_7__11__22_, connection_7__11__21_, 
        connection_7__11__20_, connection_7__11__19_, connection_7__11__18_, 
        connection_7__11__17_, connection_7__11__16_, connection_7__11__15_, 
        connection_7__11__14_, connection_7__11__13_, connection_7__11__12_, 
        connection_7__11__11_, connection_7__11__10_, connection_7__11__9_, 
        connection_7__11__8_, connection_7__11__7_, connection_7__11__6_, 
        connection_7__11__5_, connection_7__11__4_, connection_7__11__3_, 
        connection_7__11__2_, connection_7__11__1_, connection_7__11__0_}), 
        .o_valid({n1593, n1594}), .o_data_bus({n1873, n1874, n1875, n1876, 
        n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, 
        n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, 
        n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, 
        n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, 
        n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, 
        n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936}), 
        .i_en(i_en), .i_cmd(cmd_pipeline_stage_7__pipeline_i_cmd_reg[9:8]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_4 second_half_stages_7__group_sec_half_0__switch_sec_half_12__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_7__28_, 
        connection_valid_7__12_}), .i_data_bus({connection_7__28__31_, 
        connection_7__28__30_, connection_7__28__29_, connection_7__28__28_, 
        connection_7__28__27_, connection_7__28__26_, connection_7__28__25_, 
        connection_7__28__24_, connection_7__28__23_, connection_7__28__22_, 
        connection_7__28__21_, connection_7__28__20_, connection_7__28__19_, 
        connection_7__28__18_, connection_7__28__17_, connection_7__28__16_, 
        connection_7__28__15_, connection_7__28__14_, connection_7__28__13_, 
        connection_7__28__12_, connection_7__28__11_, connection_7__28__10_, 
        connection_7__28__9_, connection_7__28__8_, connection_7__28__7_, 
        connection_7__28__6_, connection_7__28__5_, connection_7__28__4_, 
        connection_7__28__3_, connection_7__28__2_, connection_7__28__1_, 
        connection_7__28__0_, connection_7__12__31_, connection_7__12__30_, 
        connection_7__12__29_, connection_7__12__28_, connection_7__12__27_, 
        connection_7__12__26_, connection_7__12__25_, connection_7__12__24_, 
        connection_7__12__23_, connection_7__12__22_, connection_7__12__21_, 
        connection_7__12__20_, connection_7__12__19_, connection_7__12__18_, 
        connection_7__12__17_, connection_7__12__16_, connection_7__12__15_, 
        connection_7__12__14_, connection_7__12__13_, connection_7__12__12_, 
        connection_7__12__11_, connection_7__12__10_, connection_7__12__9_, 
        connection_7__12__8_, connection_7__12__7_, connection_7__12__6_, 
        connection_7__12__5_, connection_7__12__4_, connection_7__12__3_, 
        connection_7__12__2_, connection_7__12__1_, connection_7__12__0_}), 
        .o_valid({n1591, n1592}), .o_data_bus({n1809, n1810, n1811, n1812, 
        n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, 
        n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, 
        n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, 
        n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, 
        n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, 
        n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872}), 
        .i_en(i_en), .i_cmd(cmd_pipeline_stage_7__pipeline_i_cmd_reg[7:6]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_3 second_half_stages_7__group_sec_half_0__switch_sec_half_13__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_7__29_, 
        connection_valid_7__13_}), .i_data_bus({connection_7__29__31_, 
        connection_7__29__30_, connection_7__29__29_, connection_7__29__28_, 
        connection_7__29__27_, connection_7__29__26_, connection_7__29__25_, 
        connection_7__29__24_, connection_7__29__23_, connection_7__29__22_, 
        connection_7__29__21_, connection_7__29__20_, connection_7__29__19_, 
        connection_7__29__18_, connection_7__29__17_, connection_7__29__16_, 
        connection_7__29__15_, connection_7__29__14_, connection_7__29__13_, 
        connection_7__29__12_, connection_7__29__11_, connection_7__29__10_, 
        connection_7__29__9_, connection_7__29__8_, connection_7__29__7_, 
        connection_7__29__6_, connection_7__29__5_, connection_7__29__4_, 
        connection_7__29__3_, connection_7__29__2_, connection_7__29__1_, 
        connection_7__29__0_, connection_7__13__31_, connection_7__13__30_, 
        connection_7__13__29_, connection_7__13__28_, connection_7__13__27_, 
        connection_7__13__26_, connection_7__13__25_, connection_7__13__24_, 
        connection_7__13__23_, connection_7__13__22_, connection_7__13__21_, 
        connection_7__13__20_, connection_7__13__19_, connection_7__13__18_, 
        connection_7__13__17_, connection_7__13__16_, connection_7__13__15_, 
        connection_7__13__14_, connection_7__13__13_, connection_7__13__12_, 
        connection_7__13__11_, connection_7__13__10_, connection_7__13__9_, 
        connection_7__13__8_, connection_7__13__7_, connection_7__13__6_, 
        connection_7__13__5_, connection_7__13__4_, connection_7__13__3_, 
        connection_7__13__2_, connection_7__13__1_, connection_7__13__0_}), 
        .o_valid({n1589, n1590}), .o_data_bus({n1745, n1746, n1747, n1748, 
        n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, 
        n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, 
        n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, 
        n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, 
        n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, 
        n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808}), 
        .i_en(i_en), .i_cmd(cmd_pipeline_stage_7__pipeline_i_cmd_reg[5:4]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_2 second_half_stages_7__group_sec_half_0__switch_sec_half_14__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_7__30_, 
        connection_valid_7__14_}), .i_data_bus({connection_7__30__31_, 
        connection_7__30__30_, connection_7__30__29_, connection_7__30__28_, 
        connection_7__30__27_, connection_7__30__26_, connection_7__30__25_, 
        connection_7__30__24_, connection_7__30__23_, connection_7__30__22_, 
        connection_7__30__21_, connection_7__30__20_, connection_7__30__19_, 
        connection_7__30__18_, connection_7__30__17_, connection_7__30__16_, 
        connection_7__30__15_, connection_7__30__14_, connection_7__30__13_, 
        connection_7__30__12_, connection_7__30__11_, connection_7__30__10_, 
        connection_7__30__9_, connection_7__30__8_, connection_7__30__7_, 
        connection_7__30__6_, connection_7__30__5_, connection_7__30__4_, 
        connection_7__30__3_, connection_7__30__2_, connection_7__30__1_, 
        connection_7__30__0_, connection_7__14__31_, connection_7__14__30_, 
        connection_7__14__29_, connection_7__14__28_, connection_7__14__27_, 
        connection_7__14__26_, connection_7__14__25_, connection_7__14__24_, 
        connection_7__14__23_, connection_7__14__22_, connection_7__14__21_, 
        connection_7__14__20_, connection_7__14__19_, connection_7__14__18_, 
        connection_7__14__17_, connection_7__14__16_, connection_7__14__15_, 
        connection_7__14__14_, connection_7__14__13_, connection_7__14__12_, 
        connection_7__14__11_, connection_7__14__10_, connection_7__14__9_, 
        connection_7__14__8_, connection_7__14__7_, connection_7__14__6_, 
        connection_7__14__5_, connection_7__14__4_, connection_7__14__3_, 
        connection_7__14__2_, connection_7__14__1_, connection_7__14__0_}), 
        .o_valid({n1587, n1588}), .o_data_bus({n1681, n1682, n1683, n1684, 
        n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, 
        n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, 
        n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, 
        n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, 
        n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, 
        n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744}), 
        .i_en(i_en), .i_cmd(cmd_pipeline_stage_7__pipeline_i_cmd_reg[3:2]) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_1 second_half_stages_7__group_sec_half_0__switch_sec_half_15__third_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_7__31_, 
        connection_valid_7__15_}), .i_data_bus({connection_7__31__31_, 
        connection_7__31__30_, connection_7__31__29_, connection_7__31__28_, 
        connection_7__31__27_, connection_7__31__26_, connection_7__31__25_, 
        connection_7__31__24_, connection_7__31__23_, connection_7__31__22_, 
        connection_7__31__21_, connection_7__31__20_, connection_7__31__19_, 
        connection_7__31__18_, connection_7__31__17_, connection_7__31__16_, 
        connection_7__31__15_, connection_7__31__14_, connection_7__31__13_, 
        connection_7__31__12_, connection_7__31__11_, connection_7__31__10_, 
        connection_7__31__9_, connection_7__31__8_, connection_7__31__7_, 
        connection_7__31__6_, connection_7__31__5_, connection_7__31__4_, 
        connection_7__31__3_, connection_7__31__2_, connection_7__31__1_, 
        connection_7__31__0_, connection_7__15__31_, connection_7__15__30_, 
        connection_7__15__29_, connection_7__15__28_, connection_7__15__27_, 
        connection_7__15__26_, connection_7__15__25_, connection_7__15__24_, 
        connection_7__15__23_, connection_7__15__22_, connection_7__15__21_, 
        connection_7__15__20_, connection_7__15__19_, connection_7__15__18_, 
        connection_7__15__17_, connection_7__15__16_, connection_7__15__15_, 
        connection_7__15__14_, connection_7__15__13_, connection_7__15__12_, 
        connection_7__15__11_, connection_7__15__10_, connection_7__15__9_, 
        connection_7__15__8_, connection_7__15__7_, connection_7__15__6_, 
        connection_7__15__5_, connection_7__15__4_, connection_7__15__3_, 
        connection_7__15__2_, connection_7__15__1_, connection_7__15__0_}), 
        .o_valid({n1585, n1586}), .o_data_bus({n1617, n1618, n1619, n1620, 
        n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, 
        n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, 
        n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, 
        n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, 
        n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, 
        n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680}), 
        .i_en(i_en), .i_cmd(cmd_pipeline_stage_7__pipeline_i_cmd_reg[1:0]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__0__1_ ( .D(
        i_cmd[65]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[223]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__0__0_ ( .D(
        i_cmd[64]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[222]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__1__1_ ( .D(
        i_cmd[67]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[221]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__1__0_ ( .D(
        i_cmd[66]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[220]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__2__1_ ( .D(
        i_cmd[69]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[219]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__2__0_ ( .D(
        i_cmd[68]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[218]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__3__1_ ( .D(
        i_cmd[71]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[217]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__3__0_ ( .D(
        i_cmd[70]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[216]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__4__1_ ( .D(
        i_cmd[73]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[215]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__4__0_ ( .D(
        i_cmd[72]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[214]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__5__1_ ( .D(
        i_cmd[75]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[213]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__5__0_ ( .D(
        i_cmd[74]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[212]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__6__1_ ( .D(
        i_cmd[77]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[211]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__6__0_ ( .D(
        i_cmd[76]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[210]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__7__1_ ( .D(
        i_cmd[79]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[209]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__7__0_ ( .D(
        i_cmd[78]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[208]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__8__1_ ( .D(
        i_cmd[81]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[207]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__8__0_ ( .D(
        i_cmd[80]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[206]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__9__1_ ( .D(
        i_cmd[83]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[205]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__9__0_ ( .D(
        i_cmd[82]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[204]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__10__1_ ( .D(
        i_cmd[85]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[203]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__10__0_ ( .D(
        i_cmd[84]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[202]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__11__1_ ( .D(
        i_cmd[87]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[201]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__11__0_ ( .D(
        i_cmd[86]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[200]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__12__1_ ( .D(
        i_cmd[89]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[199]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__12__0_ ( .D(
        i_cmd[88]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[198]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__13__1_ ( .D(
        i_cmd[91]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[197]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__13__0_ ( .D(
        i_cmd[90]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[196]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__14__1_ ( .D(
        i_cmd[93]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[195]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__14__0_ ( .D(
        i_cmd[92]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[194]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__15__1_ ( .D(
        i_cmd[95]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[193]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__15__0_ ( .D(
        i_cmd[94]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[192]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__0__1_ ( .D(
        i_cmd[97]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[191]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__0__0_ ( .D(
        i_cmd[96]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[190]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__1__1_ ( .D(
        i_cmd[99]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[189]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__1__0_ ( .D(
        i_cmd[98]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[188]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__2__1_ ( .D(
        i_cmd[101]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[187]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__2__0_ ( .D(
        i_cmd[100]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[186]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__3__1_ ( .D(
        i_cmd[103]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[185]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__3__0_ ( .D(
        i_cmd[102]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[184]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__4__1_ ( .D(
        i_cmd[105]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[183]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__4__0_ ( .D(
        i_cmd[104]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[182]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__5__1_ ( .D(
        i_cmd[107]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[181]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__5__0_ ( .D(
        i_cmd[106]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[180]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__6__1_ ( .D(
        i_cmd[109]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[179]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__6__0_ ( .D(
        i_cmd[108]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[178]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__7__1_ ( .D(
        i_cmd[111]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[177]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__7__0_ ( .D(
        i_cmd[110]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[176]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__8__1_ ( .D(
        i_cmd[113]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[175]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__8__0_ ( .D(
        i_cmd[112]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[174]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__9__1_ ( .D(
        i_cmd[115]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[173]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__9__0_ ( .D(
        i_cmd[114]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[172]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__10__1_ ( .D(
        i_cmd[117]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[171]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__10__0_ ( .D(
        i_cmd[116]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[170]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__11__1_ ( .D(
        i_cmd[119]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[169]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__11__0_ ( .D(
        i_cmd[118]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[168]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__12__1_ ( .D(
        i_cmd[121]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[167]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__12__0_ ( .D(
        i_cmd[120]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[166]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__13__1_ ( .D(
        i_cmd[123]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[165]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__13__0_ ( .D(
        i_cmd[122]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[164]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__14__1_ ( .D(
        i_cmd[125]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[163]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__14__0_ ( .D(
        i_cmd[124]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[162]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__15__1_ ( .D(
        i_cmd[127]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[161]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__15__0_ ( .D(
        i_cmd[126]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[160]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__0__1_ ( .D(
        i_cmd[129]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[159]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__0__0_ ( .D(
        i_cmd[128]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[158]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__1__1_ ( .D(
        i_cmd[131]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[157]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__1__0_ ( .D(
        i_cmd[130]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[156]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__2__1_ ( .D(
        i_cmd[133]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[155]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__2__0_ ( .D(
        i_cmd[132]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[154]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__3__1_ ( .D(
        i_cmd[135]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[153]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__3__0_ ( .D(
        i_cmd[134]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[152]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__4__1_ ( .D(
        i_cmd[137]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[151]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__4__0_ ( .D(
        i_cmd[136]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[150]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__5__1_ ( .D(
        i_cmd[139]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[149]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__5__0_ ( .D(
        i_cmd[138]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[148]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__6__1_ ( .D(
        i_cmd[141]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[147]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__6__0_ ( .D(
        i_cmd[140]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[146]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__7__1_ ( .D(
        i_cmd[143]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[145]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__7__0_ ( .D(
        i_cmd[142]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[144]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__8__1_ ( .D(
        i_cmd[145]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[143]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__8__0_ ( .D(
        i_cmd[144]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[142]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__9__1_ ( .D(
        i_cmd[147]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[141]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__9__0_ ( .D(
        i_cmd[146]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[140]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__10__1_ ( .D(
        i_cmd[149]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[139]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__10__0_ ( .D(
        i_cmd[148]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[138]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__11__1_ ( .D(
        i_cmd[151]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[137]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__11__0_ ( .D(
        i_cmd[150]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[136]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__12__1_ ( .D(
        i_cmd[153]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[135]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__12__0_ ( .D(
        i_cmd[152]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[134]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__13__1_ ( .D(
        i_cmd[155]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[133]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__13__0_ ( .D(
        i_cmd[154]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[132]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__14__1_ ( .D(
        i_cmd[157]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[131]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__14__0_ ( .D(
        i_cmd[156]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[130]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__15__1_ ( .D(
        i_cmd[159]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[129]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__15__0_ ( .D(
        i_cmd[158]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[128]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__0__1_ ( .D(
        i_cmd[161]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[127]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__0__0_ ( .D(
        i_cmd[160]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[126]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__1__1_ ( .D(
        i_cmd[163]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[125]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__1__0_ ( .D(
        i_cmd[162]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[124]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__2__1_ ( .D(
        i_cmd[165]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[123]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__2__0_ ( .D(
        i_cmd[164]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[122]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__3__1_ ( .D(
        i_cmd[167]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[121]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__3__0_ ( .D(
        i_cmd[166]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[120]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__4__1_ ( .D(
        i_cmd[169]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[119]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__4__0_ ( .D(
        i_cmd[168]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[118]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__5__1_ ( .D(
        i_cmd[171]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[117]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__5__0_ ( .D(
        i_cmd[170]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[116]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__6__1_ ( .D(
        i_cmd[173]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[115]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__6__0_ ( .D(
        i_cmd[172]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[114]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__7__1_ ( .D(
        i_cmd[175]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[113]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__7__0_ ( .D(
        i_cmd[174]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[112]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__8__1_ ( .D(
        i_cmd[177]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[111]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__8__0_ ( .D(
        i_cmd[176]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[110]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__9__1_ ( .D(
        i_cmd[179]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[109]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__9__0_ ( .D(
        i_cmd[178]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[108]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__10__1_ ( .D(
        i_cmd[181]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[107]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__10__0_ ( .D(
        i_cmd[180]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[106]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__11__1_ ( .D(
        i_cmd[183]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[105]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__11__0_ ( .D(
        i_cmd[182]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[104]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__12__1_ ( .D(
        i_cmd[185]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[103]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__12__0_ ( .D(
        i_cmd[184]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[102]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__13__1_ ( .D(
        i_cmd[187]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[101]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__13__0_ ( .D(
        i_cmd[186]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[100]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__14__1_ ( .D(
        i_cmd[189]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[99]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__14__0_ ( .D(
        i_cmd[188]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[98]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__15__1_ ( .D(
        i_cmd[191]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[97]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__15__0_ ( .D(
        i_cmd[190]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[96]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__0__1_ ( .D(
        i_cmd[193]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[95]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__0__0_ ( .D(
        i_cmd[192]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[94]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__1__1_ ( .D(
        i_cmd[195]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[93]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__1__0_ ( .D(
        i_cmd[194]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[92]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__2__1_ ( .D(
        i_cmd[197]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[91]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__2__0_ ( .D(
        i_cmd[196]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[90]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__3__1_ ( .D(
        i_cmd[199]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[89]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__3__0_ ( .D(
        i_cmd[198]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[88]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__4__1_ ( .D(
        i_cmd[201]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[87]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__4__0_ ( .D(
        i_cmd[200]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[86]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__5__1_ ( .D(
        i_cmd[203]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[85]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__5__0_ ( .D(
        i_cmd[202]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[84]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__6__1_ ( .D(
        i_cmd[205]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[83]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__6__0_ ( .D(
        i_cmd[204]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[82]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__7__1_ ( .D(
        i_cmd[207]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[81]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__7__0_ ( .D(
        i_cmd[206]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[80]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__8__1_ ( .D(
        i_cmd[209]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[79]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__8__0_ ( .D(
        i_cmd[208]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[78]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__9__1_ ( .D(
        i_cmd[211]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[77]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__9__0_ ( .D(
        i_cmd[210]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[76]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__10__1_ ( .D(
        i_cmd[213]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[75]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__10__0_ ( .D(
        i_cmd[212]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[74]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__11__1_ ( .D(
        i_cmd[215]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[73]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__11__0_ ( .D(
        i_cmd[214]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[72]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__12__1_ ( .D(
        i_cmd[217]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[71]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__12__0_ ( .D(
        i_cmd[216]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[70]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__13__1_ ( .D(
        i_cmd[219]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[69]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__13__0_ ( .D(
        i_cmd[218]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[68]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__14__1_ ( .D(
        i_cmd[221]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[67]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__14__0_ ( .D(
        i_cmd[220]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[66]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__15__1_ ( .D(
        i_cmd[223]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[65]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__15__0_ ( .D(
        i_cmd[222]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[64]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__0__1_ ( .D(
        i_cmd[225]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[63]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__0__0_ ( .D(
        i_cmd[224]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[62]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__1__1_ ( .D(
        i_cmd[227]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[61]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__1__0_ ( .D(
        i_cmd[226]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[60]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__2__1_ ( .D(
        i_cmd[229]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[59]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__2__0_ ( .D(
        i_cmd[228]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[58]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__3__1_ ( .D(
        i_cmd[231]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[57]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__3__0_ ( .D(
        i_cmd[230]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[56]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__4__1_ ( .D(
        i_cmd[233]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[55]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__4__0_ ( .D(
        i_cmd[232]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[54]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__5__1_ ( .D(
        i_cmd[235]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[53]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__5__0_ ( .D(
        i_cmd[234]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[52]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__6__1_ ( .D(
        i_cmd[237]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[51]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__6__0_ ( .D(
        i_cmd[236]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[50]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__7__1_ ( .D(
        i_cmd[239]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[49]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__7__0_ ( .D(
        i_cmd[238]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[48]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__8__1_ ( .D(
        i_cmd[241]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[47]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__8__0_ ( .D(
        i_cmd[240]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[46]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__9__1_ ( .D(
        i_cmd[243]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[45]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__9__0_ ( .D(
        i_cmd[242]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[44]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__10__1_ ( .D(
        i_cmd[245]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[43]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__10__0_ ( .D(
        i_cmd[244]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[42]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__11__1_ ( .D(
        i_cmd[247]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[41]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__11__0_ ( .D(
        i_cmd[246]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[40]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__12__1_ ( .D(
        i_cmd[249]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[39]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__12__0_ ( .D(
        i_cmd[248]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[38]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__13__1_ ( .D(
        i_cmd[251]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[37]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__13__0_ ( .D(
        i_cmd[250]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[36]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__14__1_ ( .D(
        i_cmd[253]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[35]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__14__0_ ( .D(
        i_cmd[252]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[34]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__15__1_ ( .D(
        i_cmd[255]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[33]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_6__15__0_ ( .D(
        i_cmd[254]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[32]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__0__1_ ( .D(
        i_cmd[257]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[31]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__0__0_ ( .D(
        i_cmd[256]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[30]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__1__1_ ( .D(
        i_cmd[259]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[29]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__1__0_ ( .D(
        i_cmd[258]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[28]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__2__1_ ( .D(
        i_cmd[261]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[27]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__2__0_ ( .D(
        i_cmd[260]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[26]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__3__1_ ( .D(
        i_cmd[263]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[25]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__3__0_ ( .D(
        i_cmd[262]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[24]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__4__1_ ( .D(
        i_cmd[265]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[23]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__4__0_ ( .D(
        i_cmd[264]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[22]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__5__1_ ( .D(
        i_cmd[267]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[21]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__5__0_ ( .D(
        i_cmd[266]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[20]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__6__1_ ( .D(
        i_cmd[269]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[19]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__6__0_ ( .D(
        i_cmd[268]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[18]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__7__1_ ( .D(
        i_cmd[271]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[17]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__7__0_ ( .D(
        i_cmd[270]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[16]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__8__1_ ( .D(
        i_cmd[273]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[15]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__8__0_ ( .D(
        i_cmd[272]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[14]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__9__1_ ( .D(
        i_cmd[275]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[13]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__9__0_ ( .D(
        i_cmd[274]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[12]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__10__1_ ( .D(
        i_cmd[277]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[11]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__10__0_ ( .D(
        i_cmd[276]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[10]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__11__1_ ( .D(
        i_cmd[279]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[9])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__11__0_ ( .D(
        i_cmd[278]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[8])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__12__1_ ( .D(
        i_cmd[281]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[7])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__12__0_ ( .D(
        i_cmd[280]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[6])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__13__1_ ( .D(
        i_cmd[283]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[5])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__13__0_ ( .D(
        i_cmd[282]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[4])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__14__1_ ( .D(
        i_cmd[285]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[3])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__14__0_ ( .D(
        i_cmd[284]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[2])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__15__1_ ( .D(
        i_cmd[287]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[1])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_7__15__0_ ( .D(
        i_cmd[286]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[0])
         );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__0__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[191]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[191]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__0__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[190]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[190]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__1__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[189]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[189]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__1__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[188]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[188]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__2__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[187]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[187]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__2__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[186]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[186]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__3__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[185]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[185]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__3__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[184]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[184]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__4__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[183]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[183]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__4__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[182]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[182]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__5__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[181]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[181]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__5__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[180]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[180]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__6__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[179]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[179]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__6__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[178]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[178]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__7__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[177]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[177]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__7__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[176]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[176]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__8__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[175]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[175]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__8__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[174]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[174]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__9__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[173]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[173]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__9__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[172]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[172]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__10__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[171]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[171]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__10__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[170]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[170]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__11__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[169]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[169]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__11__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[168]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[168]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__12__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[167]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[167]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__12__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[166]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[166]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__13__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[165]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[165]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__13__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[164]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[164]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__14__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[163]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[163]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__14__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[162]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[162]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__15__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[161]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[161]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__15__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[160]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[160]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__0__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[159]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[159]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__0__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[158]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[158]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__1__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[157]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[157]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__1__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[156]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[156]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__2__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[155]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[155]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__2__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[154]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[154]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__3__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[153]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[153]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__3__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[152]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[152]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__4__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[151]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[151]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__4__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[150]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[150]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__5__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[149]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[149]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__5__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[148]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[148]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__6__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[147]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[147]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__6__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[146]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[146]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__7__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[145]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[145]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__7__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[144]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[144]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__8__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[143]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[143]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__8__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[142]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[142]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__9__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[141]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[141]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__9__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[140]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[140]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__10__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[139]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[139]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__10__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[138]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[138]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__11__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[137]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[137]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__11__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[136]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[136]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__12__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[135]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[135]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__12__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[134]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[134]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__13__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[133]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[133]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__13__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[132]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[132]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__14__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[131]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[131]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__14__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[130]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[130]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__15__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[129]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[129]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__15__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[128]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[128]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__0__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[127]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[127]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__0__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[126]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[126]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__1__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[125]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[125]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__1__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[124]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[124]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__2__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[123]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[123]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__2__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[122]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[122]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__3__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[121]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[121]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__3__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[120]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[120]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__4__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[119]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[119]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__4__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[118]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[118]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__5__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[117]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[117]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__5__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[116]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[116]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__6__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[115]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[115]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__6__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[114]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[114]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__7__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[113]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[113]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__7__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[112]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[112]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__8__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[111]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[111]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__8__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[110]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[110]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__9__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[109]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[109]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__9__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[108]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[108]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__10__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[107]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[107]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__10__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[106]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[106]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__11__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[105]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[105]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__11__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[104]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[104]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__12__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[103]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[103]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__12__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[102]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[102]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__13__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[101]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[101]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__13__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[100]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[100]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__14__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[99]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[99]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__14__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[98]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[98]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__15__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[97]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[97]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__15__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[96]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[96]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__0__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[95]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[95]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__0__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[94]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[94]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__1__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[93]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[93]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__1__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[92]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[92]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__2__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[91]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[91]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__2__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[90]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[90]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__3__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[89]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[89]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__3__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[88]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[88]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__4__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[87]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[87]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__4__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[86]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[86]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__5__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[85]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[85]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__5__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[84]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[84]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__6__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[83]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[83]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__6__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[82]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[82]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__7__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[81]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[81]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__7__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[80]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[80]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__8__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[79]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[79]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__8__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[78]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[78]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__9__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[77]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[77]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__9__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[76]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[76]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__10__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[75]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[75]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__10__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[74]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[74]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__11__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[73]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[73]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__11__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[72]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[72]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__12__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[71]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[71]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__12__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[70]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[70]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__13__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[69]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[69]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__13__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[68]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[68]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__14__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[67]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[67]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__14__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[66]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[66]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__15__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[65]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[65]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__15__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[64]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[64]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__0__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[63]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[63]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__0__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[62]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[62]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__1__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[61]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[61]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__1__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[60]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[60]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__2__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[59]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[59]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__2__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[58]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[58]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__3__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[57]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[57]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__3__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[56]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[56]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__4__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[55]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[55]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__4__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[54]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[54]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__5__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[53]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[53]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__5__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[52]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[52]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__6__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[51]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[51]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__6__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[50]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[50]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__7__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[49]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[49]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__7__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[48]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[48]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__8__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[47]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[47]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__8__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[46]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[46]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__9__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[45]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[45]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__9__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[44]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[44]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__10__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[43]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[43]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__10__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[42]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[42]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__11__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[41]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[41]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__11__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[40]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[40]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__12__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[39]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[39]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__12__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[38]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[38]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__13__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[37]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[37]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__13__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[36]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[36]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__14__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[35]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[35]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__14__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[34]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[34]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__15__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[33]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[33]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_5__15__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[32]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[32]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__0__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[31]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[31]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__0__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[30]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[30]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__1__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[29]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[29]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__1__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[28]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[28]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__2__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[27]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[27]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__2__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[26]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[26]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__3__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[25]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[25]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__3__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[24]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[24]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__4__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[23]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[23]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__4__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[22]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[22]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__5__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[21]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[21]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__5__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[20]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[20]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__6__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[19]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[19]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__6__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[18]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[18]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__7__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[17]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[17]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__7__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[16]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[16]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__8__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[15]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[15]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__8__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[14]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[14]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__9__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[13]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[13]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__9__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[12]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[12]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__10__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[11]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[11]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__10__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[10]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[10]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__11__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[9]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[9]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__11__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[8]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[8]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__12__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[7]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[7]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__12__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[6]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[6]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__13__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[5]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[5]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__13__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[4]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[4]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__14__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[3]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[3]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__14__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[2]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[2]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__15__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[1]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[1]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_6__15__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[0]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[0]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__7__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[176]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[176]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__8__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[174]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[174]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__9__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[172]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[172]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__10__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[170]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[170]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__11__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[168]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[168]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__13__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[164]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[164]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__15__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[160]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[160]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__0__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[159]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[159]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__0__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[158]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[158]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__1__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[157]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[157]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__1__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[156]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[156]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__2__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[155]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[155]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__2__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[154]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[154]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__3__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[153]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[153]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__3__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[152]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[152]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__4__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[151]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[151]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__4__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[150]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[150]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__5__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[149]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[149]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__5__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[148]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[148]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__6__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[147]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[147]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__6__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[146]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[146]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__7__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[145]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[145]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__7__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[144]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[144]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__8__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[143]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[143]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__8__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[142]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[142]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__9__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[141]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[141]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__9__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[140]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[140]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__10__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[139]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[139]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__10__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[138]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[138]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__11__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[137]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[137]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__11__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[136]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[136]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__12__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[135]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[135]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__12__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[134]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[134]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__13__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[133]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[133]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__13__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[132]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[132]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__14__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[131]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[131]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__14__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[130]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[130]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__15__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[129]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[129]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__15__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[128]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[128]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__0__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[127]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[127]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__0__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[126]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[126]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__1__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[125]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[125]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__1__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[124]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[124]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__2__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[123]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[123]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__2__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[122]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[122]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__3__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[121]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[121]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__3__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[120]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[120]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__4__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[119]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[119]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__4__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[118]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[118]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__5__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[117]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[117]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__5__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[116]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[116]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__6__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[115]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[115]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__6__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[114]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[114]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__7__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[113]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[113]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__7__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[112]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[112]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__8__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[111]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[111]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__8__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[110]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[110]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__9__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[109]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[109]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__9__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[108]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[108]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__10__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[107]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[107]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__10__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[106]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[106]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__11__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[105]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[105]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__11__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[104]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[104]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__12__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[103]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[103]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__12__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[102]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[102]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__13__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[101]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[101]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__13__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[100]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[100]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__14__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[99]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[99]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__14__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[98]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[98]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__15__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[97]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[97]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__15__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[96]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[96]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__0__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[95]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[95]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__0__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[94]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[94]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__1__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[93]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[93]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__1__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[92]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[92]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__2__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[91]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[91]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__2__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[90]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[90]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__3__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[89]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[89]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__3__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[88]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[88]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__4__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[87]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[87]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__4__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[86]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[86]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__5__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[85]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[85]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__5__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[84]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[84]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__6__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[83]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[83]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__6__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[82]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[82]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__7__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[81]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[81]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__7__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[80]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[80]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__8__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[79]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[79]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__8__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[78]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[78]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__9__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[77]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[77]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__9__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[76]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[76]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__10__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[75]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[75]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__10__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[74]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[74]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__11__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[73]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[73]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__11__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[72]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[72]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__12__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[71]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[71]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__12__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[70]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[70]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__13__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[69]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[69]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__13__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[68]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[68]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__14__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[67]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[67]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__14__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[66]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[66]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__15__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[65]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[65]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__15__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[64]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[64]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__0__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[63]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[63]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__0__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[62]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[62]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__1__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[61]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[61]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__1__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[60]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[60]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__2__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[59]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[59]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__2__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[58]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[58]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__3__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[57]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[57]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__3__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[56]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[56]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__4__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[55]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[55]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__4__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[54]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[54]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__5__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[53]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[53]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__5__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[52]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[52]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__6__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[51]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[51]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__6__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[50]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[50]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__7__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[49]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[49]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__7__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[48]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[48]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__8__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[47]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[47]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__8__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[46]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[46]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__9__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[45]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[45]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__9__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[44]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[44]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__10__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[43]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[43]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__10__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[42]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[42]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__11__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[41]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[41]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__11__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[40]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[40]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__12__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[39]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[39]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__12__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[38]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[38]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__13__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[37]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[37]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__13__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[36]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[36]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__14__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[35]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[35]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__14__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[34]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[34]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__15__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[33]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[33]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_4__15__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[32]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[32]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__0__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[31]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[31]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__0__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[30]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[30]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__1__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[29]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[29]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__1__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[28]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[28]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__2__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[27]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[27]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__2__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[26]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[26]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__3__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[25]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[25]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__3__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[24]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[24]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__4__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[23]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[23]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__4__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[22]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[22]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__5__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[21]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[21]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__5__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[20]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[20]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__6__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[19]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[19]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__6__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[18]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[18]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__7__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[17]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[17]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__7__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[16]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[16]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__8__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[15]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[15]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__8__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[14]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[14]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__9__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[13]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[13]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__9__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[12]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[12]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__10__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[11]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[11]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__10__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[10]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[10]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__11__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[9]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[9]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__11__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[8]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[8]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__12__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[7]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[7]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__12__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[6]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[6]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__13__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[5]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[5]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__13__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[4]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[4]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__14__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[3]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[3]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__14__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[2]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[2]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__15__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[1]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[1]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_5__15__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[0]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[0]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__1__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[156]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[156]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__5__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[148]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[148]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__0__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[127]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[127]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__0__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[126]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[126]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__1__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[125]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[125]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__1__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[124]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[124]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__2__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[123]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[123]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__2__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[122]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[122]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__3__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[121]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[121]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__3__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[120]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[120]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__4__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[119]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[119]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__4__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[118]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[118]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__5__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[117]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[117]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__5__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[116]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[116]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__6__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[115]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[115]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__6__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[114]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[114]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__7__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[113]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[113]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__7__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[112]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[112]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__8__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[111]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[111]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__8__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[110]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[110]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__9__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[109]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[109]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__9__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[108]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[108]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__10__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[107]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[107]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__10__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[106]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[106]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__11__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[105]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[105]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__11__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[104]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[104]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__12__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[103]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[103]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__12__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[102]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[102]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__13__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[101]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[101]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__13__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[100]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[100]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__14__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[99]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[99]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__14__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[98]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[98]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__15__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[97]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[97]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__15__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[96]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[96]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__0__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[95]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[95]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__0__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[94]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[94]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__1__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[93]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[93]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__1__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[92]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[92]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__2__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[91]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[91]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__2__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[90]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[90]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__3__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[89]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[89]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__3__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[88]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[88]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__4__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[87]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[87]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__4__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[86]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[86]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__5__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[85]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[85]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__5__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[84]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[84]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__6__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[83]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[83]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__6__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[82]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[82]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__7__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[81]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[81]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__7__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[80]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[80]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__8__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[79]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[79]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__8__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[78]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[78]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__9__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[77]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[77]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__9__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[76]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[76]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__10__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[75]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[75]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__10__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[74]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[74]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__11__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[73]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[73]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__11__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[72]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[72]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__12__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[71]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[71]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__12__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[70]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[70]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__13__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[69]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[69]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__13__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[68]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[68]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__14__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[67]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[67]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__14__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[66]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[66]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__15__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[65]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[65]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__15__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[64]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[64]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__0__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[63]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[63]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__0__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[62]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[62]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__1__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[61]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[61]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__1__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[60]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[60]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__2__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[59]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[59]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__2__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[58]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[58]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__3__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[57]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[57]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__3__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[56]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[56]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__4__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[55]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[55]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__4__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[54]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[54]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__5__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[53]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[53]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__5__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[52]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[52]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__6__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[51]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[51]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__6__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[50]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[50]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__7__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[49]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[49]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__7__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[48]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[48]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__8__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[47]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[47]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__8__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[46]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[46]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__9__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[45]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[45]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__9__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[44]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[44]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__10__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[43]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[43]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__10__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[42]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[42]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__11__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[41]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[41]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__11__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[40]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[40]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__12__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[39]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[39]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__12__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[38]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[38]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__13__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[37]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[37]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__13__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[36]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[36]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__14__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[35]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[35]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__14__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[34]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[34]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__15__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[33]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[33]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_3__15__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[32]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[32]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__0__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[31]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[31]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__0__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[30]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[30]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__1__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[29]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[29]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__1__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[28]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[28]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__2__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[27]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[27]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__2__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[26]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[26]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__3__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[25]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[25]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__3__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[24]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[24]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__4__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[23]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[23]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__4__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[22]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[22]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__5__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[21]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[21]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__5__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[20]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[20]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__6__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[19]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[19]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__6__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[18]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[18]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__7__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[17]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[17]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__7__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[16]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[16]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__8__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[15]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[15]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__8__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[14]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[14]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__9__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[13]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[13]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__9__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[12]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[12]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__10__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[11]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[11]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__10__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[10]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[10]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__11__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[9]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[9]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__11__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[8]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[8]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__12__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[7]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[7]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__12__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[6]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[6]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__13__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[5]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[5]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__13__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[4]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[4]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__14__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[3]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[3]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__14__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[2]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[2]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__15__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[1]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[1]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_4__15__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[0]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[0]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__0__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[95]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[95]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__0__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[94]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[94]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__1__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[93]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[93]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__1__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[92]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[92]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__2__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[91]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[91]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__2__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[90]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[90]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__3__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[89]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[89]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__3__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[88]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[88]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__4__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[87]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[87]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__4__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[86]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[86]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__5__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[85]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[85]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__5__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[84]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[84]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__6__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[83]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[83]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__6__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[82]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[82]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__7__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[81]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[81]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__7__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[80]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[80]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__8__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[79]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[79]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__8__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[78]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[78]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__9__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[77]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[77]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__9__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[76]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[76]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__10__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[75]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[75]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__10__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[74]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[74]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__11__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[73]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[73]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__11__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[72]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[72]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__12__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[71]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[71]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__12__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[70]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[70]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__13__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[69]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[69]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__13__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[68]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[68]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__14__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[67]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[67]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__14__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[66]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[66]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__15__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[65]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[65]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__15__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[64]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[64]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__0__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[63]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[63]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__0__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[62]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[62]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__1__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[61]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[61]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__1__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[60]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[60]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__2__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[59]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[59]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__2__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[58]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[58]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__3__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[57]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[57]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__3__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[56]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[56]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__4__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[55]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[55]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__4__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[54]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[54]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__5__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[53]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[53]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__5__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[52]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[52]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__6__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[51]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[51]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__6__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[50]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[50]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__7__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[49]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[49]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__7__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[48]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[48]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__8__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[47]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[47]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__8__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[46]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[46]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__9__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[45]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[45]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__9__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[44]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[44]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__10__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[43]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[43]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__10__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[42]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[42]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__11__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[41]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[41]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__11__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[40]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[40]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__12__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[39]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[39]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__12__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[38]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[38]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__13__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[37]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[37]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__13__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[36]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[36]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__14__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[35]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[35]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__14__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[34]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[34]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__15__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[33]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[33]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_2__15__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[32]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[32]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__0__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[31]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[31]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__0__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[30]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[30]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__1__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[29]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[29]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__1__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[28]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[28]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__2__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[27]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[27]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__2__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[26]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[26]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__3__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[25]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[25]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__3__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[24]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[24]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__4__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[23]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[23]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__4__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[22]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[22]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__5__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[21]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[21]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__5__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[20]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[20]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__6__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[19]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[19]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__6__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[18]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[18]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__7__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[17]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[17]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__7__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[16]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[16]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__8__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[15]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[15]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__8__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[14]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[14]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__9__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[13]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[13]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__9__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[12]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[12]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__10__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[11]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[11]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__10__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[10]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[10]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__11__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[9]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[9]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__11__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[8]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[8]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__12__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[7]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[7]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__12__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[6]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[6]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__13__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[5]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[5]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__13__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[4]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[4]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__14__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[3]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[3]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__14__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[2]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[2]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__15__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[1]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[1]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_3__15__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[0]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[0]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__0__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[63]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[63]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__0__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[62]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[62]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__1__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[61]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[61]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__1__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[60]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[60]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__2__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[59]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[59]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__2__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[58]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[58]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__3__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[57]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[57]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__3__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[56]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[56]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__4__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[55]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[55]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__4__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[54]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[54]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__5__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[53]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[53]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__5__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[52]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[52]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__6__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[51]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[51]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__6__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[50]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[50]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__7__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[49]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[49]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__7__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[48]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[48]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__8__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[47]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[47]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__8__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[46]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[46]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__9__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[45]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[45]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__9__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[44]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[44]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__10__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[43]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[43]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__10__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[42]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[42]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__11__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[41]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[41]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__11__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[40]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[40]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__12__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[39]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[39]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__12__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[38]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[38]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__13__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[37]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[37]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__13__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[36]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[36]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__14__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[35]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[35]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__14__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[34]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[34]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__15__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[33]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[33]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_1__15__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[32]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[32]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__0__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[31]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[31]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__0__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[30]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[30]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__1__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[29]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[29]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__1__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[28]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[28]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__2__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[27]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[27]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__2__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[26]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[26]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__3__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[25]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[25]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__3__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[24]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[24]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__4__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[23]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[23]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__4__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[22]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[22]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__5__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[21]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[21]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__5__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[20]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[20]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__6__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[19]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[19]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__6__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[18]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[18]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__7__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[17]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[17]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__7__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[16]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[16]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__8__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[15]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[15]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__8__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[14]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[14]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__9__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[13]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[13]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__9__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[12]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[12]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__10__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[11]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[11]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__10__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[10]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[10]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__11__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[9]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[9]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__11__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[8]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[8]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__12__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[7]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[7]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__12__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[6]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[6]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__13__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[5]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[5]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__13__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[4]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[4]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__14__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[3]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[3]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__14__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[2]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[2]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__15__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[1]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[1]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_2__15__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[0]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[0]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__0__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[31]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[31]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__0__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[30]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[30]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__1__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[29]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[29]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__1__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[28]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[28]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__2__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[27]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[27]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__2__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[26]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[26]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__3__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[25]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[25]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__3__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[24]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[24]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__4__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[23]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[23]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__4__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[22]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[22]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__5__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[21]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[21]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__5__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[20]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[20]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__6__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[19]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[19]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__6__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[18]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[18]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__7__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[17]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[17]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__7__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[16]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[16]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__8__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[15]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[15]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__8__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[14]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[14]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__9__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[13]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[13]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__9__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[12]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[12]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__10__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[11]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[11]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__10__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[10]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[10]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__11__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[9]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[9]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__11__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[8]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[8]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__12__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[7]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[7]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__12__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[6]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[6]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__13__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[5]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[5]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__13__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[4]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[4]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__14__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[3]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[3]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__14__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[2]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[2]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__15__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[1]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[1]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_1__15__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[0]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[0]) );
  DFQD4BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__10__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[171]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[171]) );
  DFQD4BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__11__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[169]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[169]) );
  DFQD4BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__12__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[167]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[167]) );
  DFQD4BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__13__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[165]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[165]) );
  DFQD4BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__14__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[163]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[163]) );
  DFQD4BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__15__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[161]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[161]) );
  DFQD4BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__0__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[159]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[159]) );
  DFQD4BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__1__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[157]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[157]) );
  DFQD4BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__2__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[155]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[155]) );
  DFQD4BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__3__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[153]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[153]) );
  DFQD4BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__4__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[151]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[151]) );
  DFQD4BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__5__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[149]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[149]) );
  DFQD4BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__15__1_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[1]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[1]) );
  DFQD4BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__14__1_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[3]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[3]) );
  DFQD4BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__13__1_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[5]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[5]) );
  DFQD4BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__12__1_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[7]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[7]) );
  DFQD4BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__11__1_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[9]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[9]) );
  DFQD4BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__10__1_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[11]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[11]) );
  DFQD4BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__9__1_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[13]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[13]) );
  DFQD4BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__8__1_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[15]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[15]) );
  DFQD4BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__7__1_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[17]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[17]) );
  DFQD4BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__6__1_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[19]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[19]) );
  DFQD4BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__5__1_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[21]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[21]) );
  DFQD4BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__4__1_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[23]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[23]) );
  DFQD4BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__2__1_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[27]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[27]) );
  DFQD4BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__3__1_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[25]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[25]) );
  DFQD4BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__1__1_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[29]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[29]) );
  DFQD4BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__0__1_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[31]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[31]) );
  DFQD4BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__6__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[147]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[147]) );
  DFQD4BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__7__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[145]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[145]) );
  DFQD4BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__8__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[143]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[143]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__15__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[32]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[32]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__14__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[34]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[34]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__13__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[36]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[36]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__12__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[38]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[38]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__11__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[40]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[40]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__10__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[42]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[42]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__9__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[44]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[44]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__8__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[46]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[46]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__7__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[48]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[48]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__6__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[50]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[50]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__5__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[52]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[52]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__4__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[54]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[54]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__3__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[56]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[56]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__2__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[58]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[58]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__1__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[60]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[60]) );
  DFQD1BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__0__0_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[62]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[62]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__15__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[64]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[64]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__14__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[66]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[66]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__13__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[68]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[68]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__12__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[70]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[70]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__11__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[72]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[72]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__10__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[74]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[74]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__9__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[76]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[76]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__8__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[78]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[78]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__7__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[80]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[80]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__6__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[82]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[82]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__5__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[84]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[84]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__4__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[86]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[86]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__3__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[88]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[88]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__2__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[90]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[90]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__1__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[92]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[92]) );
  DFQD1BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__0__0_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[94]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[94]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__15__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[96]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[96]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__14__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[98]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[98]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__13__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[100]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[100]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__12__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[102]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[102]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__11__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[104]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[104]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__10__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[106]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[106]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__9__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[108]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[108]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__8__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[110]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[110]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__7__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[112]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[112]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__6__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[114]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[114]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__5__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[116]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[116]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__4__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[118]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[118]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__3__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[120]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[120]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__2__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[122]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[122]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__1__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[124]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[124]) );
  DFQD1BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__0__0_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[126]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[126]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__15__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[128]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[128]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__14__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[130]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[130]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__13__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[132]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[132]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__12__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[134]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[134]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__11__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[136]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[136]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__10__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[138]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[138]) );
  DFQD1BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__9__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[140]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[140]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__6__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[178]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[178]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__5__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[180]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[180]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__4__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[182]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[182]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__3__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[184]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[184]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__2__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[186]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[186]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__1__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[188]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[188]) );
  DFQD1BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__0__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[190]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[190]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__15__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[192]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[192]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__14__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[194]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[194]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__13__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[196]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[196]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__12__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[198]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[198]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__11__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[200]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[200]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__10__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[202]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[202]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__9__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[204]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[204]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__8__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[206]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[206]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__7__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[208]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[208]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__6__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[210]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[210]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__5__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[212]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[212]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__4__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[214]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[214]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__3__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[216]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[216]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__2__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[218]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[218]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__1__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[220]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[220]) );
  DFQD1BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__0__0_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[222]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[222]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__15__0_ ( .D(
        i_cmd[62]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[224]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__14__0_ ( .D(
        i_cmd[60]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[226]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__13__0_ ( .D(
        i_cmd[58]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[228]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__12__0_ ( .D(
        i_cmd[56]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[230]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__11__0_ ( .D(
        i_cmd[54]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[232]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__10__0_ ( .D(
        i_cmd[52]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[234]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__9__0_ ( .D(
        i_cmd[50]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[236]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__8__0_ ( .D(
        i_cmd[48]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[238]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__7__0_ ( .D(
        i_cmd[46]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[240]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__6__0_ ( .D(
        i_cmd[44]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[242]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__5__0_ ( .D(
        i_cmd[42]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[244]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__4__0_ ( .D(
        i_cmd[40]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[246]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__3__0_ ( .D(
        i_cmd[38]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[248]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__2__0_ ( .D(
        i_cmd[36]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[250]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__1__0_ ( .D(
        i_cmd[34]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[252]) );
  DFQD1BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__0__0_ ( .D(
        i_cmd[32]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[254]) );
  DFQD2BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__1__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[189]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[189]) );
  DFQD2BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__3__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[185]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[185]) );
  DFQD2BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__5__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[181]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[181]) );
  DFQD2BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__12__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[166]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[166]) );
  DFQD2BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__14__0_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[162]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[162]) );
  DFQD2BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__0__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[158]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[158]) );
  DFQD2BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__2__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[154]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[154]) );
  DFQD2BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__3__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[152]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[152]) );
  DFQD2BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__4__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[150]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[150]) );
  DFQD2BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__8__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[142]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[142]) );
  DFQD2BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__7__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[144]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[144]) );
  DFQD2BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__6__0_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[146]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[146]) );
  DFQD2BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__15__0_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[0]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[0]) );
  DFQD2BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__10__0_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[10]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[10]) );
  DFQD2BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__11__0_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[8]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[8]) );
  DFQD2BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__13__0_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[4]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[4]) );
  DFQD2BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__0__0_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[30]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[30]) );
  DFQD2BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__1__0_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[28]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[28]) );
  DFQD2BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__2__0_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[26]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[26]) );
  DFQD2BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__4__0_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[22]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[22]) );
  DFQD2BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__5__0_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[20]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[20]) );
  DFQD2BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__6__0_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[18]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[18]) );
  DFQD2BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__7__0_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[16]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[16]) );
  DFQD2BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__9__0_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[12]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[12]) );
  DFQD2BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__12__0_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[6]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[6]) );
  DFQD2BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__14__0_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[2]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[2]) );
  DFQD2BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__3__0_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[24]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[24]) );
  DFQD2BWP30P140 cmd_pipeline_stage_7__pipeline_i_cmd_reg_reg_0__8__0_ ( .D(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[14]), .CP(clk), .Q(
        cmd_pipeline_stage_7__pipeline_i_cmd_reg[14]) );
  DFQD2BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__7__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[177]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[177]) );
  DFQD2BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__8__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[175]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[175]) );
  DFQD2BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__9__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[173]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[173]) );
  DFQD2BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__0__1_ ( .D(
        i_cmd[33]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[255]) );
  DFQD2BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__2__1_ ( .D(
        i_cmd[37]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[251]) );
  DFQD2BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__3__1_ ( .D(
        i_cmd[39]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[249]) );
  DFQD2BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__4__1_ ( .D(
        i_cmd[41]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[247]) );
  DFQD2BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__6__1_ ( .D(
        i_cmd[45]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[243]) );
  DFQD2BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__7__1_ ( .D(
        i_cmd[47]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[241]) );
  DFQD2BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__8__1_ ( .D(
        i_cmd[49]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[239]) );
  DFQD2BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__10__1_ ( .D(
        i_cmd[53]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[235]) );
  DFQD2BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__12__1_ ( .D(
        i_cmd[57]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[231]) );
  DFQD2BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__14__1_ ( .D(
        i_cmd[61]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[227]) );
  DFQD2BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__0__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[223]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[223]) );
  DFQD2BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__2__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[219]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[219]) );
  DFQD2BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__4__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[215]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[215]) );
  DFQD2BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__6__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[211]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[211]) );
  DFQD2BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__8__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[207]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[207]) );
  DFQD2BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__9__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[205]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[205]) );
  DFQD2BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__10__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[203]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[203]) );
  DFQD2BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__11__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[201]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[201]) );
  DFQD2BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__12__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[199]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[199]) );
  DFQD2BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__14__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[195]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[195]) );
  DFQD2BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__15__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[193]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[193]) );
  DFQD2BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__0__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[191]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[191]) );
  DFQD2BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__2__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[187]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[187]) );
  DFQD2BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__4__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[183]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[183]) );
  DFQD2BWP30P140 cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__6__1_ ( .D(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[179]), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[179]) );
  DFQD2BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__1__1_ ( .D(
        i_cmd[35]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[253]) );
  DFQD2BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__5__1_ ( .D(
        i_cmd[43]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[245]) );
  DFQD2BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__9__1_ ( .D(
        i_cmd[51]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[237]) );
  DFQD2BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__11__1_ ( .D(
        i_cmd[55]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[233]) );
  DFQD2BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__13__1_ ( .D(
        i_cmd[59]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[229]) );
  DFQD2BWP30P140 cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__15__1_ ( .D(
        i_cmd[63]), .CP(clk), .Q(cmd_pipeline_stage_0__pipeline_i_cmd_reg[225]) );
  DFQD2BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__1__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[221]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[221]) );
  DFQD2BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__3__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[217]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[217]) );
  DFQD2BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__5__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[213]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[213]) );
  DFQD2BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__7__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[209]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[209]) );
  DFQD2BWP30P140 cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__13__1_ ( .D(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg[197]), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg[197]) );
  DFQD2BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__9__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[141]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[141]) );
  DFQD2BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__10__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[139]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[139]) );
  DFQD2BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__11__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[137]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[137]) );
  DFQD2BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__12__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[135]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[135]) );
  DFQD2BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__13__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[133]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[133]) );
  DFQD2BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__14__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[131]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[131]) );
  DFQD2BWP30P140 cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__15__1_ ( .D(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg[129]), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[129]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__0__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[127]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[127]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__1__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[125]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[125]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__2__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[123]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[123]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__3__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[121]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[121]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__4__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[119]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[119]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__5__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[117]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[117]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__6__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[115]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[115]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__7__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[113]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[113]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__8__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[111]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[111]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__9__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[109]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[109]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__10__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[107]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[107]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__11__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[105]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[105]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__12__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[103]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[103]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__13__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[101]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[101]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__14__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[99]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[99]) );
  DFQD2BWP30P140 cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__15__1_ ( .D(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[97]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[97]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__0__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[95]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[95]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__1__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[93]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[93]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__2__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[91]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[91]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__3__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[89]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[89]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__4__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[87]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[87]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__5__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[85]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[85]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__6__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[83]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[83]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__7__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[81]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[81]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__8__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[79]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[79]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__9__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[77]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[77]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__10__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[75]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[75]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__11__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[73]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[73]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__12__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[71]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[71]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__13__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[69]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[69]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__14__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[67]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[67]) );
  DFQD2BWP30P140 cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__15__1_ ( .D(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[65]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[65]) );
  DFQD2BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__0__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[63]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[63]) );
  DFQD2BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__1__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[61]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[61]) );
  DFQD2BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__2__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[59]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[59]) );
  DFQD2BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__3__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[57]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[57]) );
  DFQD2BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__4__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[55]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[55]) );
  DFQD2BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__5__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[53]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[53]) );
  DFQD2BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__6__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[51]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[51]) );
  DFQD2BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__7__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[49]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[49]) );
  DFQD2BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__8__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[47]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[47]) );
  DFQD2BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__9__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[45]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[45]) );
  DFQD2BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__10__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[43]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[43]) );
  DFQD2BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__11__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[41]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[41]) );
  DFQD2BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__12__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[39]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[39]) );
  DFQD2BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__13__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[37]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[37]) );
  DFQD2BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__14__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[35]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[35]) );
  DFQD2BWP30P140 cmd_pipeline_stage_6__pipeline_i_cmd_reg_reg_0__15__1_ ( .D(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[33]), .CP(clk), .Q(
        cmd_pipeline_stage_6__pipeline_i_cmd_reg[33]) );
  INVD6BWP30P140 U5 ( .I(n2315), .ZN(n174) );
  INVD6BWP30P140 U6 ( .I(n2063), .ZN(n292) );
  INVD6BWP30P140 U7 ( .I(n2034), .ZN(n321) );
  INVD6BWP30P140 U8 ( .I(n2313), .ZN(n177) );
  INVD6BWP30P140 U9 ( .I(n2371), .ZN(n12) );
  INVD6BWP30P140 U10 ( .I(n2314), .ZN(n176) );
  INVD6BWP30P140 U11 ( .I(n2064), .ZN(n291) );
  INVD6BWP30P140 U12 ( .I(n2059), .ZN(n296) );
  INVD6BWP30P140 U13 ( .I(n2319), .ZN(n170) );
  INVD6BWP30P140 U14 ( .I(n2368), .ZN(n9) );
  INVD6BWP30P140 U15 ( .I(n2058), .ZN(n297) );
  INVD6BWP30P140 U16 ( .I(n2320), .ZN(n169) );
  INVD6BWP30P140 U17 ( .I(n2356), .ZN(n137) );
  INVD6BWP30P140 U18 ( .I(n2036), .ZN(n319) );
  INVD6BWP30P140 U19 ( .I(n2062), .ZN(n293) );
  INVD6BWP30P140 U20 ( .I(n2316), .ZN(n173) );
  INVD6BWP30P140 U21 ( .I(n2370), .ZN(n11) );
  INVD6BWP30P140 U22 ( .I(n2355), .ZN(n138) );
  INVD6BWP30P140 U23 ( .I(n2035), .ZN(n320) );
  INVD6BWP30P140 U24 ( .I(n2061), .ZN(n294) );
  INVD6BWP30P140 U25 ( .I(n2317), .ZN(n172) );
  INVD6BWP30P140 U26 ( .I(n2369), .ZN(n10) );
  INVD6BWP30P140 U27 ( .I(n2060), .ZN(n295) );
  INVD6BWP30P140 U28 ( .I(n2318), .ZN(n171) );
  INVD6BWP30P140 U29 ( .I(n2000), .ZN(n323) );
  INVD6BWP30P140 U30 ( .I(n2376), .ZN(n17) );
  INVD6BWP30P140 U31 ( .I(n2375), .ZN(n16) );
  INVD6BWP30P140 U32 ( .I(n1996), .ZN(n327) );
  INVD6BWP30P140 U33 ( .I(n2378), .ZN(n19) );
  INVD6BWP30P140 U34 ( .I(n2309), .ZN(n181) );
  INVD6BWP30P140 U35 ( .I(n1997), .ZN(n326) );
  INVD6BWP30P140 U36 ( .I(n1998), .ZN(n325) );
  INVD6BWP30P140 U37 ( .I(n2377), .ZN(n18) );
  INVD6BWP30P140 U38 ( .I(n1999), .ZN(n324) );
  INVD6BWP30P140 U39 ( .I(n2310), .ZN(n180) );
  INVD6BWP30P140 U40 ( .I(n2373), .ZN(n14) );
  INVD6BWP30P140 U41 ( .I(n2311), .ZN(n179) );
  INVD6BWP30P140 U42 ( .I(n2354), .ZN(n139) );
  INVD6BWP30P140 U43 ( .I(n2372), .ZN(n13) );
  INVD6BWP30P140 U44 ( .I(n2312), .ZN(n178) );
  INVD6BWP30P140 U45 ( .I(n2353), .ZN(n140) );
  INVD6BWP30P140 U46 ( .I(n2308), .ZN(n182) );
  INVD6BWP30P140 U47 ( .I(n2374), .ZN(n15) );
  INVD6BWP30P140 U48 ( .I(n2033), .ZN(n322) );
  INVD6BWP30P140 U49 ( .I(n2366), .ZN(n7) );
  INVD6BWP30P140 U50 ( .I(n2040), .ZN(n315) );
  INVD6BWP30P140 U51 ( .I(n2365), .ZN(n6) );
  INVD6BWP30P140 U52 ( .I(n2041), .ZN(n314) );
  INVD6BWP30P140 U53 ( .I(n2360), .ZN(n133) );
  INVD6BWP30P140 U54 ( .I(n2359), .ZN(n134) );
  INVD6BWP30P140 U55 ( .I(n2363), .ZN(n4) );
  INVD6BWP30P140 U56 ( .I(n2046), .ZN(n309) );
  INVD6BWP30P140 U57 ( .I(n2043), .ZN(n312) );
  INVD6BWP30P140 U58 ( .I(n2361), .ZN(n132) );
  INVD6BWP30P140 U59 ( .I(n2045), .ZN(n310) );
  INVD6BWP30P140 U60 ( .I(n2362), .ZN(n131) );
  INVD6BWP30P140 U61 ( .I(n2044), .ZN(n311) );
  INVD6BWP30P140 U62 ( .I(n2049), .ZN(n306) );
  INVD6BWP30P140 U63 ( .I(n2048), .ZN(n307) );
  INVD6BWP30P140 U64 ( .I(n2364), .ZN(n5) );
  INVD6BWP30P140 U65 ( .I(n2042), .ZN(n313) );
  INVD6BWP30P140 U66 ( .I(n2047), .ZN(n308) );
  INVD6BWP30P140 U67 ( .I(n2037), .ZN(n318) );
  INVD6BWP30P140 U68 ( .I(n2054), .ZN(n301) );
  INVD6BWP30P140 U69 ( .I(n2357), .ZN(n136) );
  INVD6BWP30P140 U70 ( .I(n2057), .ZN(n298) );
  INVD6BWP30P140 U71 ( .I(n2056), .ZN(n299) );
  INVD6BWP30P140 U72 ( .I(n2055), .ZN(n300) );
  INVD6BWP30P140 U73 ( .I(n2050), .ZN(n305) );
  INVD6BWP30P140 U74 ( .I(n2039), .ZN(n316) );
  INVD6BWP30P140 U75 ( .I(n2367), .ZN(n8) );
  INVD6BWP30P140 U76 ( .I(n2053), .ZN(n302) );
  INVD6BWP30P140 U77 ( .I(n2038), .ZN(n317) );
  INVD6BWP30P140 U78 ( .I(n2052), .ZN(n303) );
  INVD6BWP30P140 U79 ( .I(n2358), .ZN(n135) );
  INVD6BWP30P140 U80 ( .I(n2051), .ZN(n304) );
  INVD6BWP30P140 U81 ( .I(n2232), .ZN(n130) );
  INVD6BWP30P140 U82 ( .I(n2634), .ZN(n197) );
  INVD6BWP30P140 U83 ( .I(n2231), .ZN(n129) );
  INVD6BWP30P140 U84 ( .I(n2230), .ZN(n128) );
  INVD6BWP30P140 U85 ( .I(n2161), .ZN(n175) );
  INVD6BWP30P140 U86 ( .I(n2229), .ZN(n127) );
  INVD6BWP30P140 U87 ( .I(n2635), .ZN(n196) );
  INVD6BWP30P140 U88 ( .I(n2632), .ZN(n199) );
  INVD6BWP30P140 U89 ( .I(n2233), .ZN(n190) );
  INVD6BWP30P140 U90 ( .I(n2633), .ZN(n198) );
  INVD6BWP30P140 U91 ( .I(n2166), .ZN(n71) );
  INVD6BWP30P140 U92 ( .I(n2228), .ZN(n126) );
  INVD6BWP30P140 U93 ( .I(n2162), .ZN(n67) );
  INVD6BWP30P140 U94 ( .I(n2227), .ZN(n125) );
  INVD6BWP30P140 U95 ( .I(n2163), .ZN(n68) );
  INVD6BWP30P140 U96 ( .I(n2226), .ZN(n124) );
  INVD6BWP30P140 U97 ( .I(n2164), .ZN(n69) );
  INVD6BWP30P140 U98 ( .I(n2225), .ZN(n100) );
  INVD6BWP30P140 U99 ( .I(n2165), .ZN(n70) );
  INVD6BWP30P140 U100 ( .I(n2243), .ZN(n114) );
  INVD6BWP30P140 U101 ( .I(n2242), .ZN(n115) );
  INVD6BWP30P140 U102 ( .I(n2241), .ZN(n116) );
  INVD6BWP30P140 U103 ( .I(n2240), .ZN(n117) );
  INVD6BWP30P140 U104 ( .I(n2626), .ZN(n205) );
  INVD6BWP30P140 U105 ( .I(n2247), .ZN(n110) );
  INVD6BWP30P140 U106 ( .I(n2246), .ZN(n111) );
  INVD6BWP30P140 U107 ( .I(n2245), .ZN(n112) );
  INVD6BWP30P140 U108 ( .I(n2244), .ZN(n113) );
  INVD6BWP30P140 U109 ( .I(n2627), .ZN(n204) );
  INVD6BWP30P140 U110 ( .I(n2630), .ZN(n201) );
  INVD6BWP30P140 U111 ( .I(n2631), .ZN(n200) );
  INVD6BWP30P140 U112 ( .I(n2239), .ZN(n118) );
  INVD6BWP30P140 U113 ( .I(n2628), .ZN(n203) );
  INVD6BWP30P140 U114 ( .I(n2238), .ZN(n119) );
  INVD6BWP30P140 U115 ( .I(n2237), .ZN(n120) );
  INVD6BWP30P140 U116 ( .I(n2236), .ZN(n121) );
  INVD6BWP30P140 U117 ( .I(n2629), .ZN(n202) );
  INVD6BWP30P140 U118 ( .I(n2235), .ZN(n122) );
  INVD6BWP30P140 U119 ( .I(n2234), .ZN(n123) );
  INVD6BWP30P140 U120 ( .I(n2637), .ZN(n194) );
  INVD6BWP30P140 U121 ( .I(n2175), .ZN(n80) );
  INVD6BWP30P140 U122 ( .I(n2638), .ZN(n193) );
  INVD6BWP30P140 U123 ( .I(n2192), .ZN(n97) );
  INVD6BWP30P140 U124 ( .I(n2176), .ZN(n81) );
  INVD6BWP30P140 U125 ( .I(n2636), .ZN(n195) );
  INVD6BWP30P140 U126 ( .I(n2182), .ZN(n87) );
  INVD6BWP30P140 U127 ( .I(n2191), .ZN(n96) );
  INVD6BWP30P140 U128 ( .I(n2183), .ZN(n88) );
  INVD6BWP30P140 U129 ( .I(n2184), .ZN(n89) );
  INVD6BWP30P140 U130 ( .I(n2190), .ZN(n95) );
  INVD6BWP30P140 U131 ( .I(n2185), .ZN(n90) );
  INVD6BWP30P140 U132 ( .I(n2189), .ZN(n94) );
  INVD6BWP30P140 U133 ( .I(n2186), .ZN(n91) );
  INVD6BWP30P140 U134 ( .I(n2188), .ZN(n93) );
  INVD6BWP30P140 U135 ( .I(n2187), .ZN(n92) );
  INVD6BWP30P140 U136 ( .I(n2177), .ZN(n82) );
  INVD6BWP30P140 U137 ( .I(n2639), .ZN(n192) );
  INVD6BWP30P140 U138 ( .I(n2178), .ZN(n83) );
  INVD6BWP30P140 U139 ( .I(n2179), .ZN(n84) );
  INVD6BWP30P140 U140 ( .I(n2640), .ZN(n191) );
  INVD6BWP30P140 U141 ( .I(n2180), .ZN(n85) );
  INVD6BWP30P140 U142 ( .I(n2181), .ZN(n86) );
  INVD6BWP30P140 U143 ( .I(n2167), .ZN(n72) );
  INVD6BWP30P140 U144 ( .I(n2168), .ZN(n73) );
  INVD6BWP30P140 U145 ( .I(n2173), .ZN(n78) );
  INVD6BWP30P140 U146 ( .I(n2174), .ZN(n79) );
  INVD6BWP30P140 U147 ( .I(n2169), .ZN(n74) );
  INVD6BWP30P140 U148 ( .I(n2170), .ZN(n75) );
  INVD6BWP30P140 U149 ( .I(n2171), .ZN(n76) );
  INVD6BWP30P140 U150 ( .I(n2172), .ZN(n77) );
  INVD6BWP30P140 U151 ( .I(n2617), .ZN(n214) );
  INVD6BWP30P140 U152 ( .I(n2097), .ZN(n290) );
  INVD6BWP30P140 U153 ( .I(n2292), .ZN(n64) );
  INVD6BWP30P140 U154 ( .I(n2098), .ZN(n289) );
  INVD6BWP30P140 U155 ( .I(n2291), .ZN(n65) );
  INVD6BWP30P140 U156 ( .I(n2099), .ZN(n288) );
  INVD6BWP30P140 U157 ( .I(n2290), .ZN(n66) );
  INVD6BWP30P140 U158 ( .I(n2100), .ZN(n287) );
  INVD6BWP30P140 U159 ( .I(n2289), .ZN(n98) );
  INVD6BWP30P140 U160 ( .I(n2615), .ZN(n216) );
  INVD6BWP30P140 U161 ( .I(n2616), .ZN(n215) );
  INVD6BWP30P140 U162 ( .I(n2106), .ZN(n146) );
  INVD6BWP30P140 U163 ( .I(n2619), .ZN(n212) );
  INVD6BWP30P140 U164 ( .I(n2107), .ZN(n147) );
  INVD6BWP30P140 U165 ( .I(n2105), .ZN(n145) );
  INVD6BWP30P140 U166 ( .I(n2618), .ZN(n213) );
  INVD6BWP30P140 U167 ( .I(n2101), .ZN(n141) );
  INVD6BWP30P140 U168 ( .I(n2102), .ZN(n142) );
  INVD6BWP30P140 U169 ( .I(n2103), .ZN(n143) );
  INVD6BWP30P140 U170 ( .I(n2104), .ZN(n144) );
  INVD6BWP30P140 U171 ( .I(n2303), .ZN(n187) );
  INVD6BWP30P140 U172 ( .I(n2302), .ZN(n188) );
  INVD6BWP30P140 U173 ( .I(n2301), .ZN(n189) );
  INVD6BWP30P140 U174 ( .I(n2610), .ZN(n221) );
  INVD6BWP30P140 U175 ( .I(n2300), .ZN(n99) );
  INVD6BWP30P140 U176 ( .I(n2307), .ZN(n183) );
  INVD6BWP30P140 U177 ( .I(n2306), .ZN(n184) );
  INVD6BWP30P140 U178 ( .I(n2305), .ZN(n185) );
  INVD6BWP30P140 U179 ( .I(n2609), .ZN(n222) );
  INVD6BWP30P140 U180 ( .I(n2304), .ZN(n186) );
  INVD6BWP30P140 U181 ( .I(n2294), .ZN(n62) );
  INVD6BWP30P140 U182 ( .I(n2613), .ZN(n218) );
  INVD6BWP30P140 U183 ( .I(n2293), .ZN(n63) );
  INVD6BWP30P140 U184 ( .I(n2614), .ZN(n217) );
  INVD6BWP30P140 U185 ( .I(n2299), .ZN(n57) );
  INVD6BWP30P140 U186 ( .I(n2298), .ZN(n58) );
  INVD6BWP30P140 U187 ( .I(n2297), .ZN(n59) );
  INVD6BWP30P140 U188 ( .I(n2611), .ZN(n220) );
  INVD6BWP30P140 U189 ( .I(n2296), .ZN(n60) );
  INVD6BWP30P140 U190 ( .I(n2612), .ZN(n219) );
  INVD6BWP30P140 U191 ( .I(n2295), .ZN(n61) );
  INVD6BWP30P140 U192 ( .I(n2255), .ZN(n102) );
  INVD6BWP30P140 U193 ( .I(n2124), .ZN(n164) );
  INVD6BWP30P140 U194 ( .I(n2621), .ZN(n210) );
  INVD6BWP30P140 U195 ( .I(n2254), .ZN(n103) );
  INVD6BWP30P140 U196 ( .I(n2253), .ZN(n104) );
  INVD6BWP30P140 U197 ( .I(n2252), .ZN(n105) );
  INVD6BWP30P140 U198 ( .I(n2622), .ZN(n209) );
  INVD6BWP30P140 U199 ( .I(n2251), .ZN(n106) );
  INVD6BWP30P140 U200 ( .I(n2120), .ZN(n160) );
  INVD6BWP30P140 U201 ( .I(n2121), .ZN(n161) );
  INVD6BWP30P140 U202 ( .I(n2122), .ZN(n162) );
  INVD6BWP30P140 U203 ( .I(n2123), .ZN(n163) );
  INVD6BWP30P140 U204 ( .I(n2620), .ZN(n211) );
  INVD6BWP30P140 U205 ( .I(n2256), .ZN(n101) );
  INVD6BWP30P140 U206 ( .I(n2127), .ZN(n167) );
  INVD6BWP30P140 U207 ( .I(n2128), .ZN(n168) );
  INVD6BWP30P140 U208 ( .I(n2625), .ZN(n206) );
  INVD6BWP30P140 U209 ( .I(n2250), .ZN(n107) );
  INVD6BWP30P140 U210 ( .I(n2249), .ZN(n108) );
  INVD6BWP30P140 U211 ( .I(n2248), .ZN(n109) );
  INVD6BWP30P140 U212 ( .I(n2623), .ZN(n208) );
  INVD6BWP30P140 U213 ( .I(n2125), .ZN(n165) );
  INVD6BWP30P140 U214 ( .I(n2624), .ZN(n207) );
  INVD6BWP30P140 U215 ( .I(n2126), .ZN(n166) );
  INVD6BWP30P140 U216 ( .I(n2108), .ZN(n148) );
  INVD6BWP30P140 U217 ( .I(n2109), .ZN(n149) );
  INVD6BWP30P140 U218 ( .I(n2115), .ZN(n155) );
  INVD6BWP30P140 U219 ( .I(n2116), .ZN(n156) );
  INVD6BWP30P140 U220 ( .I(n2117), .ZN(n157) );
  INVD6BWP30P140 U221 ( .I(n2118), .ZN(n158) );
  INVD6BWP30P140 U222 ( .I(n2119), .ZN(n159) );
  INVD6BWP30P140 U223 ( .I(n2110), .ZN(n150) );
  INVD6BWP30P140 U224 ( .I(n2111), .ZN(n151) );
  INVD6BWP30P140 U225 ( .I(n2112), .ZN(n152) );
  INVD6BWP30P140 U226 ( .I(n2113), .ZN(n153) );
  INVD6BWP30P140 U227 ( .I(n2114), .ZN(n154) );
  INVD6BWP30P140 U228 ( .I(n2424), .ZN(n50) );
  INVD6BWP30P140 U229 ( .I(n2569), .ZN(n262) );
  INVD6BWP30P140 U230 ( .I(n1799), .ZN(n428) );
  INVD6BWP30P140 U231 ( .I(n2546), .ZN(n285) );
  INVD6BWP30P140 U232 ( .I(n2425), .ZN(n49) );
  INVD6BWP30P140 U233 ( .I(n1724), .ZN(n471) );
  INVD6BWP30P140 U234 ( .I(n1800), .ZN(n427) );
  INVD6BWP30P140 U235 ( .I(n2568), .ZN(n263) );
  INVD6BWP30P140 U236 ( .I(n2426), .ZN(n48) );
  INVD6BWP30P140 U237 ( .I(n2421), .ZN(n53) );
  INVD6BWP30P140 U238 ( .I(n2484), .ZN(n251) );
  INVD6BWP30P140 U239 ( .I(n1797), .ZN(n430) );
  INVD6BWP30P140 U240 ( .I(n2422), .ZN(n52) );
  INVD6BWP30P140 U241 ( .I(n1726), .ZN(n469) );
  INVD6BWP30P140 U242 ( .I(n2559), .ZN(n272) );
  INVD6BWP30P140 U243 ( .I(n2570), .ZN(n261) );
  INVD6BWP30P140 U244 ( .I(n2423), .ZN(n51) );
  INVD6BWP30P140 U245 ( .I(n1725), .ZN(n470) );
  INVD6BWP30P140 U246 ( .I(n1798), .ZN(n429) );
  INVD6BWP30P140 U247 ( .I(n1802), .ZN(n425) );
  INVD6BWP30P140 U248 ( .I(n2545), .ZN(n284) );
  INVD6BWP30P140 U249 ( .I(n1803), .ZN(n424) );
  INVD6BWP30P140 U250 ( .I(n1721), .ZN(n474) );
  INVD6BWP30P140 U251 ( .I(n2500), .ZN(n235) );
  INVD6BWP30P140 U252 ( .I(n1872), .ZN(n387) );
  INVD6BWP30P140 U253 ( .I(n2567), .ZN(n264) );
  INVD6BWP30P140 U254 ( .I(n1801), .ZN(n426) );
  INVD6BWP30P140 U255 ( .I(n1723), .ZN(n472) );
  INVD6BWP30P140 U256 ( .I(n2501), .ZN(n234) );
  INVD6BWP30P140 U257 ( .I(n2566), .ZN(n265) );
  INVD6BWP30P140 U258 ( .I(n1722), .ZN(n473) );
  INVD6BWP30P140 U259 ( .I(n1791), .ZN(n436) );
  INVD6BWP30P140 U260 ( .I(n1917), .ZN(n374) );
  INVD6BWP30P140 U261 ( .I(n1916), .ZN(n375) );
  INVD6BWP30P140 U262 ( .I(n2503), .ZN(n232) );
  INVD6BWP30P140 U263 ( .I(n1915), .ZN(n376) );
  INVD6BWP30P140 U264 ( .I(n1914), .ZN(n377) );
  INVD6BWP30P140 U265 ( .I(n1913), .ZN(n378) );
  INVD6BWP30P140 U266 ( .I(n2502), .ZN(n233) );
  INVD6BWP30P140 U267 ( .I(n2547), .ZN(n286) );
  INVD6BWP30P140 U268 ( .I(n1912), .ZN(n379) );
  INVD6BWP30P140 U269 ( .I(n2482), .ZN(n253) );
  INVD6BWP30P140 U270 ( .I(n2506), .ZN(n229) );
  INVD6BWP30P140 U271 ( .I(n1922), .ZN(n369) );
  INVD6BWP30P140 U272 ( .I(n1921), .ZN(n370) );
  INVD6BWP30P140 U273 ( .I(n1790), .ZN(n437) );
  INVD6BWP30P140 U274 ( .I(n1920), .ZN(n371) );
  INVD6BWP30P140 U275 ( .I(n2573), .ZN(n258) );
  INVD6BWP30P140 U276 ( .I(n2505), .ZN(n230) );
  INVD6BWP30P140 U277 ( .I(n1919), .ZN(n372) );
  INVD6BWP30P140 U278 ( .I(n1918), .ZN(n373) );
  INVD6BWP30P140 U279 ( .I(n2557), .ZN(n274) );
  INVD6BWP30P140 U280 ( .I(n2504), .ZN(n231) );
  INVD6BWP30P140 U281 ( .I(n2419), .ZN(n55) );
  INVD6BWP30P140 U282 ( .I(n1905), .ZN(n386) );
  INVD6BWP30P140 U283 ( .I(n1729), .ZN(n466) );
  INVD6BWP30P140 U284 ( .I(n1794), .ZN(n433) );
  INVD6BWP30P140 U285 ( .I(n1728), .ZN(n467) );
  INVD6BWP30P140 U286 ( .I(n2420), .ZN(n54) );
  INVD6BWP30P140 U287 ( .I(n1795), .ZN(n432) );
  INVD6BWP30P140 U288 ( .I(n2571), .ZN(n260) );
  INVD6BWP30P140 U289 ( .I(n1727), .ZN(n468) );
  INVD6BWP30P140 U290 ( .I(n1796), .ZN(n431) );
  INVD6BWP30P140 U291 ( .I(n1731), .ZN(n464) );
  INVD6BWP30P140 U292 ( .I(n1792), .ZN(n435) );
  INVD6BWP30P140 U293 ( .I(n1911), .ZN(n380) );
  INVD6BWP30P140 U294 ( .I(n2483), .ZN(n252) );
  INVD6BWP30P140 U295 ( .I(n1910), .ZN(n381) );
  INVD6BWP30P140 U296 ( .I(n2417), .ZN(n3) );
  INVD6BWP30P140 U297 ( .I(n1909), .ZN(n382) );
  INVD6BWP30P140 U298 ( .I(n1908), .ZN(n383) );
  INVD6BWP30P140 U299 ( .I(n1907), .ZN(n384) );
  INVD6BWP30P140 U300 ( .I(n2418), .ZN(n56) );
  INVD6BWP30P140 U301 ( .I(n2558), .ZN(n273) );
  INVD6BWP30P140 U302 ( .I(n1793), .ZN(n434) );
  INVD6BWP30P140 U303 ( .I(n2572), .ZN(n259) );
  INVD6BWP30P140 U304 ( .I(n1730), .ZN(n465) );
  INVD6BWP30P140 U305 ( .I(n1906), .ZN(n385) );
  INVD6BWP30P140 U306 ( .I(n2490), .ZN(n245) );
  INVD6BWP30P140 U307 ( .I(n1843), .ZN(n416) );
  INVD6BWP30P140 U308 ( .I(n2438), .ZN(n36) );
  INVD6BWP30P140 U309 ( .I(n1842), .ZN(n417) );
  INVD6BWP30P140 U310 ( .I(n1717), .ZN(n478) );
  INVD6BWP30P140 U311 ( .I(n1841), .ZN(n418) );
  INVD6BWP30P140 U312 ( .I(n2489), .ZN(n246) );
  INVD6BWP30P140 U313 ( .I(n2439), .ZN(n35) );
  INVD6BWP30P140 U314 ( .I(n1716), .ZN(n479) );
  INVD6BWP30P140 U315 ( .I(n1848), .ZN(n411) );
  INVD6BWP30P140 U316 ( .I(n2561), .ZN(n270) );
  INVD6BWP30P140 U317 ( .I(n2436), .ZN(n38) );
  INVD6BWP30P140 U318 ( .I(n1847), .ZN(n412) );
  INVD6BWP30P140 U319 ( .I(n2491), .ZN(n244) );
  INVD6BWP30P140 U320 ( .I(n1846), .ZN(n413) );
  INVD6BWP30P140 U321 ( .I(n2437), .ZN(n37) );
  INVD6BWP30P140 U322 ( .I(n1845), .ZN(n414) );
  INVD6BWP30P140 U323 ( .I(n1844), .ZN(n415) );
  INVD6BWP30P140 U324 ( .I(n2442), .ZN(n32) );
  INVD6BWP30P140 U325 ( .I(n1714), .ZN(n481) );
  INVD6BWP30P140 U326 ( .I(n2486), .ZN(n249) );
  INVD6BWP30P140 U327 ( .I(n2485), .ZN(n250) );
  INVD6BWP30P140 U328 ( .I(n2443), .ZN(n31) );
  INVD6BWP30P140 U329 ( .I(n1713), .ZN(n482) );
  INVD6BWP30P140 U330 ( .I(n2440), .ZN(n34) );
  INVD6BWP30P140 U331 ( .I(n2488), .ZN(n247) );
  INVD6BWP30P140 U332 ( .I(n2441), .ZN(n33) );
  INVD6BWP30P140 U333 ( .I(n1715), .ZN(n480) );
  INVD6BWP30P140 U334 ( .I(n2487), .ZN(n248) );
  INVD6BWP30P140 U335 ( .I(n1865), .ZN(n394) );
  INVD6BWP30P140 U336 ( .I(n2427), .ZN(n47) );
  INVD6BWP30P140 U337 ( .I(n2446), .ZN(n28) );
  INVD6BWP30P140 U338 ( .I(n1864), .ZN(n395) );
  INVD6BWP30P140 U339 ( .I(n1807), .ZN(n420) );
  INVD6BWP30P140 U340 ( .I(n1719), .ZN(n476) );
  INVD6BWP30P140 U341 ( .I(n2496), .ZN(n239) );
  INVD6BWP30P140 U342 ( .I(n1863), .ZN(n396) );
  INVD6BWP30P140 U343 ( .I(n1862), .ZN(n397) );
  INVD6BWP30P140 U344 ( .I(n1861), .ZN(n398) );
  INVD6BWP30P140 U345 ( .I(n1808), .ZN(n419) );
  INVD6BWP30P140 U346 ( .I(n2445), .ZN(n29) );
  INVD6BWP30P140 U347 ( .I(n2428), .ZN(n46) );
  INVD6BWP30P140 U348 ( .I(n1860), .ZN(n399) );
  INVD6BWP30P140 U349 ( .I(n2495), .ZN(n240) );
  INVD6BWP30P140 U350 ( .I(n2564), .ZN(n267) );
  INVD6BWP30P140 U351 ( .I(n2565), .ZN(n266) );
  INVD6BWP30P140 U352 ( .I(n1871), .ZN(n388) );
  INVD6BWP30P140 U353 ( .I(n2560), .ZN(n271) );
  INVD6BWP30P140 U354 ( .I(n1804), .ZN(n423) );
  INVD6BWP30P140 U355 ( .I(n2448), .ZN(n26) );
  INVD6BWP30P140 U356 ( .I(n1720), .ZN(n475) );
  INVD6BWP30P140 U357 ( .I(n1870), .ZN(n389) );
  INVD6BWP30P140 U358 ( .I(n2499), .ZN(n236) );
  INVD6BWP30P140 U359 ( .I(n1869), .ZN(n390) );
  INVD6BWP30P140 U360 ( .I(n1868), .ZN(n391) );
  INVD6BWP30P140 U361 ( .I(n1805), .ZN(n422) );
  INVD6BWP30P140 U362 ( .I(n2498), .ZN(n237) );
  INVD6BWP30P140 U363 ( .I(n2447), .ZN(n27) );
  INVD6BWP30P140 U364 ( .I(n1867), .ZN(n392) );
  INVD6BWP30P140 U365 ( .I(n1866), .ZN(n393) );
  INVD6BWP30P140 U366 ( .I(n1806), .ZN(n421) );
  INVD6BWP30P140 U367 ( .I(n2497), .ZN(n238) );
  INVD6BWP30P140 U368 ( .I(n2432), .ZN(n42) );
  INVD6BWP30P140 U369 ( .I(n1853), .ZN(n406) );
  INVD6BWP30P140 U370 ( .I(n1852), .ZN(n407) );
  INVD6BWP30P140 U371 ( .I(n2433), .ZN(n41) );
  INVD6BWP30P140 U372 ( .I(n2562), .ZN(n269) );
  INVD6BWP30P140 U373 ( .I(n1851), .ZN(n408) );
  INVD6BWP30P140 U374 ( .I(n2434), .ZN(n40) );
  INVD6BWP30P140 U375 ( .I(n2492), .ZN(n243) );
  INVD6BWP30P140 U376 ( .I(n1850), .ZN(n409) );
  INVD6BWP30P140 U377 ( .I(n1849), .ZN(n410) );
  INVD6BWP30P140 U378 ( .I(n2435), .ZN(n39) );
  INVD6BWP30P140 U379 ( .I(n2429), .ZN(n45) );
  INVD6BWP30P140 U380 ( .I(n1859), .ZN(n400) );
  INVD6BWP30P140 U381 ( .I(n2494), .ZN(n241) );
  INVD6BWP30P140 U382 ( .I(n1858), .ZN(n401) );
  INVD6BWP30P140 U383 ( .I(n1857), .ZN(n402) );
  INVD6BWP30P140 U384 ( .I(n2430), .ZN(n44) );
  INVD6BWP30P140 U385 ( .I(n1856), .ZN(n403) );
  INVD6BWP30P140 U386 ( .I(n2563), .ZN(n268) );
  INVD6BWP30P140 U387 ( .I(n1718), .ZN(n477) );
  INVD6BWP30P140 U388 ( .I(n2444), .ZN(n30) );
  INVD6BWP30P140 U389 ( .I(n2431), .ZN(n43) );
  INVD6BWP30P140 U390 ( .I(n1855), .ZN(n404) );
  INVD6BWP30P140 U391 ( .I(n2493), .ZN(n242) );
  INVD6BWP30P140 U392 ( .I(n1854), .ZN(n405) );
  INVD6BWP30P140 U393 ( .I(n1976), .ZN(n347) );
  INVD6BWP30P140 U394 ( .I(n1975), .ZN(n348) );
  INVD6BWP30P140 U395 ( .I(n1974), .ZN(n349) );
  INVD6BWP30P140 U396 ( .I(n1973), .ZN(n350) );
  INVD6BWP30P140 U397 ( .I(n1742), .ZN(n453) );
  INVD6BWP30P140 U398 ( .I(n1979), .ZN(n344) );
  INVD6BWP30P140 U399 ( .I(n1978), .ZN(n345) );
  INVD6BWP30P140 U400 ( .I(n1743), .ZN(n452) );
  INVD6BWP30P140 U401 ( .I(n1977), .ZN(n346) );
  INVD6BWP30P140 U402 ( .I(n1740), .ZN(n455) );
  INVD6BWP30P140 U403 ( .I(n2548), .ZN(n283) );
  INVD6BWP30P140 U404 ( .I(n1972), .ZN(n351) );
  INVD6BWP30P140 U405 ( .I(n2553), .ZN(n278) );
  INVD6BWP30P140 U406 ( .I(n1971), .ZN(n352) );
  INVD6BWP30P140 U407 ( .I(n1970), .ZN(n353) );
  INVD6BWP30P140 U408 ( .I(n1969), .ZN(n354) );
  INVD6BWP30P140 U409 ( .I(n1741), .ZN(n454) );
  INVD6BWP30P140 U410 ( .I(n2381), .ZN(n22) );
  INVD6BWP30P140 U411 ( .I(n1990), .ZN(n333) );
  INVD6BWP30P140 U412 ( .I(n1989), .ZN(n334) );
  INVD6BWP30P140 U413 ( .I(n2551), .ZN(n280) );
  INVD6BWP30P140 U414 ( .I(n2382), .ZN(n23) );
  INVD6BWP30P140 U415 ( .I(n1988), .ZN(n335) );
  INVD6BWP30P140 U416 ( .I(n1987), .ZN(n336) );
  INVD6BWP30P140 U417 ( .I(n2383), .ZN(n24) );
  INVD6BWP30P140 U418 ( .I(n1995), .ZN(n328) );
  INVD6BWP30P140 U419 ( .I(n2550), .ZN(n281) );
  INVD6BWP30P140 U420 ( .I(n1994), .ZN(n329) );
  INVD6BWP30P140 U421 ( .I(n2379), .ZN(n20) );
  INVD6BWP30P140 U422 ( .I(n1993), .ZN(n330) );
  INVD6BWP30P140 U423 ( .I(n1992), .ZN(n331) );
  INVD6BWP30P140 U424 ( .I(n2380), .ZN(n21) );
  INVD6BWP30P140 U425 ( .I(n1991), .ZN(n332) );
  INVD6BWP30P140 U426 ( .I(n1982), .ZN(n341) );
  INVD6BWP30P140 U427 ( .I(n1981), .ZN(n342) );
  INVD6BWP30P140 U428 ( .I(n1744), .ZN(n451) );
  INVD6BWP30P140 U429 ( .I(n1980), .ZN(n343) );
  INVD6BWP30P140 U430 ( .I(n2552), .ZN(n279) );
  INVD6BWP30P140 U431 ( .I(n1986), .ZN(n337) );
  INVD6BWP30P140 U432 ( .I(n1985), .ZN(n338) );
  INVD6BWP30P140 U433 ( .I(n2384), .ZN(n25) );
  INVD6BWP30P140 U434 ( .I(n1984), .ZN(n339) );
  INVD6BWP30P140 U435 ( .I(n1983), .ZN(n340) );
  INVD6BWP30P140 U436 ( .I(n2549), .ZN(n282) );
  INVD6BWP30P140 U437 ( .I(n1735), .ZN(n460) );
  INVD6BWP30P140 U438 ( .I(n1782), .ZN(n445) );
  INVD6BWP30P140 U439 ( .I(n2510), .ZN(n225) );
  INVD6BWP30P140 U440 ( .I(n1936), .ZN(n355) );
  INVD6BWP30P140 U441 ( .I(n2481), .ZN(n254) );
  INVD6BWP30P140 U442 ( .I(n1783), .ZN(n444) );
  INVD6BWP30P140 U443 ( .I(n1935), .ZN(n356) );
  INVD6BWP30P140 U444 ( .I(n1934), .ZN(n357) );
  INVD6BWP30P140 U445 ( .I(n1784), .ZN(n443) );
  INVD6BWP30P140 U446 ( .I(n1933), .ZN(n358) );
  INVD6BWP30P140 U447 ( .I(n1736), .ZN(n459) );
  INVD6BWP30P140 U448 ( .I(n1780), .ZN(n447) );
  INVD6BWP30P140 U449 ( .I(n2511), .ZN(n224) );
  INVD6BWP30P140 U450 ( .I(n2555), .ZN(n276) );
  INVD6BWP30P140 U451 ( .I(n2576), .ZN(n255) );
  INVD6BWP30P140 U452 ( .I(n1781), .ZN(n446) );
  INVD6BWP30P140 U453 ( .I(n1932), .ZN(n359) );
  INVD6BWP30P140 U454 ( .I(n2508), .ZN(n227) );
  INVD6BWP30P140 U455 ( .I(n2574), .ZN(n257) );
  INVD6BWP30P140 U456 ( .I(n1787), .ZN(n440) );
  INVD6BWP30P140 U457 ( .I(n1733), .ZN(n462) );
  INVD6BWP30P140 U458 ( .I(n1927), .ZN(n364) );
  INVD6BWP30P140 U459 ( .I(n1788), .ZN(n439) );
  INVD6BWP30P140 U460 ( .I(n1926), .ZN(n365) );
  INVD6BWP30P140 U461 ( .I(n1928), .ZN(n363) );
  INVD6BWP30P140 U462 ( .I(n1925), .ZN(n366) );
  INVD6BWP30P140 U463 ( .I(n2507), .ZN(n228) );
  INVD6BWP30P140 U464 ( .I(n1789), .ZN(n438) );
  INVD6BWP30P140 U465 ( .I(n1924), .ZN(n367) );
  INVD6BWP30P140 U466 ( .I(n1732), .ZN(n463) );
  INVD6BWP30P140 U467 ( .I(n1923), .ZN(n368) );
  INVD6BWP30P140 U468 ( .I(n1734), .ZN(n461) );
  INVD6BWP30P140 U469 ( .I(n2509), .ZN(n226) );
  INVD6BWP30P140 U470 ( .I(n2575), .ZN(n256) );
  INVD6BWP30P140 U471 ( .I(n1785), .ZN(n442) );
  INVD6BWP30P140 U472 ( .I(n1931), .ZN(n360) );
  INVD6BWP30P140 U473 ( .I(n1786), .ZN(n441) );
  INVD6BWP30P140 U474 ( .I(n2556), .ZN(n275) );
  INVD6BWP30P140 U475 ( .I(n1930), .ZN(n361) );
  INVD6BWP30P140 U476 ( .I(n1929), .ZN(n362) );
  INVD6BWP30P140 U477 ( .I(n1738), .ZN(n457) );
  INVD6BWP30P140 U478 ( .I(n2512), .ZN(n223) );
  INVD6BWP30P140 U479 ( .I(n1778), .ZN(n449) );
  INVD6BWP30P140 U480 ( .I(n1777), .ZN(n450) );
  INVD6BWP30P140 U481 ( .I(n1737), .ZN(n458) );
  INVD6BWP30P140 U482 ( .I(n2554), .ZN(n277) );
  INVD6BWP30P140 U483 ( .I(n1779), .ZN(n448) );
  INVD6BWP30P140 U484 ( .I(n1739), .ZN(n456) );
  INVD2BWP30P140 U485 ( .I(n1680), .ZN(n483) );
  INVD2BWP30P140 U486 ( .I(n1679), .ZN(n484) );
  INVD2BWP30P140 U487 ( .I(n1678), .ZN(n485) );
  INVD2BWP30P140 U488 ( .I(n1677), .ZN(n486) );
  INVD2BWP30P140 U489 ( .I(n1676), .ZN(n487) );
  INVD2BWP30P140 U490 ( .I(n1675), .ZN(n488) );
  INVD2BWP30P140 U491 ( .I(n1674), .ZN(n489) );
  INVD2BWP30P140 U492 ( .I(n1673), .ZN(n490) );
  INVD2BWP30P140 U493 ( .I(n1672), .ZN(n491) );
  INVD2BWP30P140 U494 ( .I(n1671), .ZN(n492) );
  INVD2BWP30P140 U495 ( .I(n1670), .ZN(n493) );
  INVD2BWP30P140 U496 ( .I(n1669), .ZN(n494) );
  INVD2BWP30P140 U497 ( .I(n1668), .ZN(n495) );
  INVD2BWP30P140 U498 ( .I(n1667), .ZN(n496) );
  INVD2BWP30P140 U499 ( .I(n1666), .ZN(n497) );
  INVD2BWP30P140 U500 ( .I(n1665), .ZN(n498) );
  INVD2BWP30P140 U501 ( .I(n1664), .ZN(n499) );
  INVD2BWP30P140 U502 ( .I(n1663), .ZN(n500) );
  INVD2BWP30P140 U503 ( .I(n1662), .ZN(n501) );
  INVD2BWP30P140 U504 ( .I(n1661), .ZN(n502) );
  INVD2BWP30P140 U505 ( .I(n1660), .ZN(n503) );
  INVD2BWP30P140 U506 ( .I(n1659), .ZN(n504) );
  INVD2BWP30P140 U507 ( .I(n1658), .ZN(n505) );
  INVD2BWP30P140 U508 ( .I(n1657), .ZN(n506) );
  INVD2BWP30P140 U509 ( .I(n1656), .ZN(n507) );
  INVD2BWP30P140 U510 ( .I(n1655), .ZN(n508) );
  INVD2BWP30P140 U511 ( .I(n1654), .ZN(n509) );
  INVD2BWP30P140 U512 ( .I(n1653), .ZN(n510) );
  INVD2BWP30P140 U513 ( .I(n1652), .ZN(n511) );
  INVD2BWP30P140 U514 ( .I(n1651), .ZN(n512) );
  INVD15BWP30P140 U515 ( .I(n3), .ZN(o_data_bus[223]) );
  INVD15BWP30P140 U516 ( .I(n4), .ZN(o_data_bus[277]) );
  INVD15BWP30P140 U517 ( .I(n5), .ZN(o_data_bus[276]) );
  INVD15BWP30P140 U518 ( .I(n6), .ZN(o_data_bus[275]) );
  INVD15BWP30P140 U519 ( .I(n7), .ZN(o_data_bus[274]) );
  INVD15BWP30P140 U520 ( .I(n8), .ZN(o_data_bus[273]) );
  INVD15BWP30P140 U521 ( .I(n9), .ZN(o_data_bus[272]) );
  INVD15BWP30P140 U522 ( .I(n10), .ZN(o_data_bus[271]) );
  INVD15BWP30P140 U523 ( .I(n11), .ZN(o_data_bus[270]) );
  INVD15BWP30P140 U524 ( .I(n12), .ZN(o_data_bus[269]) );
  INVD15BWP30P140 U525 ( .I(n13), .ZN(o_data_bus[268]) );
  INVD15BWP30P140 U526 ( .I(n14), .ZN(o_data_bus[267]) );
  INVD15BWP30P140 U527 ( .I(n15), .ZN(o_data_bus[266]) );
  INVD15BWP30P140 U528 ( .I(n16), .ZN(o_data_bus[265]) );
  INVD15BWP30P140 U529 ( .I(n17), .ZN(o_data_bus[264]) );
  INVD15BWP30P140 U530 ( .I(n18), .ZN(o_data_bus[263]) );
  INVD15BWP30P140 U531 ( .I(n19), .ZN(o_data_bus[262]) );
  INVD15BWP30P140 U532 ( .I(n20), .ZN(o_data_bus[261]) );
  INVD15BWP30P140 U533 ( .I(n21), .ZN(o_data_bus[260]) );
  INVD15BWP30P140 U534 ( .I(n22), .ZN(o_data_bus[259]) );
  INVD15BWP30P140 U535 ( .I(n23), .ZN(o_data_bus[258]) );
  INVD15BWP30P140 U536 ( .I(n24), .ZN(o_data_bus[257]) );
  INVD15BWP30P140 U537 ( .I(n25), .ZN(o_data_bus[256]) );
  INVD15BWP30P140 U538 ( .I(n26), .ZN(o_data_bus[192]) );
  INVD15BWP30P140 U539 ( .I(n27), .ZN(o_data_bus[193]) );
  INVD15BWP30P140 U540 ( .I(n28), .ZN(o_data_bus[194]) );
  INVD15BWP30P140 U541 ( .I(n29), .ZN(o_data_bus[195]) );
  INVD15BWP30P140 U542 ( .I(n30), .ZN(o_data_bus[196]) );
  INVD15BWP30P140 U543 ( .I(n31), .ZN(o_data_bus[197]) );
  INVD15BWP30P140 U544 ( .I(n32), .ZN(o_data_bus[198]) );
  INVD15BWP30P140 U545 ( .I(n33), .ZN(o_data_bus[199]) );
  INVD15BWP30P140 U546 ( .I(n34), .ZN(o_data_bus[200]) );
  INVD15BWP30P140 U547 ( .I(n35), .ZN(o_data_bus[201]) );
  INVD15BWP30P140 U548 ( .I(n36), .ZN(o_data_bus[202]) );
  INVD15BWP30P140 U549 ( .I(n37), .ZN(o_data_bus[203]) );
  INVD15BWP30P140 U550 ( .I(n38), .ZN(o_data_bus[204]) );
  INVD15BWP30P140 U551 ( .I(n39), .ZN(o_data_bus[205]) );
  INVD15BWP30P140 U552 ( .I(n40), .ZN(o_data_bus[206]) );
  INVD15BWP30P140 U553 ( .I(n41), .ZN(o_data_bus[207]) );
  INVD15BWP30P140 U554 ( .I(n42), .ZN(o_data_bus[208]) );
  INVD15BWP30P140 U555 ( .I(n43), .ZN(o_data_bus[209]) );
  INVD15BWP30P140 U556 ( .I(n44), .ZN(o_data_bus[210]) );
  INVD15BWP30P140 U557 ( .I(n45), .ZN(o_data_bus[211]) );
  INVD15BWP30P140 U558 ( .I(n46), .ZN(o_data_bus[212]) );
  INVD15BWP30P140 U559 ( .I(n47), .ZN(o_data_bus[213]) );
  INVD15BWP30P140 U560 ( .I(n48), .ZN(o_data_bus[214]) );
  INVD15BWP30P140 U561 ( .I(n49), .ZN(o_data_bus[215]) );
  INVD15BWP30P140 U562 ( .I(n50), .ZN(o_data_bus[216]) );
  INVD15BWP30P140 U563 ( .I(n51), .ZN(o_data_bus[217]) );
  INVD15BWP30P140 U564 ( .I(n52), .ZN(o_data_bus[218]) );
  INVD15BWP30P140 U565 ( .I(n53), .ZN(o_data_bus[219]) );
  INVD15BWP30P140 U566 ( .I(n54), .ZN(o_data_bus[220]) );
  INVD15BWP30P140 U567 ( .I(n55), .ZN(o_data_bus[221]) );
  INVD15BWP30P140 U568 ( .I(n56), .ZN(o_data_bus[222]) );
  INVD15BWP30P140 U569 ( .I(n57), .ZN(o_data_bus[341]) );
  INVD15BWP30P140 U570 ( .I(n58), .ZN(o_data_bus[342]) );
  INVD15BWP30P140 U571 ( .I(n59), .ZN(o_data_bus[343]) );
  INVD15BWP30P140 U572 ( .I(n60), .ZN(o_data_bus[344]) );
  INVD15BWP30P140 U573 ( .I(n61), .ZN(o_data_bus[345]) );
  INVD15BWP30P140 U574 ( .I(n62), .ZN(o_data_bus[346]) );
  INVD15BWP30P140 U575 ( .I(n63), .ZN(o_data_bus[347]) );
  INVD15BWP30P140 U576 ( .I(n64), .ZN(o_data_bus[348]) );
  INVD15BWP30P140 U577 ( .I(n65), .ZN(o_data_bus[349]) );
  INVD15BWP30P140 U578 ( .I(n66), .ZN(o_data_bus[350]) );
  INVD15BWP30P140 U579 ( .I(n67), .ZN(o_data_bus[478]) );
  INVD15BWP30P140 U580 ( .I(n68), .ZN(o_data_bus[477]) );
  INVD15BWP30P140 U581 ( .I(n69), .ZN(o_data_bus[476]) );
  INVD15BWP30P140 U582 ( .I(n70), .ZN(o_data_bus[475]) );
  INVD15BWP30P140 U583 ( .I(n71), .ZN(o_data_bus[474]) );
  INVD15BWP30P140 U584 ( .I(n72), .ZN(o_data_bus[473]) );
  INVD15BWP30P140 U585 ( .I(n73), .ZN(o_data_bus[472]) );
  INVD15BWP30P140 U586 ( .I(n74), .ZN(o_data_bus[471]) );
  INVD15BWP30P140 U587 ( .I(n75), .ZN(o_data_bus[470]) );
  INVD15BWP30P140 U588 ( .I(n76), .ZN(o_data_bus[469]) );
  INVD15BWP30P140 U589 ( .I(n77), .ZN(o_data_bus[468]) );
  INVD15BWP30P140 U590 ( .I(n78), .ZN(o_data_bus[467]) );
  INVD15BWP30P140 U591 ( .I(n79), .ZN(o_data_bus[466]) );
  INVD15BWP30P140 U592 ( .I(n80), .ZN(o_data_bus[465]) );
  INVD15BWP30P140 U593 ( .I(n81), .ZN(o_data_bus[464]) );
  INVD15BWP30P140 U594 ( .I(n82), .ZN(o_data_bus[463]) );
  INVD15BWP30P140 U595 ( .I(n83), .ZN(o_data_bus[462]) );
  INVD15BWP30P140 U596 ( .I(n84), .ZN(o_data_bus[461]) );
  INVD15BWP30P140 U597 ( .I(n85), .ZN(o_data_bus[460]) );
  INVD15BWP30P140 U598 ( .I(n86), .ZN(o_data_bus[459]) );
  INVD15BWP30P140 U599 ( .I(n87), .ZN(o_data_bus[458]) );
  INVD15BWP30P140 U600 ( .I(n88), .ZN(o_data_bus[457]) );
  INVD15BWP30P140 U601 ( .I(n89), .ZN(o_data_bus[456]) );
  INVD15BWP30P140 U602 ( .I(n90), .ZN(o_data_bus[455]) );
  INVD15BWP30P140 U603 ( .I(n91), .ZN(o_data_bus[454]) );
  INVD15BWP30P140 U604 ( .I(n92), .ZN(o_data_bus[453]) );
  INVD15BWP30P140 U605 ( .I(n93), .ZN(o_data_bus[452]) );
  INVD15BWP30P140 U606 ( .I(n94), .ZN(o_data_bus[451]) );
  INVD15BWP30P140 U607 ( .I(n95), .ZN(o_data_bus[450]) );
  INVD15BWP30P140 U608 ( .I(n96), .ZN(o_data_bus[449]) );
  INVD15BWP30P140 U609 ( .I(n97), .ZN(o_data_bus[448]) );
  INVD15BWP30P140 U610 ( .I(n98), .ZN(o_data_bus[351]) );
  INVD15BWP30P140 U611 ( .I(n99), .ZN(o_data_bus[340]) );
  INVD15BWP30P140 U612 ( .I(n100), .ZN(o_data_bus[415]) );
  INVD15BWP30P140 U613 ( .I(n101), .ZN(o_data_bus[384]) );
  INVD15BWP30P140 U614 ( .I(n102), .ZN(o_data_bus[385]) );
  INVD15BWP30P140 U615 ( .I(n103), .ZN(o_data_bus[386]) );
  INVD15BWP30P140 U616 ( .I(n104), .ZN(o_data_bus[387]) );
  INVD15BWP30P140 U617 ( .I(n105), .ZN(o_data_bus[388]) );
  INVD15BWP30P140 U618 ( .I(n106), .ZN(o_data_bus[389]) );
  INVD15BWP30P140 U619 ( .I(n107), .ZN(o_data_bus[390]) );
  INVD15BWP30P140 U620 ( .I(n108), .ZN(o_data_bus[391]) );
  INVD15BWP30P140 U621 ( .I(n109), .ZN(o_data_bus[392]) );
  INVD15BWP30P140 U622 ( .I(n110), .ZN(o_data_bus[393]) );
  INVD15BWP30P140 U623 ( .I(n111), .ZN(o_data_bus[394]) );
  INVD15BWP30P140 U624 ( .I(n112), .ZN(o_data_bus[395]) );
  INVD15BWP30P140 U625 ( .I(n113), .ZN(o_data_bus[396]) );
  INVD15BWP30P140 U626 ( .I(n114), .ZN(o_data_bus[397]) );
  INVD15BWP30P140 U627 ( .I(n115), .ZN(o_data_bus[398]) );
  INVD15BWP30P140 U628 ( .I(n116), .ZN(o_data_bus[399]) );
  INVD15BWP30P140 U629 ( .I(n117), .ZN(o_data_bus[400]) );
  INVD15BWP30P140 U630 ( .I(n118), .ZN(o_data_bus[401]) );
  INVD15BWP30P140 U631 ( .I(n119), .ZN(o_data_bus[402]) );
  INVD15BWP30P140 U632 ( .I(n120), .ZN(o_data_bus[403]) );
  INVD15BWP30P140 U633 ( .I(n121), .ZN(o_data_bus[404]) );
  INVD15BWP30P140 U634 ( .I(n122), .ZN(o_data_bus[405]) );
  INVD15BWP30P140 U635 ( .I(n123), .ZN(o_data_bus[406]) );
  INVD15BWP30P140 U636 ( .I(n124), .ZN(o_data_bus[414]) );
  INVD15BWP30P140 U637 ( .I(n125), .ZN(o_data_bus[413]) );
  INVD15BWP30P140 U638 ( .I(n126), .ZN(o_data_bus[412]) );
  INVD15BWP30P140 U639 ( .I(n127), .ZN(o_data_bus[411]) );
  INVD15BWP30P140 U640 ( .I(n128), .ZN(o_data_bus[410]) );
  INVD15BWP30P140 U641 ( .I(n129), .ZN(o_data_bus[409]) );
  INVD15BWP30P140 U642 ( .I(n130), .ZN(o_data_bus[408]) );
  INVD15BWP30P140 U643 ( .I(n131), .ZN(o_data_bus[278]) );
  INVD15BWP30P140 U644 ( .I(n132), .ZN(o_data_bus[279]) );
  INVD15BWP30P140 U645 ( .I(n133), .ZN(o_data_bus[280]) );
  INVD15BWP30P140 U646 ( .I(n134), .ZN(o_data_bus[281]) );
  INVD15BWP30P140 U647 ( .I(n135), .ZN(o_data_bus[282]) );
  INVD15BWP30P140 U648 ( .I(n136), .ZN(o_data_bus[283]) );
  INVD15BWP30P140 U649 ( .I(n137), .ZN(o_data_bus[284]) );
  INVD15BWP30P140 U650 ( .I(n138), .ZN(o_data_bus[285]) );
  INVD15BWP30P140 U651 ( .I(n139), .ZN(o_data_bus[286]) );
  INVD15BWP30P140 U652 ( .I(n140), .ZN(o_data_bus[287]) );
  INVD15BWP30P140 U653 ( .I(n141), .ZN(o_data_bus[539]) );
  INVD15BWP30P140 U654 ( .I(n142), .ZN(o_data_bus[538]) );
  INVD15BWP30P140 U655 ( .I(n143), .ZN(o_data_bus[537]) );
  INVD15BWP30P140 U656 ( .I(n144), .ZN(o_data_bus[536]) );
  INVD15BWP30P140 U657 ( .I(n145), .ZN(o_data_bus[535]) );
  INVD15BWP30P140 U658 ( .I(n146), .ZN(o_data_bus[534]) );
  INVD15BWP30P140 U659 ( .I(n147), .ZN(o_data_bus[533]) );
  INVD15BWP30P140 U660 ( .I(n148), .ZN(o_data_bus[532]) );
  INVD15BWP30P140 U661 ( .I(n149), .ZN(o_data_bus[531]) );
  INVD15BWP30P140 U662 ( .I(n150), .ZN(o_data_bus[530]) );
  INVD15BWP30P140 U663 ( .I(n151), .ZN(o_data_bus[529]) );
  INVD15BWP30P140 U664 ( .I(n152), .ZN(o_data_bus[528]) );
  INVD15BWP30P140 U665 ( .I(n153), .ZN(o_data_bus[527]) );
  INVD15BWP30P140 U666 ( .I(n154), .ZN(o_data_bus[526]) );
  INVD15BWP30P140 U667 ( .I(n155), .ZN(o_data_bus[525]) );
  INVD15BWP30P140 U668 ( .I(n156), .ZN(o_data_bus[524]) );
  INVD15BWP30P140 U669 ( .I(n157), .ZN(o_data_bus[523]) );
  INVD15BWP30P140 U670 ( .I(n158), .ZN(o_data_bus[522]) );
  INVD15BWP30P140 U671 ( .I(n159), .ZN(o_data_bus[521]) );
  INVD15BWP30P140 U672 ( .I(n160), .ZN(o_data_bus[520]) );
  INVD15BWP30P140 U673 ( .I(n161), .ZN(o_data_bus[519]) );
  INVD15BWP30P140 U674 ( .I(n162), .ZN(o_data_bus[518]) );
  INVD15BWP30P140 U675 ( .I(n163), .ZN(o_data_bus[517]) );
  INVD15BWP30P140 U676 ( .I(n164), .ZN(o_data_bus[516]) );
  INVD15BWP30P140 U677 ( .I(n165), .ZN(o_data_bus[515]) );
  INVD15BWP30P140 U678 ( .I(n166), .ZN(o_data_bus[514]) );
  INVD15BWP30P140 U679 ( .I(n167), .ZN(o_data_bus[513]) );
  INVD15BWP30P140 U680 ( .I(n168), .ZN(o_data_bus[512]) );
  INVD15BWP30P140 U681 ( .I(n169), .ZN(o_data_bus[320]) );
  INVD15BWP30P140 U682 ( .I(n170), .ZN(o_data_bus[321]) );
  INVD15BWP30P140 U683 ( .I(n171), .ZN(o_data_bus[322]) );
  INVD15BWP30P140 U684 ( .I(n172), .ZN(o_data_bus[323]) );
  INVD15BWP30P140 U685 ( .I(n173), .ZN(o_data_bus[324]) );
  INVD15BWP30P140 U686 ( .I(n174), .ZN(o_data_bus[325]) );
  INVD15BWP30P140 U687 ( .I(n175), .ZN(o_data_bus[479]) );
  INVD15BWP30P140 U688 ( .I(n176), .ZN(o_data_bus[326]) );
  INVD15BWP30P140 U689 ( .I(n177), .ZN(o_data_bus[327]) );
  INVD15BWP30P140 U690 ( .I(n178), .ZN(o_data_bus[328]) );
  INVD15BWP30P140 U691 ( .I(n179), .ZN(o_data_bus[329]) );
  INVD15BWP30P140 U692 ( .I(n180), .ZN(o_data_bus[330]) );
  INVD15BWP30P140 U693 ( .I(n181), .ZN(o_data_bus[331]) );
  INVD15BWP30P140 U694 ( .I(n182), .ZN(o_data_bus[332]) );
  INVD15BWP30P140 U695 ( .I(n183), .ZN(o_data_bus[333]) );
  INVD15BWP30P140 U696 ( .I(n184), .ZN(o_data_bus[334]) );
  INVD15BWP30P140 U697 ( .I(n185), .ZN(o_data_bus[335]) );
  INVD15BWP30P140 U698 ( .I(n186), .ZN(o_data_bus[336]) );
  INVD15BWP30P140 U699 ( .I(n187), .ZN(o_data_bus[337]) );
  INVD15BWP30P140 U700 ( .I(n188), .ZN(o_data_bus[338]) );
  INVD15BWP30P140 U701 ( .I(n189), .ZN(o_data_bus[339]) );
  INVD15BWP30P140 U702 ( .I(n190), .ZN(o_data_bus[407]) );
  INVD15BWP30P140 U703 ( .I(n191), .ZN(o_data_bus[0]) );
  INVD15BWP30P140 U704 ( .I(n192), .ZN(o_data_bus[1]) );
  INVD15BWP30P140 U705 ( .I(n193), .ZN(o_data_bus[2]) );
  INVD15BWP30P140 U706 ( .I(n194), .ZN(o_data_bus[3]) );
  INVD15BWP30P140 U707 ( .I(n195), .ZN(o_data_bus[4]) );
  INVD15BWP30P140 U708 ( .I(n196), .ZN(o_data_bus[5]) );
  INVD15BWP30P140 U709 ( .I(n197), .ZN(o_data_bus[6]) );
  INVD15BWP30P140 U710 ( .I(n198), .ZN(o_data_bus[7]) );
  INVD15BWP30P140 U711 ( .I(n199), .ZN(o_data_bus[8]) );
  INVD15BWP30P140 U712 ( .I(n200), .ZN(o_data_bus[9]) );
  INVD15BWP30P140 U713 ( .I(n201), .ZN(o_data_bus[10]) );
  INVD15BWP30P140 U714 ( .I(n202), .ZN(o_data_bus[11]) );
  INVD15BWP30P140 U715 ( .I(n203), .ZN(o_data_bus[12]) );
  INVD15BWP30P140 U716 ( .I(n204), .ZN(o_data_bus[13]) );
  INVD15BWP30P140 U717 ( .I(n205), .ZN(o_data_bus[14]) );
  INVD15BWP30P140 U718 ( .I(n206), .ZN(o_data_bus[15]) );
  INVD15BWP30P140 U719 ( .I(n207), .ZN(o_data_bus[16]) );
  INVD15BWP30P140 U720 ( .I(n208), .ZN(o_data_bus[17]) );
  INVD15BWP30P140 U721 ( .I(n209), .ZN(o_data_bus[18]) );
  INVD15BWP30P140 U722 ( .I(n210), .ZN(o_data_bus[19]) );
  INVD15BWP30P140 U723 ( .I(n211), .ZN(o_data_bus[20]) );
  INVD15BWP30P140 U724 ( .I(n212), .ZN(o_data_bus[21]) );
  INVD15BWP30P140 U725 ( .I(n213), .ZN(o_data_bus[22]) );
  INVD15BWP30P140 U726 ( .I(n214), .ZN(o_data_bus[23]) );
  INVD15BWP30P140 U727 ( .I(n215), .ZN(o_data_bus[24]) );
  INVD15BWP30P140 U728 ( .I(n216), .ZN(o_data_bus[25]) );
  INVD15BWP30P140 U729 ( .I(n217), .ZN(o_data_bus[26]) );
  INVD15BWP30P140 U730 ( .I(n218), .ZN(o_data_bus[27]) );
  INVD15BWP30P140 U731 ( .I(n219), .ZN(o_data_bus[28]) );
  INVD15BWP30P140 U732 ( .I(n220), .ZN(o_data_bus[29]) );
  INVD15BWP30P140 U733 ( .I(n221), .ZN(o_data_bus[30]) );
  INVD15BWP30P140 U734 ( .I(n222), .ZN(o_data_bus[31]) );
  INVD15BWP30P140 U735 ( .I(n223), .ZN(o_data_bus[128]) );
  INVD15BWP30P140 U736 ( .I(n224), .ZN(o_data_bus[129]) );
  INVD15BWP30P140 U737 ( .I(n225), .ZN(o_data_bus[130]) );
  INVD15BWP30P140 U738 ( .I(n226), .ZN(o_data_bus[131]) );
  INVD15BWP30P140 U739 ( .I(n227), .ZN(o_data_bus[132]) );
  INVD15BWP30P140 U740 ( .I(n228), .ZN(o_data_bus[133]) );
  INVD15BWP30P140 U741 ( .I(n229), .ZN(o_data_bus[134]) );
  INVD15BWP30P140 U742 ( .I(n230), .ZN(o_data_bus[135]) );
  INVD15BWP30P140 U743 ( .I(n231), .ZN(o_data_bus[136]) );
  INVD15BWP30P140 U744 ( .I(n232), .ZN(o_data_bus[137]) );
  INVD15BWP30P140 U745 ( .I(n233), .ZN(o_data_bus[138]) );
  INVD15BWP30P140 U746 ( .I(n234), .ZN(o_data_bus[139]) );
  INVD15BWP30P140 U747 ( .I(n235), .ZN(o_data_bus[140]) );
  INVD15BWP30P140 U748 ( .I(n236), .ZN(o_data_bus[141]) );
  INVD15BWP30P140 U749 ( .I(n237), .ZN(o_data_bus[142]) );
  INVD15BWP30P140 U750 ( .I(n238), .ZN(o_data_bus[143]) );
  INVD15BWP30P140 U751 ( .I(n239), .ZN(o_data_bus[144]) );
  INVD15BWP30P140 U752 ( .I(n240), .ZN(o_data_bus[145]) );
  INVD15BWP30P140 U753 ( .I(n241), .ZN(o_data_bus[146]) );
  INVD15BWP30P140 U754 ( .I(n242), .ZN(o_data_bus[147]) );
  INVD15BWP30P140 U755 ( .I(n243), .ZN(o_data_bus[148]) );
  INVD15BWP30P140 U756 ( .I(n244), .ZN(o_data_bus[149]) );
  INVD15BWP30P140 U757 ( .I(n245), .ZN(o_data_bus[150]) );
  INVD15BWP30P140 U758 ( .I(n246), .ZN(o_data_bus[151]) );
  INVD15BWP30P140 U759 ( .I(n247), .ZN(o_data_bus[152]) );
  INVD15BWP30P140 U760 ( .I(n248), .ZN(o_data_bus[153]) );
  INVD15BWP30P140 U761 ( .I(n249), .ZN(o_data_bus[154]) );
  INVD15BWP30P140 U762 ( .I(n250), .ZN(o_data_bus[155]) );
  INVD15BWP30P140 U763 ( .I(n251), .ZN(o_data_bus[156]) );
  INVD15BWP30P140 U764 ( .I(n252), .ZN(o_data_bus[157]) );
  INVD15BWP30P140 U765 ( .I(n253), .ZN(o_data_bus[158]) );
  INVD15BWP30P140 U766 ( .I(n254), .ZN(o_data_bus[159]) );
  INVD15BWP30P140 U767 ( .I(n255), .ZN(o_data_bus[64]) );
  INVD15BWP30P140 U768 ( .I(n256), .ZN(o_data_bus[65]) );
  INVD15BWP30P140 U769 ( .I(n257), .ZN(o_data_bus[66]) );
  INVD15BWP30P140 U770 ( .I(n258), .ZN(o_data_bus[67]) );
  INVD15BWP30P140 U771 ( .I(n259), .ZN(o_data_bus[68]) );
  INVD15BWP30P140 U772 ( .I(n260), .ZN(o_data_bus[69]) );
  INVD15BWP30P140 U773 ( .I(n261), .ZN(o_data_bus[70]) );
  INVD15BWP30P140 U774 ( .I(n262), .ZN(o_data_bus[71]) );
  INVD15BWP30P140 U775 ( .I(n263), .ZN(o_data_bus[72]) );
  INVD15BWP30P140 U776 ( .I(n264), .ZN(o_data_bus[73]) );
  INVD15BWP30P140 U777 ( .I(n265), .ZN(o_data_bus[74]) );
  INVD15BWP30P140 U778 ( .I(n266), .ZN(o_data_bus[75]) );
  INVD15BWP30P140 U779 ( .I(n267), .ZN(o_data_bus[76]) );
  INVD15BWP30P140 U780 ( .I(n268), .ZN(o_data_bus[77]) );
  INVD15BWP30P140 U781 ( .I(n269), .ZN(o_data_bus[78]) );
  INVD15BWP30P140 U782 ( .I(n270), .ZN(o_data_bus[79]) );
  INVD15BWP30P140 U783 ( .I(n271), .ZN(o_data_bus[80]) );
  INVD15BWP30P140 U784 ( .I(n272), .ZN(o_data_bus[81]) );
  INVD15BWP30P140 U785 ( .I(n273), .ZN(o_data_bus[82]) );
  INVD15BWP30P140 U786 ( .I(n274), .ZN(o_data_bus[83]) );
  INVD15BWP30P140 U787 ( .I(n275), .ZN(o_data_bus[84]) );
  INVD15BWP30P140 U788 ( .I(n276), .ZN(o_data_bus[85]) );
  INVD15BWP30P140 U789 ( .I(n277), .ZN(o_data_bus[86]) );
  INVD15BWP30P140 U790 ( .I(n278), .ZN(o_data_bus[87]) );
  INVD15BWP30P140 U791 ( .I(n279), .ZN(o_data_bus[88]) );
  INVD15BWP30P140 U792 ( .I(n280), .ZN(o_data_bus[89]) );
  INVD15BWP30P140 U793 ( .I(n281), .ZN(o_data_bus[90]) );
  INVD15BWP30P140 U794 ( .I(n282), .ZN(o_data_bus[91]) );
  INVD15BWP30P140 U795 ( .I(n283), .ZN(o_data_bus[92]) );
  INVD15BWP30P140 U796 ( .I(n284), .ZN(o_data_bus[95]) );
  INVD15BWP30P140 U797 ( .I(n285), .ZN(o_data_bus[94]) );
  INVD15BWP30P140 U798 ( .I(n286), .ZN(o_data_bus[93]) );
  INVD15BWP30P140 U799 ( .I(n287), .ZN(o_data_bus[540]) );
  INVD15BWP30P140 U800 ( .I(n288), .ZN(o_data_bus[541]) );
  INVD15BWP30P140 U801 ( .I(n289), .ZN(o_data_bus[542]) );
  INVD15BWP30P140 U802 ( .I(n290), .ZN(o_data_bus[543]) );
  INVD15BWP30P140 U803 ( .I(n291), .ZN(o_data_bus[576]) );
  INVD15BWP30P140 U804 ( .I(n292), .ZN(o_data_bus[577]) );
  INVD15BWP30P140 U805 ( .I(n293), .ZN(o_data_bus[578]) );
  INVD15BWP30P140 U806 ( .I(n294), .ZN(o_data_bus[579]) );
  INVD15BWP30P140 U807 ( .I(n295), .ZN(o_data_bus[580]) );
  INVD15BWP30P140 U808 ( .I(n296), .ZN(o_data_bus[581]) );
  INVD15BWP30P140 U809 ( .I(n297), .ZN(o_data_bus[582]) );
  INVD15BWP30P140 U810 ( .I(n298), .ZN(o_data_bus[583]) );
  INVD15BWP30P140 U811 ( .I(n299), .ZN(o_data_bus[584]) );
  INVD15BWP30P140 U812 ( .I(n300), .ZN(o_data_bus[585]) );
  INVD15BWP30P140 U813 ( .I(n301), .ZN(o_data_bus[586]) );
  INVD15BWP30P140 U814 ( .I(n302), .ZN(o_data_bus[587]) );
  INVD15BWP30P140 U815 ( .I(n303), .ZN(o_data_bus[588]) );
  INVD15BWP30P140 U816 ( .I(n304), .ZN(o_data_bus[589]) );
  INVD15BWP30P140 U817 ( .I(n305), .ZN(o_data_bus[590]) );
  INVD15BWP30P140 U818 ( .I(n306), .ZN(o_data_bus[591]) );
  INVD15BWP30P140 U819 ( .I(n307), .ZN(o_data_bus[592]) );
  INVD15BWP30P140 U820 ( .I(n308), .ZN(o_data_bus[593]) );
  INVD15BWP30P140 U821 ( .I(n309), .ZN(o_data_bus[594]) );
  INVD15BWP30P140 U822 ( .I(n310), .ZN(o_data_bus[595]) );
  INVD15BWP30P140 U823 ( .I(n311), .ZN(o_data_bus[596]) );
  INVD15BWP30P140 U824 ( .I(n312), .ZN(o_data_bus[597]) );
  INVD15BWP30P140 U825 ( .I(n313), .ZN(o_data_bus[598]) );
  INVD15BWP30P140 U826 ( .I(n314), .ZN(o_data_bus[599]) );
  INVD15BWP30P140 U827 ( .I(n315), .ZN(o_data_bus[600]) );
  INVD15BWP30P140 U828 ( .I(n316), .ZN(o_data_bus[601]) );
  INVD15BWP30P140 U829 ( .I(n317), .ZN(o_data_bus[602]) );
  INVD15BWP30P140 U830 ( .I(n318), .ZN(o_data_bus[603]) );
  INVD15BWP30P140 U831 ( .I(n319), .ZN(o_data_bus[604]) );
  INVD15BWP30P140 U832 ( .I(n320), .ZN(o_data_bus[605]) );
  INVD15BWP30P140 U833 ( .I(n321), .ZN(o_data_bus[606]) );
  INVD15BWP30P140 U834 ( .I(n322), .ZN(o_data_bus[607]) );
  INVD15BWP30P140 U835 ( .I(n323), .ZN(o_data_bus[640]) );
  INVD15BWP30P140 U836 ( .I(n324), .ZN(o_data_bus[641]) );
  INVD15BWP30P140 U837 ( .I(n325), .ZN(o_data_bus[642]) );
  INVD15BWP30P140 U838 ( .I(n326), .ZN(o_data_bus[643]) );
  INVD15BWP30P140 U839 ( .I(n327), .ZN(o_data_bus[644]) );
  INVD15BWP30P140 U840 ( .I(n328), .ZN(o_data_bus[645]) );
  INVD15BWP30P140 U841 ( .I(n329), .ZN(o_data_bus[646]) );
  INVD15BWP30P140 U842 ( .I(n330), .ZN(o_data_bus[647]) );
  INVD15BWP30P140 U843 ( .I(n331), .ZN(o_data_bus[648]) );
  INVD15BWP30P140 U844 ( .I(n332), .ZN(o_data_bus[649]) );
  INVD15BWP30P140 U845 ( .I(n333), .ZN(o_data_bus[650]) );
  INVD15BWP30P140 U846 ( .I(n334), .ZN(o_data_bus[651]) );
  INVD15BWP30P140 U847 ( .I(n335), .ZN(o_data_bus[652]) );
  INVD15BWP30P140 U848 ( .I(n336), .ZN(o_data_bus[653]) );
  INVD15BWP30P140 U849 ( .I(n337), .ZN(o_data_bus[654]) );
  INVD15BWP30P140 U850 ( .I(n338), .ZN(o_data_bus[655]) );
  INVD15BWP30P140 U851 ( .I(n339), .ZN(o_data_bus[656]) );
  INVD15BWP30P140 U852 ( .I(n340), .ZN(o_data_bus[657]) );
  INVD15BWP30P140 U853 ( .I(n341), .ZN(o_data_bus[658]) );
  INVD15BWP30P140 U854 ( .I(n342), .ZN(o_data_bus[659]) );
  INVD15BWP30P140 U855 ( .I(n343), .ZN(o_data_bus[660]) );
  INVD15BWP30P140 U856 ( .I(n344), .ZN(o_data_bus[661]) );
  INVD15BWP30P140 U857 ( .I(n345), .ZN(o_data_bus[662]) );
  INVD15BWP30P140 U858 ( .I(n346), .ZN(o_data_bus[663]) );
  INVD15BWP30P140 U859 ( .I(n347), .ZN(o_data_bus[664]) );
  INVD15BWP30P140 U860 ( .I(n348), .ZN(o_data_bus[665]) );
  INVD15BWP30P140 U861 ( .I(n349), .ZN(o_data_bus[666]) );
  INVD15BWP30P140 U862 ( .I(n350), .ZN(o_data_bus[667]) );
  INVD15BWP30P140 U863 ( .I(n351), .ZN(o_data_bus[668]) );
  INVD15BWP30P140 U864 ( .I(n352), .ZN(o_data_bus[669]) );
  INVD15BWP30P140 U865 ( .I(n353), .ZN(o_data_bus[670]) );
  INVD15BWP30P140 U866 ( .I(n354), .ZN(o_data_bus[671]) );
  INVD15BWP30P140 U867 ( .I(n355), .ZN(o_data_bus[704]) );
  INVD15BWP30P140 U868 ( .I(n356), .ZN(o_data_bus[705]) );
  INVD15BWP30P140 U869 ( .I(n357), .ZN(o_data_bus[706]) );
  INVD15BWP30P140 U870 ( .I(n358), .ZN(o_data_bus[707]) );
  INVD15BWP30P140 U871 ( .I(n359), .ZN(o_data_bus[708]) );
  INVD15BWP30P140 U872 ( .I(n360), .ZN(o_data_bus[709]) );
  INVD15BWP30P140 U873 ( .I(n361), .ZN(o_data_bus[710]) );
  INVD15BWP30P140 U874 ( .I(n362), .ZN(o_data_bus[711]) );
  INVD15BWP30P140 U875 ( .I(n363), .ZN(o_data_bus[712]) );
  INVD15BWP30P140 U876 ( .I(n364), .ZN(o_data_bus[713]) );
  INVD15BWP30P140 U877 ( .I(n365), .ZN(o_data_bus[714]) );
  INVD15BWP30P140 U878 ( .I(n366), .ZN(o_data_bus[715]) );
  INVD15BWP30P140 U879 ( .I(n367), .ZN(o_data_bus[716]) );
  INVD15BWP30P140 U880 ( .I(n368), .ZN(o_data_bus[717]) );
  INVD15BWP30P140 U881 ( .I(n369), .ZN(o_data_bus[718]) );
  INVD15BWP30P140 U882 ( .I(n370), .ZN(o_data_bus[719]) );
  INVD15BWP30P140 U883 ( .I(n371), .ZN(o_data_bus[720]) );
  INVD15BWP30P140 U884 ( .I(n372), .ZN(o_data_bus[721]) );
  INVD15BWP30P140 U885 ( .I(n373), .ZN(o_data_bus[722]) );
  INVD15BWP30P140 U886 ( .I(n374), .ZN(o_data_bus[723]) );
  INVD15BWP30P140 U887 ( .I(n375), .ZN(o_data_bus[724]) );
  INVD15BWP30P140 U888 ( .I(n376), .ZN(o_data_bus[725]) );
  INVD15BWP30P140 U889 ( .I(n377), .ZN(o_data_bus[726]) );
  INVD15BWP30P140 U890 ( .I(n378), .ZN(o_data_bus[727]) );
  INVD15BWP30P140 U891 ( .I(n379), .ZN(o_data_bus[728]) );
  INVD15BWP30P140 U892 ( .I(n380), .ZN(o_data_bus[729]) );
  INVD15BWP30P140 U893 ( .I(n381), .ZN(o_data_bus[730]) );
  INVD15BWP30P140 U894 ( .I(n382), .ZN(o_data_bus[731]) );
  INVD15BWP30P140 U895 ( .I(n383), .ZN(o_data_bus[732]) );
  INVD15BWP30P140 U896 ( .I(n384), .ZN(o_data_bus[733]) );
  INVD15BWP30P140 U897 ( .I(n385), .ZN(o_data_bus[734]) );
  INVD15BWP30P140 U898 ( .I(n386), .ZN(o_data_bus[735]) );
  INVD15BWP30P140 U899 ( .I(n387), .ZN(o_data_bus[768]) );
  INVD15BWP30P140 U900 ( .I(n388), .ZN(o_data_bus[769]) );
  INVD15BWP30P140 U901 ( .I(n389), .ZN(o_data_bus[770]) );
  INVD15BWP30P140 U902 ( .I(n390), .ZN(o_data_bus[771]) );
  INVD15BWP30P140 U903 ( .I(n391), .ZN(o_data_bus[772]) );
  INVD15BWP30P140 U904 ( .I(n392), .ZN(o_data_bus[773]) );
  INVD15BWP30P140 U905 ( .I(n393), .ZN(o_data_bus[774]) );
  INVD15BWP30P140 U906 ( .I(n394), .ZN(o_data_bus[775]) );
  INVD15BWP30P140 U907 ( .I(n395), .ZN(o_data_bus[776]) );
  INVD15BWP30P140 U908 ( .I(n396), .ZN(o_data_bus[777]) );
  INVD15BWP30P140 U909 ( .I(n397), .ZN(o_data_bus[778]) );
  INVD15BWP30P140 U910 ( .I(n398), .ZN(o_data_bus[779]) );
  INVD15BWP30P140 U911 ( .I(n399), .ZN(o_data_bus[780]) );
  INVD15BWP30P140 U912 ( .I(n400), .ZN(o_data_bus[781]) );
  INVD15BWP30P140 U913 ( .I(n401), .ZN(o_data_bus[782]) );
  INVD15BWP30P140 U914 ( .I(n402), .ZN(o_data_bus[783]) );
  INVD15BWP30P140 U915 ( .I(n403), .ZN(o_data_bus[784]) );
  INVD15BWP30P140 U916 ( .I(n404), .ZN(o_data_bus[785]) );
  INVD15BWP30P140 U917 ( .I(n405), .ZN(o_data_bus[786]) );
  INVD15BWP30P140 U918 ( .I(n406), .ZN(o_data_bus[787]) );
  INVD15BWP30P140 U919 ( .I(n407), .ZN(o_data_bus[788]) );
  INVD15BWP30P140 U920 ( .I(n408), .ZN(o_data_bus[789]) );
  INVD15BWP30P140 U921 ( .I(n409), .ZN(o_data_bus[790]) );
  INVD15BWP30P140 U922 ( .I(n410), .ZN(o_data_bus[791]) );
  INVD15BWP30P140 U923 ( .I(n411), .ZN(o_data_bus[792]) );
  INVD15BWP30P140 U924 ( .I(n412), .ZN(o_data_bus[793]) );
  INVD15BWP30P140 U925 ( .I(n413), .ZN(o_data_bus[794]) );
  INVD15BWP30P140 U926 ( .I(n414), .ZN(o_data_bus[795]) );
  INVD15BWP30P140 U927 ( .I(n415), .ZN(o_data_bus[796]) );
  INVD15BWP30P140 U928 ( .I(n416), .ZN(o_data_bus[797]) );
  INVD15BWP30P140 U929 ( .I(n417), .ZN(o_data_bus[798]) );
  INVD15BWP30P140 U930 ( .I(n418), .ZN(o_data_bus[799]) );
  INVD15BWP30P140 U931 ( .I(n419), .ZN(o_data_bus[832]) );
  INVD15BWP30P140 U932 ( .I(n420), .ZN(o_data_bus[833]) );
  INVD15BWP30P140 U933 ( .I(n421), .ZN(o_data_bus[834]) );
  INVD15BWP30P140 U934 ( .I(n422), .ZN(o_data_bus[835]) );
  INVD15BWP30P140 U935 ( .I(n423), .ZN(o_data_bus[836]) );
  INVD15BWP30P140 U936 ( .I(n424), .ZN(o_data_bus[837]) );
  INVD15BWP30P140 U937 ( .I(n425), .ZN(o_data_bus[838]) );
  INVD15BWP30P140 U938 ( .I(n426), .ZN(o_data_bus[839]) );
  INVD15BWP30P140 U939 ( .I(n427), .ZN(o_data_bus[840]) );
  INVD15BWP30P140 U940 ( .I(n428), .ZN(o_data_bus[841]) );
  INVD15BWP30P140 U941 ( .I(n429), .ZN(o_data_bus[842]) );
  INVD15BWP30P140 U942 ( .I(n430), .ZN(o_data_bus[843]) );
  INVD15BWP30P140 U943 ( .I(n431), .ZN(o_data_bus[844]) );
  INVD15BWP30P140 U944 ( .I(n432), .ZN(o_data_bus[845]) );
  INVD15BWP30P140 U945 ( .I(n433), .ZN(o_data_bus[846]) );
  INVD15BWP30P140 U946 ( .I(n434), .ZN(o_data_bus[847]) );
  INVD15BWP30P140 U947 ( .I(n435), .ZN(o_data_bus[848]) );
  INVD15BWP30P140 U948 ( .I(n436), .ZN(o_data_bus[849]) );
  INVD15BWP30P140 U949 ( .I(n437), .ZN(o_data_bus[850]) );
  INVD15BWP30P140 U950 ( .I(n438), .ZN(o_data_bus[851]) );
  INVD15BWP30P140 U951 ( .I(n439), .ZN(o_data_bus[852]) );
  INVD15BWP30P140 U952 ( .I(n440), .ZN(o_data_bus[853]) );
  INVD15BWP30P140 U953 ( .I(n441), .ZN(o_data_bus[854]) );
  INVD15BWP30P140 U954 ( .I(n442), .ZN(o_data_bus[855]) );
  INVD15BWP30P140 U955 ( .I(n443), .ZN(o_data_bus[856]) );
  INVD15BWP30P140 U956 ( .I(n444), .ZN(o_data_bus[857]) );
  INVD15BWP30P140 U957 ( .I(n445), .ZN(o_data_bus[858]) );
  INVD15BWP30P140 U958 ( .I(n446), .ZN(o_data_bus[859]) );
  INVD15BWP30P140 U959 ( .I(n447), .ZN(o_data_bus[860]) );
  INVD15BWP30P140 U960 ( .I(n448), .ZN(o_data_bus[861]) );
  INVD15BWP30P140 U961 ( .I(n449), .ZN(o_data_bus[862]) );
  INVD15BWP30P140 U962 ( .I(n450), .ZN(o_data_bus[863]) );
  INVD15BWP30P140 U963 ( .I(n451), .ZN(o_data_bus[896]) );
  INVD15BWP30P140 U964 ( .I(n452), .ZN(o_data_bus[897]) );
  INVD15BWP30P140 U965 ( .I(n453), .ZN(o_data_bus[898]) );
  INVD15BWP30P140 U966 ( .I(n454), .ZN(o_data_bus[899]) );
  INVD15BWP30P140 U967 ( .I(n455), .ZN(o_data_bus[900]) );
  INVD15BWP30P140 U968 ( .I(n456), .ZN(o_data_bus[901]) );
  INVD15BWP30P140 U969 ( .I(n457), .ZN(o_data_bus[902]) );
  INVD15BWP30P140 U970 ( .I(n458), .ZN(o_data_bus[903]) );
  INVD15BWP30P140 U971 ( .I(n459), .ZN(o_data_bus[904]) );
  INVD15BWP30P140 U972 ( .I(n460), .ZN(o_data_bus[905]) );
  INVD15BWP30P140 U973 ( .I(n461), .ZN(o_data_bus[906]) );
  INVD15BWP30P140 U974 ( .I(n462), .ZN(o_data_bus[907]) );
  INVD15BWP30P140 U975 ( .I(n463), .ZN(o_data_bus[908]) );
  INVD15BWP30P140 U976 ( .I(n464), .ZN(o_data_bus[909]) );
  INVD15BWP30P140 U977 ( .I(n465), .ZN(o_data_bus[910]) );
  INVD15BWP30P140 U978 ( .I(n466), .ZN(o_data_bus[911]) );
  INVD15BWP30P140 U979 ( .I(n467), .ZN(o_data_bus[912]) );
  INVD15BWP30P140 U980 ( .I(n468), .ZN(o_data_bus[913]) );
  INVD15BWP30P140 U981 ( .I(n469), .ZN(o_data_bus[914]) );
  INVD15BWP30P140 U982 ( .I(n470), .ZN(o_data_bus[915]) );
  INVD15BWP30P140 U983 ( .I(n471), .ZN(o_data_bus[916]) );
  INVD15BWP30P140 U984 ( .I(n472), .ZN(o_data_bus[917]) );
  INVD15BWP30P140 U985 ( .I(n473), .ZN(o_data_bus[918]) );
  INVD15BWP30P140 U986 ( .I(n474), .ZN(o_data_bus[919]) );
  INVD15BWP30P140 U987 ( .I(n475), .ZN(o_data_bus[920]) );
  INVD15BWP30P140 U988 ( .I(n476), .ZN(o_data_bus[921]) );
  INVD15BWP30P140 U989 ( .I(n477), .ZN(o_data_bus[922]) );
  INVD15BWP30P140 U990 ( .I(n478), .ZN(o_data_bus[923]) );
  INVD15BWP30P140 U991 ( .I(n479), .ZN(o_data_bus[924]) );
  INVD15BWP30P140 U992 ( .I(n480), .ZN(o_data_bus[925]) );
  INVD15BWP30P140 U993 ( .I(n481), .ZN(o_data_bus[926]) );
  INVD15BWP30P140 U994 ( .I(n482), .ZN(o_data_bus[927]) );
  INVD12BWP30P140 U995 ( .I(n483), .ZN(o_data_bus[960]) );
  INVD12BWP30P140 U996 ( .I(n484), .ZN(o_data_bus[961]) );
  INVD12BWP30P140 U997 ( .I(n485), .ZN(o_data_bus[962]) );
  INVD12BWP30P140 U998 ( .I(n486), .ZN(o_data_bus[963]) );
  INVD12BWP30P140 U999 ( .I(n487), .ZN(o_data_bus[964]) );
  INVD12BWP30P140 U1000 ( .I(n488), .ZN(o_data_bus[965]) );
  INVD12BWP30P140 U1001 ( .I(n489), .ZN(o_data_bus[966]) );
  INVD12BWP30P140 U1002 ( .I(n490), .ZN(o_data_bus[967]) );
  INVD12BWP30P140 U1003 ( .I(n491), .ZN(o_data_bus[968]) );
  INVD12BWP30P140 U1004 ( .I(n492), .ZN(o_data_bus[969]) );
  INVD12BWP30P140 U1005 ( .I(n493), .ZN(o_data_bus[970]) );
  INVD12BWP30P140 U1006 ( .I(n494), .ZN(o_data_bus[971]) );
  INVD12BWP30P140 U1007 ( .I(n495), .ZN(o_data_bus[972]) );
  INVD12BWP30P140 U1008 ( .I(n496), .ZN(o_data_bus[973]) );
  INVD12BWP30P140 U1009 ( .I(n497), .ZN(o_data_bus[974]) );
  INVD12BWP30P140 U1010 ( .I(n498), .ZN(o_data_bus[975]) );
  INVD12BWP30P140 U1011 ( .I(n499), .ZN(o_data_bus[976]) );
  INVD12BWP30P140 U1012 ( .I(n500), .ZN(o_data_bus[977]) );
  INVD12BWP30P140 U1013 ( .I(n501), .ZN(o_data_bus[978]) );
  INVD12BWP30P140 U1014 ( .I(n502), .ZN(o_data_bus[979]) );
  INVD12BWP30P140 U1015 ( .I(n503), .ZN(o_data_bus[980]) );
  INVD12BWP30P140 U1016 ( .I(n504), .ZN(o_data_bus[981]) );
  INVD12BWP30P140 U1017 ( .I(n505), .ZN(o_data_bus[982]) );
  INVD12BWP30P140 U1018 ( .I(n506), .ZN(o_data_bus[983]) );
  INVD12BWP30P140 U1019 ( .I(n507), .ZN(o_data_bus[984]) );
  INVD12BWP30P140 U1020 ( .I(n508), .ZN(o_data_bus[985]) );
  INVD12BWP30P140 U1021 ( .I(n509), .ZN(o_data_bus[986]) );
  INVD12BWP30P140 U1022 ( .I(n510), .ZN(o_data_bus[987]) );
  INVD12BWP30P140 U1023 ( .I(n511), .ZN(o_data_bus[988]) );
  INVD12BWP30P140 U1024 ( .I(n512), .ZN(o_data_bus[989]) );
  BUFFD12BWP30P140 U1025 ( .I(n2600), .Z(o_data_bus[40]) );
  BUFFD12BWP30P140 U1026 ( .I(n2599), .Z(o_data_bus[41]) );
  BUFFD12BWP30P140 U1027 ( .I(n2598), .Z(o_data_bus[42]) );
  BUFFD12BWP30P140 U1028 ( .I(n2597), .Z(o_data_bus[43]) );
  BUFFD12BWP30P140 U1029 ( .I(n2596), .Z(o_data_bus[44]) );
  BUFFD12BWP30P140 U1030 ( .I(n2595), .Z(o_data_bus[45]) );
  BUFFD12BWP30P140 U1031 ( .I(n2594), .Z(o_data_bus[46]) );
  BUFFD12BWP30P140 U1032 ( .I(n2593), .Z(o_data_bus[47]) );
  BUFFD12BWP30P140 U1033 ( .I(n2592), .Z(o_data_bus[48]) );
  BUFFD12BWP30P140 U1034 ( .I(n2591), .Z(o_data_bus[49]) );
  BUFFD12BWP30P140 U1035 ( .I(n2590), .Z(o_data_bus[50]) );
  BUFFD12BWP30P140 U1036 ( .I(n2589), .Z(o_data_bus[51]) );
  BUFFD12BWP30P140 U1037 ( .I(n2588), .Z(o_data_bus[52]) );
  BUFFD12BWP30P140 U1038 ( .I(n2587), .Z(o_data_bus[53]) );
  BUFFD12BWP30P140 U1039 ( .I(n2586), .Z(o_data_bus[54]) );
  BUFFD12BWP30P140 U1040 ( .I(n2585), .Z(o_data_bus[55]) );
  BUFFD12BWP30P140 U1041 ( .I(n2584), .Z(o_data_bus[56]) );
  BUFFD12BWP30P140 U1042 ( .I(n2583), .Z(o_data_bus[57]) );
  BUFFD12BWP30P140 U1043 ( .I(n2582), .Z(o_data_bus[58]) );
  BUFFD12BWP30P140 U1044 ( .I(n2581), .Z(o_data_bus[59]) );
  BUFFD12BWP30P140 U1045 ( .I(n2580), .Z(o_data_bus[60]) );
  BUFFD12BWP30P140 U1046 ( .I(n2579), .Z(o_data_bus[61]) );
  BUFFD12BWP30P140 U1047 ( .I(n2578), .Z(o_data_bus[62]) );
  BUFFD12BWP30P140 U1048 ( .I(n2577), .Z(o_data_bus[63]) );
  BUFFD12BWP30P140 U1049 ( .I(n2536), .Z(o_data_bus[104]) );
  BUFFD12BWP30P140 U1050 ( .I(n2535), .Z(o_data_bus[105]) );
  BUFFD12BWP30P140 U1051 ( .I(n2534), .Z(o_data_bus[106]) );
  BUFFD12BWP30P140 U1052 ( .I(n2533), .Z(o_data_bus[107]) );
  BUFFD12BWP30P140 U1053 ( .I(n2532), .Z(o_data_bus[108]) );
  BUFFD12BWP30P140 U1054 ( .I(n2531), .Z(o_data_bus[109]) );
  BUFFD12BWP30P140 U1055 ( .I(n2530), .Z(o_data_bus[110]) );
  BUFFD12BWP30P140 U1056 ( .I(n2529), .Z(o_data_bus[111]) );
  BUFFD12BWP30P140 U1057 ( .I(n2528), .Z(o_data_bus[112]) );
  BUFFD12BWP30P140 U1058 ( .I(n2527), .Z(o_data_bus[113]) );
  BUFFD12BWP30P140 U1059 ( .I(n2526), .Z(o_data_bus[114]) );
  BUFFD12BWP30P140 U1060 ( .I(n2525), .Z(o_data_bus[115]) );
  BUFFD12BWP30P140 U1061 ( .I(n2524), .Z(o_data_bus[116]) );
  BUFFD12BWP30P140 U1062 ( .I(n2523), .Z(o_data_bus[117]) );
  BUFFD12BWP30P140 U1063 ( .I(n2522), .Z(o_data_bus[118]) );
  BUFFD12BWP30P140 U1064 ( .I(n2521), .Z(o_data_bus[119]) );
  BUFFD12BWP30P140 U1065 ( .I(n2520), .Z(o_data_bus[120]) );
  BUFFD12BWP30P140 U1066 ( .I(n2519), .Z(o_data_bus[121]) );
  BUFFD12BWP30P140 U1067 ( .I(n2518), .Z(o_data_bus[122]) );
  BUFFD12BWP30P140 U1068 ( .I(n2517), .Z(o_data_bus[123]) );
  BUFFD12BWP30P140 U1069 ( .I(n2516), .Z(o_data_bus[124]) );
  BUFFD12BWP30P140 U1070 ( .I(n2515), .Z(o_data_bus[125]) );
  BUFFD12BWP30P140 U1071 ( .I(n2514), .Z(o_data_bus[126]) );
  BUFFD12BWP30P140 U1072 ( .I(n2513), .Z(o_data_bus[127]) );
  BUFFD12BWP30P140 U1073 ( .I(n2472), .Z(o_data_bus[168]) );
  BUFFD12BWP30P140 U1074 ( .I(n2471), .Z(o_data_bus[169]) );
  BUFFD12BWP30P140 U1075 ( .I(n2470), .Z(o_data_bus[170]) );
  BUFFD12BWP30P140 U1076 ( .I(n2469), .Z(o_data_bus[171]) );
  BUFFD12BWP30P140 U1077 ( .I(n2468), .Z(o_data_bus[172]) );
  BUFFD12BWP30P140 U1078 ( .I(n2467), .Z(o_data_bus[173]) );
  BUFFD12BWP30P140 U1079 ( .I(n2466), .Z(o_data_bus[174]) );
  BUFFD12BWP30P140 U1080 ( .I(n2465), .Z(o_data_bus[175]) );
  BUFFD12BWP30P140 U1081 ( .I(n2464), .Z(o_data_bus[176]) );
  BUFFD12BWP30P140 U1082 ( .I(n2463), .Z(o_data_bus[177]) );
  BUFFD12BWP30P140 U1083 ( .I(n2462), .Z(o_data_bus[178]) );
  BUFFD12BWP30P140 U1084 ( .I(n2461), .Z(o_data_bus[179]) );
  BUFFD12BWP30P140 U1085 ( .I(n2460), .Z(o_data_bus[180]) );
  BUFFD12BWP30P140 U1086 ( .I(n2459), .Z(o_data_bus[181]) );
  BUFFD12BWP30P140 U1087 ( .I(n2458), .Z(o_data_bus[182]) );
  BUFFD12BWP30P140 U1088 ( .I(n2457), .Z(o_data_bus[183]) );
  BUFFD12BWP30P140 U1089 ( .I(n2456), .Z(o_data_bus[184]) );
  BUFFD12BWP30P140 U1090 ( .I(n2455), .Z(o_data_bus[185]) );
  BUFFD12BWP30P140 U1091 ( .I(n2454), .Z(o_data_bus[186]) );
  BUFFD12BWP30P140 U1092 ( .I(n2453), .Z(o_data_bus[187]) );
  BUFFD12BWP30P140 U1093 ( .I(n2452), .Z(o_data_bus[188]) );
  BUFFD12BWP30P140 U1094 ( .I(n2451), .Z(o_data_bus[189]) );
  BUFFD12BWP30P140 U1095 ( .I(n2450), .Z(o_data_bus[190]) );
  BUFFD12BWP30P140 U1096 ( .I(n2449), .Z(o_data_bus[191]) );
  BUFFD12BWP30P140 U1097 ( .I(n2408), .Z(o_data_bus[232]) );
  BUFFD12BWP30P140 U1098 ( .I(n2407), .Z(o_data_bus[233]) );
  BUFFD12BWP30P140 U1099 ( .I(n2406), .Z(o_data_bus[234]) );
  BUFFD12BWP30P140 U1100 ( .I(n2405), .Z(o_data_bus[235]) );
  BUFFD12BWP30P140 U1101 ( .I(n2404), .Z(o_data_bus[236]) );
  BUFFD12BWP30P140 U1102 ( .I(n2403), .Z(o_data_bus[237]) );
  BUFFD12BWP30P140 U1103 ( .I(n2402), .Z(o_data_bus[238]) );
  BUFFD12BWP30P140 U1104 ( .I(n2401), .Z(o_data_bus[239]) );
  BUFFD12BWP30P140 U1105 ( .I(n2400), .Z(o_data_bus[240]) );
  BUFFD12BWP30P140 U1106 ( .I(n2399), .Z(o_data_bus[241]) );
  BUFFD12BWP30P140 U1107 ( .I(n2398), .Z(o_data_bus[242]) );
  BUFFD12BWP30P140 U1108 ( .I(n2397), .Z(o_data_bus[243]) );
  BUFFD12BWP30P140 U1109 ( .I(n2396), .Z(o_data_bus[244]) );
  BUFFD12BWP30P140 U1110 ( .I(n2395), .Z(o_data_bus[245]) );
  BUFFD12BWP30P140 U1111 ( .I(n2394), .Z(o_data_bus[246]) );
  BUFFD12BWP30P140 U1112 ( .I(n2393), .Z(o_data_bus[247]) );
  BUFFD12BWP30P140 U1113 ( .I(n2392), .Z(o_data_bus[248]) );
  BUFFD12BWP30P140 U1114 ( .I(n2391), .Z(o_data_bus[249]) );
  BUFFD12BWP30P140 U1115 ( .I(n2390), .Z(o_data_bus[250]) );
  BUFFD12BWP30P140 U1116 ( .I(n2389), .Z(o_data_bus[251]) );
  BUFFD12BWP30P140 U1117 ( .I(n2388), .Z(o_data_bus[252]) );
  BUFFD12BWP30P140 U1118 ( .I(n2387), .Z(o_data_bus[253]) );
  BUFFD12BWP30P140 U1119 ( .I(n2386), .Z(o_data_bus[254]) );
  BUFFD12BWP30P140 U1120 ( .I(n2385), .Z(o_data_bus[255]) );
  BUFFD12BWP30P140 U1121 ( .I(n2344), .Z(o_data_bus[296]) );
  BUFFD12BWP30P140 U1122 ( .I(n2343), .Z(o_data_bus[297]) );
  BUFFD12BWP30P140 U1123 ( .I(n2342), .Z(o_data_bus[298]) );
  BUFFD12BWP30P140 U1124 ( .I(n2341), .Z(o_data_bus[299]) );
  BUFFD12BWP30P140 U1125 ( .I(n2340), .Z(o_data_bus[300]) );
  BUFFD12BWP30P140 U1126 ( .I(n2339), .Z(o_data_bus[301]) );
  BUFFD12BWP30P140 U1127 ( .I(n2338), .Z(o_data_bus[302]) );
  BUFFD12BWP30P140 U1128 ( .I(n2337), .Z(o_data_bus[303]) );
  BUFFD12BWP30P140 U1129 ( .I(n2336), .Z(o_data_bus[304]) );
  BUFFD12BWP30P140 U1130 ( .I(n2335), .Z(o_data_bus[305]) );
  BUFFD12BWP30P140 U1131 ( .I(n2334), .Z(o_data_bus[306]) );
  BUFFD12BWP30P140 U1132 ( .I(n2333), .Z(o_data_bus[307]) );
  BUFFD12BWP30P140 U1133 ( .I(n2332), .Z(o_data_bus[308]) );
  BUFFD12BWP30P140 U1134 ( .I(n2331), .Z(o_data_bus[309]) );
  BUFFD12BWP30P140 U1135 ( .I(n2330), .Z(o_data_bus[310]) );
  BUFFD12BWP30P140 U1136 ( .I(n2329), .Z(o_data_bus[311]) );
  BUFFD12BWP30P140 U1137 ( .I(n2328), .Z(o_data_bus[312]) );
  BUFFD12BWP30P140 U1138 ( .I(n2327), .Z(o_data_bus[313]) );
  BUFFD12BWP30P140 U1139 ( .I(n2326), .Z(o_data_bus[314]) );
  BUFFD12BWP30P140 U1140 ( .I(n2325), .Z(o_data_bus[315]) );
  BUFFD12BWP30P140 U1141 ( .I(n2324), .Z(o_data_bus[316]) );
  BUFFD12BWP30P140 U1142 ( .I(n2323), .Z(o_data_bus[317]) );
  BUFFD12BWP30P140 U1143 ( .I(n2322), .Z(o_data_bus[318]) );
  BUFFD12BWP30P140 U1144 ( .I(n2321), .Z(o_data_bus[319]) );
  BUFFD12BWP30P140 U1145 ( .I(n2280), .Z(o_data_bus[360]) );
  BUFFD12BWP30P140 U1146 ( .I(n2279), .Z(o_data_bus[361]) );
  BUFFD12BWP30P140 U1147 ( .I(n2278), .Z(o_data_bus[362]) );
  BUFFD12BWP30P140 U1148 ( .I(n2277), .Z(o_data_bus[363]) );
  BUFFD12BWP30P140 U1149 ( .I(n2276), .Z(o_data_bus[364]) );
  BUFFD12BWP30P140 U1150 ( .I(n2275), .Z(o_data_bus[365]) );
  BUFFD12BWP30P140 U1151 ( .I(n2274), .Z(o_data_bus[366]) );
  BUFFD12BWP30P140 U1152 ( .I(n2273), .Z(o_data_bus[367]) );
  BUFFD12BWP30P140 U1153 ( .I(n2272), .Z(o_data_bus[368]) );
  BUFFD12BWP30P140 U1154 ( .I(n2271), .Z(o_data_bus[369]) );
  BUFFD12BWP30P140 U1155 ( .I(n2270), .Z(o_data_bus[370]) );
  BUFFD12BWP30P140 U1156 ( .I(n2269), .Z(o_data_bus[371]) );
  BUFFD12BWP30P140 U1157 ( .I(n2268), .Z(o_data_bus[372]) );
  BUFFD12BWP30P140 U1158 ( .I(n2267), .Z(o_data_bus[373]) );
  BUFFD12BWP30P140 U1159 ( .I(n2266), .Z(o_data_bus[374]) );
  BUFFD12BWP30P140 U1160 ( .I(n2265), .Z(o_data_bus[375]) );
  BUFFD12BWP30P140 U1161 ( .I(n2264), .Z(o_data_bus[376]) );
  BUFFD12BWP30P140 U1162 ( .I(n2263), .Z(o_data_bus[377]) );
  BUFFD12BWP30P140 U1163 ( .I(n2262), .Z(o_data_bus[378]) );
  BUFFD12BWP30P140 U1164 ( .I(n2261), .Z(o_data_bus[379]) );
  BUFFD12BWP30P140 U1165 ( .I(n2260), .Z(o_data_bus[380]) );
  BUFFD12BWP30P140 U1166 ( .I(n2259), .Z(o_data_bus[381]) );
  BUFFD12BWP30P140 U1167 ( .I(n2258), .Z(o_data_bus[382]) );
  BUFFD12BWP30P140 U1168 ( .I(n2257), .Z(o_data_bus[383]) );
  BUFFD12BWP30P140 U1169 ( .I(n2216), .Z(o_data_bus[424]) );
  BUFFD12BWP30P140 U1170 ( .I(n2215), .Z(o_data_bus[425]) );
  BUFFD12BWP30P140 U1171 ( .I(n2214), .Z(o_data_bus[426]) );
  BUFFD12BWP30P140 U1172 ( .I(n2213), .Z(o_data_bus[427]) );
  BUFFD12BWP30P140 U1173 ( .I(n2212), .Z(o_data_bus[428]) );
  BUFFD12BWP30P140 U1174 ( .I(n2211), .Z(o_data_bus[429]) );
  BUFFD12BWP30P140 U1175 ( .I(n2210), .Z(o_data_bus[430]) );
  BUFFD12BWP30P140 U1176 ( .I(n2209), .Z(o_data_bus[431]) );
  BUFFD12BWP30P140 U1177 ( .I(n2208), .Z(o_data_bus[432]) );
  BUFFD12BWP30P140 U1178 ( .I(n2207), .Z(o_data_bus[433]) );
  BUFFD12BWP30P140 U1179 ( .I(n2206), .Z(o_data_bus[434]) );
  BUFFD12BWP30P140 U1180 ( .I(n2205), .Z(o_data_bus[435]) );
  BUFFD12BWP30P140 U1181 ( .I(n2204), .Z(o_data_bus[436]) );
  BUFFD12BWP30P140 U1182 ( .I(n2203), .Z(o_data_bus[437]) );
  BUFFD12BWP30P140 U1183 ( .I(n2202), .Z(o_data_bus[438]) );
  BUFFD12BWP30P140 U1184 ( .I(n2201), .Z(o_data_bus[439]) );
  BUFFD12BWP30P140 U1185 ( .I(n2200), .Z(o_data_bus[440]) );
  BUFFD12BWP30P140 U1186 ( .I(n2199), .Z(o_data_bus[441]) );
  BUFFD12BWP30P140 U1187 ( .I(n2198), .Z(o_data_bus[442]) );
  BUFFD12BWP30P140 U1188 ( .I(n2197), .Z(o_data_bus[443]) );
  BUFFD12BWP30P140 U1189 ( .I(n2196), .Z(o_data_bus[444]) );
  BUFFD12BWP30P140 U1190 ( .I(n2195), .Z(o_data_bus[445]) );
  BUFFD12BWP30P140 U1191 ( .I(n2194), .Z(o_data_bus[446]) );
  BUFFD12BWP30P140 U1192 ( .I(n2193), .Z(o_data_bus[447]) );
  BUFFD12BWP30P140 U1193 ( .I(n2152), .Z(o_data_bus[488]) );
  BUFFD12BWP30P140 U1194 ( .I(n2151), .Z(o_data_bus[489]) );
  BUFFD12BWP30P140 U1195 ( .I(n2150), .Z(o_data_bus[490]) );
  BUFFD12BWP30P140 U1196 ( .I(n2149), .Z(o_data_bus[491]) );
  BUFFD12BWP30P140 U1197 ( .I(n2148), .Z(o_data_bus[492]) );
  BUFFD12BWP30P140 U1198 ( .I(n2147), .Z(o_data_bus[493]) );
  BUFFD12BWP30P140 U1199 ( .I(n2146), .Z(o_data_bus[494]) );
  BUFFD12BWP30P140 U1200 ( .I(n2145), .Z(o_data_bus[495]) );
  BUFFD12BWP30P140 U1201 ( .I(n2144), .Z(o_data_bus[496]) );
  BUFFD12BWP30P140 U1202 ( .I(n2143), .Z(o_data_bus[497]) );
  BUFFD12BWP30P140 U1203 ( .I(n2142), .Z(o_data_bus[498]) );
  BUFFD12BWP30P140 U1204 ( .I(n2141), .Z(o_data_bus[499]) );
  BUFFD12BWP30P140 U1205 ( .I(n2140), .Z(o_data_bus[500]) );
  BUFFD12BWP30P140 U1206 ( .I(n2139), .Z(o_data_bus[501]) );
  BUFFD12BWP30P140 U1207 ( .I(n2138), .Z(o_data_bus[502]) );
  BUFFD12BWP30P140 U1208 ( .I(n2137), .Z(o_data_bus[503]) );
  BUFFD12BWP30P140 U1209 ( .I(n2136), .Z(o_data_bus[504]) );
  BUFFD12BWP30P140 U1210 ( .I(n2135), .Z(o_data_bus[505]) );
  BUFFD12BWP30P140 U1211 ( .I(n2134), .Z(o_data_bus[506]) );
  BUFFD12BWP30P140 U1212 ( .I(n2133), .Z(o_data_bus[507]) );
  BUFFD12BWP30P140 U1213 ( .I(n2132), .Z(o_data_bus[508]) );
  BUFFD12BWP30P140 U1214 ( .I(n2131), .Z(o_data_bus[509]) );
  BUFFD12BWP30P140 U1215 ( .I(n2130), .Z(o_data_bus[510]) );
  BUFFD12BWP30P140 U1216 ( .I(n2129), .Z(o_data_bus[511]) );
  INVD12BWP30P140 U1217 ( .I(n1547), .ZN(o_valid[7]) );
  INVD12BWP30P140 U1218 ( .I(n1538), .ZN(o_valid[1]) );
  INVD12BWP30P140 U1219 ( .I(n1553), .ZN(o_valid[11]) );
  INVD12BWP30P140 U1220 ( .I(n1550), .ZN(o_valid[9]) );
  INVD12BWP30P140 U1221 ( .I(n1580), .ZN(o_valid[29]) );
  INVD12BWP30P140 U1222 ( .I(n1577), .ZN(o_valid[27]) );
  INVD12BWP30P140 U1223 ( .I(n1574), .ZN(o_valid[25]) );
  INVD12BWP30P140 U1224 ( .I(n1544), .ZN(o_valid[5]) );
  INVD12BWP30P140 U1225 ( .I(n1541), .ZN(o_valid[3]) );
  INVD12BWP30P140 U1226 ( .I(n1568), .ZN(o_valid[21]) );
  INVD12BWP30P140 U1227 ( .I(n1565), .ZN(o_valid[19]) );
  INVD12BWP30P140 U1228 ( .I(n1562), .ZN(o_valid[17]) );
  INVD12BWP30P140 U1229 ( .I(n1559), .ZN(o_valid[15]) );
  INVD12BWP30P140 U1230 ( .I(n1556), .ZN(o_valid[13]) );
  INVD12BWP30P140 U1231 ( .I(n1571), .ZN(o_valid[23]) );
  INVD12BWP30P140 U1232 ( .I(n1583), .ZN(o_valid[31]) );
  BUFFD12BWP30P140 U1233 ( .I(n2409), .Z(o_data_bus[231]) );
  BUFFD12BWP30P140 U1234 ( .I(n2410), .Z(o_data_bus[230]) );
  BUFFD12BWP30P140 U1235 ( .I(n2413), .Z(o_data_bus[227]) );
  BUFFD12BWP30P140 U1236 ( .I(n2414), .Z(o_data_bus[226]) );
  BUFFD12BWP30P140 U1237 ( .I(n2411), .Z(o_data_bus[229]) );
  BUFFD12BWP30P140 U1238 ( .I(n2416), .Z(o_data_bus[224]) );
  BUFFD12BWP30P140 U1239 ( .I(n2415), .Z(o_data_bus[225]) );
  BUFFD12BWP30P140 U1240 ( .I(n2412), .Z(o_data_bus[228]) );
  BUFFD12BWP30P140 U1241 ( .I(n2477), .Z(o_data_bus[163]) );
  BUFFD12BWP30P140 U1242 ( .I(n2475), .Z(o_data_bus[165]) );
  BUFFD12BWP30P140 U1243 ( .I(n2474), .Z(o_data_bus[166]) );
  BUFFD12BWP30P140 U1244 ( .I(n2473), .Z(o_data_bus[167]) );
  BUFFD12BWP30P140 U1245 ( .I(n2476), .Z(o_data_bus[164]) );
  BUFFD12BWP30P140 U1246 ( .I(n2288), .Z(o_data_bus[352]) );
  BUFFD12BWP30P140 U1247 ( .I(n2287), .Z(o_data_bus[353]) );
  BUFFD12BWP30P140 U1248 ( .I(n2286), .Z(o_data_bus[354]) );
  BUFFD12BWP30P140 U1249 ( .I(n2285), .Z(o_data_bus[355]) );
  BUFFD12BWP30P140 U1250 ( .I(n2284), .Z(o_data_bus[356]) );
  BUFFD12BWP30P140 U1251 ( .I(n2283), .Z(o_data_bus[357]) );
  BUFFD12BWP30P140 U1252 ( .I(n2282), .Z(o_data_bus[358]) );
  BUFFD12BWP30P140 U1253 ( .I(n2281), .Z(o_data_bus[359]) );
  BUFFD12BWP30P140 U1254 ( .I(n2217), .Z(o_data_bus[423]) );
  BUFFD12BWP30P140 U1255 ( .I(n2218), .Z(o_data_bus[422]) );
  BUFFD12BWP30P140 U1256 ( .I(n2219), .Z(o_data_bus[421]) );
  BUFFD12BWP30P140 U1257 ( .I(n2220), .Z(o_data_bus[420]) );
  BUFFD12BWP30P140 U1258 ( .I(n2221), .Z(o_data_bus[419]) );
  BUFFD12BWP30P140 U1259 ( .I(n2222), .Z(o_data_bus[418]) );
  BUFFD12BWP30P140 U1260 ( .I(n2223), .Z(o_data_bus[417]) );
  BUFFD12BWP30P140 U1261 ( .I(n2224), .Z(o_data_bus[416]) );
  BUFFD12BWP30P140 U1262 ( .I(n2352), .Z(o_data_bus[288]) );
  BUFFD12BWP30P140 U1263 ( .I(n2351), .Z(o_data_bus[289]) );
  BUFFD12BWP30P140 U1264 ( .I(n2350), .Z(o_data_bus[290]) );
  BUFFD12BWP30P140 U1265 ( .I(n2349), .Z(o_data_bus[291]) );
  BUFFD12BWP30P140 U1266 ( .I(n2348), .Z(o_data_bus[292]) );
  BUFFD12BWP30P140 U1267 ( .I(n2347), .Z(o_data_bus[293]) );
  BUFFD12BWP30P140 U1268 ( .I(n2346), .Z(o_data_bus[294]) );
  BUFFD12BWP30P140 U1269 ( .I(n2345), .Z(o_data_bus[295]) );
  BUFFD12BWP30P140 U1270 ( .I(n2153), .Z(o_data_bus[487]) );
  BUFFD12BWP30P140 U1271 ( .I(n2154), .Z(o_data_bus[486]) );
  BUFFD12BWP30P140 U1272 ( .I(n2155), .Z(o_data_bus[485]) );
  BUFFD12BWP30P140 U1273 ( .I(n2156), .Z(o_data_bus[484]) );
  BUFFD12BWP30P140 U1274 ( .I(n2157), .Z(o_data_bus[483]) );
  BUFFD12BWP30P140 U1275 ( .I(n2158), .Z(o_data_bus[482]) );
  BUFFD12BWP30P140 U1276 ( .I(n2159), .Z(o_data_bus[481]) );
  BUFFD12BWP30P140 U1277 ( .I(n2160), .Z(o_data_bus[480]) );
  BUFFD12BWP30P140 U1278 ( .I(n2608), .Z(o_data_bus[32]) );
  BUFFD12BWP30P140 U1279 ( .I(n2607), .Z(o_data_bus[33]) );
  BUFFD12BWP30P140 U1280 ( .I(n2606), .Z(o_data_bus[34]) );
  BUFFD12BWP30P140 U1281 ( .I(n2605), .Z(o_data_bus[35]) );
  BUFFD12BWP30P140 U1282 ( .I(n2604), .Z(o_data_bus[36]) );
  BUFFD12BWP30P140 U1283 ( .I(n2603), .Z(o_data_bus[37]) );
  BUFFD12BWP30P140 U1284 ( .I(n2602), .Z(o_data_bus[38]) );
  BUFFD12BWP30P140 U1285 ( .I(n2601), .Z(o_data_bus[39]) );
  BUFFD12BWP30P140 U1286 ( .I(n2539), .Z(o_data_bus[101]) );
  BUFFD12BWP30P140 U1287 ( .I(n2538), .Z(o_data_bus[102]) );
  BUFFD12BWP30P140 U1288 ( .I(n2537), .Z(o_data_bus[103]) );
  BUFFD12BWP30P140 U1289 ( .I(n2540), .Z(o_data_bus[100]) );
  BUFFD12BWP30P140 U1290 ( .I(n2480), .Z(o_data_bus[160]) );
  BUFFD12BWP30P140 U1291 ( .I(n2479), .Z(o_data_bus[161]) );
  BUFFD12BWP30P140 U1292 ( .I(n2478), .Z(o_data_bus[162]) );
  BUFFD12BWP30P140 U1293 ( .I(n2544), .Z(o_data_bus[96]) );
  BUFFD12BWP30P140 U1294 ( .I(n2542), .Z(o_data_bus[98]) );
  BUFFD12BWP30P140 U1295 ( .I(n2541), .Z(o_data_bus[99]) );
  BUFFD12BWP30P140 U1296 ( .I(n2543), .Z(o_data_bus[97]) );
  BUFFD12BWP30P140 U1297 ( .I(n2096), .Z(o_data_bus[544]) );
  BUFFD12BWP30P140 U1298 ( .I(n2095), .Z(o_data_bus[545]) );
  BUFFD12BWP30P140 U1299 ( .I(n2094), .Z(o_data_bus[546]) );
  BUFFD12BWP30P140 U1300 ( .I(n2093), .Z(o_data_bus[547]) );
  BUFFD12BWP30P140 U1301 ( .I(n2092), .Z(o_data_bus[548]) );
  BUFFD12BWP30P140 U1302 ( .I(n2091), .Z(o_data_bus[549]) );
  BUFFD12BWP30P140 U1303 ( .I(n2090), .Z(o_data_bus[550]) );
  BUFFD12BWP30P140 U1304 ( .I(n2089), .Z(o_data_bus[551]) );
  BUFFD12BWP30P140 U1305 ( .I(n2088), .Z(o_data_bus[552]) );
  BUFFD12BWP30P140 U1306 ( .I(n2087), .Z(o_data_bus[553]) );
  BUFFD12BWP30P140 U1307 ( .I(n2086), .Z(o_data_bus[554]) );
  BUFFD12BWP30P140 U1308 ( .I(n2085), .Z(o_data_bus[555]) );
  BUFFD12BWP30P140 U1309 ( .I(n2084), .Z(o_data_bus[556]) );
  BUFFD12BWP30P140 U1310 ( .I(n2083), .Z(o_data_bus[557]) );
  BUFFD12BWP30P140 U1311 ( .I(n2082), .Z(o_data_bus[558]) );
  BUFFD12BWP30P140 U1312 ( .I(n2081), .Z(o_data_bus[559]) );
  BUFFD12BWP30P140 U1313 ( .I(n2080), .Z(o_data_bus[560]) );
  BUFFD12BWP30P140 U1314 ( .I(n2079), .Z(o_data_bus[561]) );
  BUFFD12BWP30P140 U1315 ( .I(n2078), .Z(o_data_bus[562]) );
  BUFFD12BWP30P140 U1316 ( .I(n2077), .Z(o_data_bus[563]) );
  BUFFD12BWP30P140 U1317 ( .I(n2076), .Z(o_data_bus[564]) );
  BUFFD12BWP30P140 U1318 ( .I(n2075), .Z(o_data_bus[565]) );
  BUFFD12BWP30P140 U1319 ( .I(n2074), .Z(o_data_bus[566]) );
  BUFFD12BWP30P140 U1320 ( .I(n2073), .Z(o_data_bus[567]) );
  BUFFD12BWP30P140 U1321 ( .I(n2072), .Z(o_data_bus[568]) );
  BUFFD12BWP30P140 U1322 ( .I(n2071), .Z(o_data_bus[569]) );
  BUFFD12BWP30P140 U1323 ( .I(n2070), .Z(o_data_bus[570]) );
  BUFFD12BWP30P140 U1324 ( .I(n2069), .Z(o_data_bus[571]) );
  BUFFD12BWP30P140 U1325 ( .I(n2068), .Z(o_data_bus[572]) );
  BUFFD12BWP30P140 U1326 ( .I(n2067), .Z(o_data_bus[573]) );
  BUFFD12BWP30P140 U1327 ( .I(n2066), .Z(o_data_bus[574]) );
  BUFFD12BWP30P140 U1328 ( .I(n2065), .Z(o_data_bus[575]) );
  BUFFD12BWP30P140 U1329 ( .I(n2032), .Z(o_data_bus[608]) );
  BUFFD12BWP30P140 U1330 ( .I(n2031), .Z(o_data_bus[609]) );
  BUFFD12BWP30P140 U1331 ( .I(n2030), .Z(o_data_bus[610]) );
  BUFFD12BWP30P140 U1332 ( .I(n2029), .Z(o_data_bus[611]) );
  BUFFD12BWP30P140 U1333 ( .I(n2028), .Z(o_data_bus[612]) );
  BUFFD12BWP30P140 U1334 ( .I(n2027), .Z(o_data_bus[613]) );
  BUFFD12BWP30P140 U1335 ( .I(n2026), .Z(o_data_bus[614]) );
  BUFFD12BWP30P140 U1336 ( .I(n2025), .Z(o_data_bus[615]) );
  BUFFD12BWP30P140 U1337 ( .I(n2024), .Z(o_data_bus[616]) );
  BUFFD12BWP30P140 U1338 ( .I(n2023), .Z(o_data_bus[617]) );
  BUFFD12BWP30P140 U1339 ( .I(n2022), .Z(o_data_bus[618]) );
  BUFFD12BWP30P140 U1340 ( .I(n2021), .Z(o_data_bus[619]) );
  BUFFD12BWP30P140 U1341 ( .I(n2020), .Z(o_data_bus[620]) );
  BUFFD12BWP30P140 U1342 ( .I(n2019), .Z(o_data_bus[621]) );
  BUFFD12BWP30P140 U1343 ( .I(n2018), .Z(o_data_bus[622]) );
  BUFFD12BWP30P140 U1344 ( .I(n2017), .Z(o_data_bus[623]) );
  BUFFD12BWP30P140 U1345 ( .I(n2016), .Z(o_data_bus[624]) );
  BUFFD12BWP30P140 U1346 ( .I(n2015), .Z(o_data_bus[625]) );
  BUFFD12BWP30P140 U1347 ( .I(n2014), .Z(o_data_bus[626]) );
  BUFFD12BWP30P140 U1348 ( .I(n2013), .Z(o_data_bus[627]) );
  BUFFD12BWP30P140 U1349 ( .I(n2012), .Z(o_data_bus[628]) );
  BUFFD12BWP30P140 U1350 ( .I(n2011), .Z(o_data_bus[629]) );
  BUFFD12BWP30P140 U1351 ( .I(n2010), .Z(o_data_bus[630]) );
  BUFFD12BWP30P140 U1352 ( .I(n2009), .Z(o_data_bus[631]) );
  BUFFD12BWP30P140 U1353 ( .I(n2008), .Z(o_data_bus[632]) );
  BUFFD12BWP30P140 U1354 ( .I(n2007), .Z(o_data_bus[633]) );
  BUFFD12BWP30P140 U1355 ( .I(n2006), .Z(o_data_bus[634]) );
  BUFFD12BWP30P140 U1356 ( .I(n2005), .Z(o_data_bus[635]) );
  BUFFD12BWP30P140 U1357 ( .I(n2004), .Z(o_data_bus[636]) );
  BUFFD12BWP30P140 U1358 ( .I(n2003), .Z(o_data_bus[637]) );
  BUFFD12BWP30P140 U1359 ( .I(n2002), .Z(o_data_bus[638]) );
  BUFFD12BWP30P140 U1360 ( .I(n2001), .Z(o_data_bus[639]) );
  BUFFD12BWP30P140 U1361 ( .I(n1968), .Z(o_data_bus[672]) );
  BUFFD12BWP30P140 U1362 ( .I(n1967), .Z(o_data_bus[673]) );
  BUFFD12BWP30P140 U1363 ( .I(n1966), .Z(o_data_bus[674]) );
  BUFFD12BWP30P140 U1364 ( .I(n1965), .Z(o_data_bus[675]) );
  BUFFD12BWP30P140 U1365 ( .I(n1964), .Z(o_data_bus[676]) );
  BUFFD12BWP30P140 U1366 ( .I(n1963), .Z(o_data_bus[677]) );
  BUFFD12BWP30P140 U1367 ( .I(n1962), .Z(o_data_bus[678]) );
  BUFFD12BWP30P140 U1368 ( .I(n1961), .Z(o_data_bus[679]) );
  BUFFD12BWP30P140 U1369 ( .I(n1960), .Z(o_data_bus[680]) );
  BUFFD12BWP30P140 U1370 ( .I(n1959), .Z(o_data_bus[681]) );
  BUFFD12BWP30P140 U1371 ( .I(n1958), .Z(o_data_bus[682]) );
  BUFFD12BWP30P140 U1372 ( .I(n1957), .Z(o_data_bus[683]) );
  BUFFD12BWP30P140 U1373 ( .I(n1956), .Z(o_data_bus[684]) );
  BUFFD12BWP30P140 U1374 ( .I(n1955), .Z(o_data_bus[685]) );
  BUFFD12BWP30P140 U1375 ( .I(n1954), .Z(o_data_bus[686]) );
  BUFFD12BWP30P140 U1376 ( .I(n1953), .Z(o_data_bus[687]) );
  BUFFD12BWP30P140 U1377 ( .I(n1952), .Z(o_data_bus[688]) );
  BUFFD12BWP30P140 U1378 ( .I(n1951), .Z(o_data_bus[689]) );
  BUFFD12BWP30P140 U1379 ( .I(n1950), .Z(o_data_bus[690]) );
  BUFFD12BWP30P140 U1380 ( .I(n1949), .Z(o_data_bus[691]) );
  BUFFD12BWP30P140 U1381 ( .I(n1948), .Z(o_data_bus[692]) );
  BUFFD12BWP30P140 U1382 ( .I(n1947), .Z(o_data_bus[693]) );
  BUFFD12BWP30P140 U1383 ( .I(n1946), .Z(o_data_bus[694]) );
  BUFFD12BWP30P140 U1384 ( .I(n1945), .Z(o_data_bus[695]) );
  BUFFD12BWP30P140 U1385 ( .I(n1944), .Z(o_data_bus[696]) );
  BUFFD12BWP30P140 U1386 ( .I(n1943), .Z(o_data_bus[697]) );
  BUFFD12BWP30P140 U1387 ( .I(n1942), .Z(o_data_bus[698]) );
  BUFFD12BWP30P140 U1388 ( .I(n1941), .Z(o_data_bus[699]) );
  BUFFD12BWP30P140 U1389 ( .I(n1940), .Z(o_data_bus[700]) );
  BUFFD12BWP30P140 U1390 ( .I(n1939), .Z(o_data_bus[701]) );
  BUFFD12BWP30P140 U1391 ( .I(n1938), .Z(o_data_bus[702]) );
  BUFFD12BWP30P140 U1392 ( .I(n1937), .Z(o_data_bus[703]) );
  BUFFD12BWP30P140 U1393 ( .I(n1904), .Z(o_data_bus[736]) );
  BUFFD12BWP30P140 U1394 ( .I(n1903), .Z(o_data_bus[737]) );
  BUFFD12BWP30P140 U1395 ( .I(n1902), .Z(o_data_bus[738]) );
  BUFFD12BWP30P140 U1396 ( .I(n1901), .Z(o_data_bus[739]) );
  BUFFD12BWP30P140 U1397 ( .I(n1900), .Z(o_data_bus[740]) );
  BUFFD12BWP30P140 U1398 ( .I(n1899), .Z(o_data_bus[741]) );
  BUFFD12BWP30P140 U1399 ( .I(n1898), .Z(o_data_bus[742]) );
  BUFFD12BWP30P140 U1400 ( .I(n1897), .Z(o_data_bus[743]) );
  BUFFD12BWP30P140 U1401 ( .I(n1896), .Z(o_data_bus[744]) );
  BUFFD12BWP30P140 U1402 ( .I(n1895), .Z(o_data_bus[745]) );
  BUFFD12BWP30P140 U1403 ( .I(n1894), .Z(o_data_bus[746]) );
  BUFFD12BWP30P140 U1404 ( .I(n1893), .Z(o_data_bus[747]) );
  BUFFD12BWP30P140 U1405 ( .I(n1892), .Z(o_data_bus[748]) );
  BUFFD12BWP30P140 U1406 ( .I(n1891), .Z(o_data_bus[749]) );
  BUFFD12BWP30P140 U1407 ( .I(n1890), .Z(o_data_bus[750]) );
  BUFFD12BWP30P140 U1408 ( .I(n1889), .Z(o_data_bus[751]) );
  BUFFD12BWP30P140 U1409 ( .I(n1888), .Z(o_data_bus[752]) );
  BUFFD12BWP30P140 U1410 ( .I(n1887), .Z(o_data_bus[753]) );
  BUFFD12BWP30P140 U1411 ( .I(n1886), .Z(o_data_bus[754]) );
  BUFFD12BWP30P140 U1412 ( .I(n1885), .Z(o_data_bus[755]) );
  BUFFD12BWP30P140 U1413 ( .I(n1884), .Z(o_data_bus[756]) );
  BUFFD12BWP30P140 U1414 ( .I(n1883), .Z(o_data_bus[757]) );
  BUFFD12BWP30P140 U1415 ( .I(n1882), .Z(o_data_bus[758]) );
  BUFFD12BWP30P140 U1416 ( .I(n1881), .Z(o_data_bus[759]) );
  BUFFD12BWP30P140 U1417 ( .I(n1880), .Z(o_data_bus[760]) );
  BUFFD12BWP30P140 U1418 ( .I(n1879), .Z(o_data_bus[761]) );
  BUFFD12BWP30P140 U1419 ( .I(n1878), .Z(o_data_bus[762]) );
  BUFFD12BWP30P140 U1420 ( .I(n1877), .Z(o_data_bus[763]) );
  BUFFD12BWP30P140 U1421 ( .I(n1876), .Z(o_data_bus[764]) );
  BUFFD12BWP30P140 U1422 ( .I(n1875), .Z(o_data_bus[765]) );
  BUFFD12BWP30P140 U1423 ( .I(n1874), .Z(o_data_bus[766]) );
  BUFFD12BWP30P140 U1424 ( .I(n1873), .Z(o_data_bus[767]) );
  BUFFD12BWP30P140 U1425 ( .I(n1840), .Z(o_data_bus[800]) );
  BUFFD12BWP30P140 U1426 ( .I(n1839), .Z(o_data_bus[801]) );
  BUFFD12BWP30P140 U1427 ( .I(n1838), .Z(o_data_bus[802]) );
  BUFFD12BWP30P140 U1428 ( .I(n1837), .Z(o_data_bus[803]) );
  BUFFD12BWP30P140 U1429 ( .I(n1836), .Z(o_data_bus[804]) );
  BUFFD12BWP30P140 U1430 ( .I(n1835), .Z(o_data_bus[805]) );
  BUFFD12BWP30P140 U1431 ( .I(n1834), .Z(o_data_bus[806]) );
  BUFFD12BWP30P140 U1432 ( .I(n1833), .Z(o_data_bus[807]) );
  BUFFD12BWP30P140 U1433 ( .I(n1832), .Z(o_data_bus[808]) );
  BUFFD12BWP30P140 U1434 ( .I(n1831), .Z(o_data_bus[809]) );
  BUFFD12BWP30P140 U1435 ( .I(n1830), .Z(o_data_bus[810]) );
  BUFFD12BWP30P140 U1436 ( .I(n1829), .Z(o_data_bus[811]) );
  BUFFD12BWP30P140 U1437 ( .I(n1828), .Z(o_data_bus[812]) );
  BUFFD12BWP30P140 U1438 ( .I(n1827), .Z(o_data_bus[813]) );
  BUFFD12BWP30P140 U1439 ( .I(n1826), .Z(o_data_bus[814]) );
  BUFFD12BWP30P140 U1440 ( .I(n1825), .Z(o_data_bus[815]) );
  BUFFD12BWP30P140 U1441 ( .I(n1824), .Z(o_data_bus[816]) );
  BUFFD12BWP30P140 U1442 ( .I(n1823), .Z(o_data_bus[817]) );
  BUFFD12BWP30P140 U1443 ( .I(n1822), .Z(o_data_bus[818]) );
  BUFFD12BWP30P140 U1444 ( .I(n1821), .Z(o_data_bus[819]) );
  BUFFD12BWP30P140 U1445 ( .I(n1820), .Z(o_data_bus[820]) );
  BUFFD12BWP30P140 U1446 ( .I(n1819), .Z(o_data_bus[821]) );
  BUFFD12BWP30P140 U1447 ( .I(n1818), .Z(o_data_bus[822]) );
  BUFFD12BWP30P140 U1448 ( .I(n1817), .Z(o_data_bus[823]) );
  BUFFD12BWP30P140 U1449 ( .I(n1816), .Z(o_data_bus[824]) );
  BUFFD12BWP30P140 U1450 ( .I(n1815), .Z(o_data_bus[825]) );
  BUFFD12BWP30P140 U1451 ( .I(n1814), .Z(o_data_bus[826]) );
  BUFFD12BWP30P140 U1452 ( .I(n1813), .Z(o_data_bus[827]) );
  BUFFD12BWP30P140 U1453 ( .I(n1812), .Z(o_data_bus[828]) );
  BUFFD12BWP30P140 U1454 ( .I(n1811), .Z(o_data_bus[829]) );
  BUFFD12BWP30P140 U1455 ( .I(n1810), .Z(o_data_bus[830]) );
  BUFFD12BWP30P140 U1456 ( .I(n1809), .Z(o_data_bus[831]) );
  BUFFD12BWP30P140 U1457 ( .I(n1776), .Z(o_data_bus[864]) );
  BUFFD12BWP30P140 U1458 ( .I(n1775), .Z(o_data_bus[865]) );
  BUFFD12BWP30P140 U1459 ( .I(n1774), .Z(o_data_bus[866]) );
  BUFFD12BWP30P140 U1460 ( .I(n1773), .Z(o_data_bus[867]) );
  BUFFD12BWP30P140 U1461 ( .I(n1772), .Z(o_data_bus[868]) );
  BUFFD12BWP30P140 U1462 ( .I(n1771), .Z(o_data_bus[869]) );
  BUFFD12BWP30P140 U1463 ( .I(n1770), .Z(o_data_bus[870]) );
  BUFFD12BWP30P140 U1464 ( .I(n1769), .Z(o_data_bus[871]) );
  BUFFD12BWP30P140 U1465 ( .I(n1768), .Z(o_data_bus[872]) );
  BUFFD12BWP30P140 U1466 ( .I(n1767), .Z(o_data_bus[873]) );
  BUFFD12BWP30P140 U1467 ( .I(n1766), .Z(o_data_bus[874]) );
  BUFFD12BWP30P140 U1468 ( .I(n1765), .Z(o_data_bus[875]) );
  BUFFD12BWP30P140 U1469 ( .I(n1764), .Z(o_data_bus[876]) );
  BUFFD12BWP30P140 U1470 ( .I(n1763), .Z(o_data_bus[877]) );
  BUFFD12BWP30P140 U1471 ( .I(n1762), .Z(o_data_bus[878]) );
  BUFFD12BWP30P140 U1472 ( .I(n1761), .Z(o_data_bus[879]) );
  BUFFD12BWP30P140 U1473 ( .I(n1760), .Z(o_data_bus[880]) );
  BUFFD12BWP30P140 U1474 ( .I(n1759), .Z(o_data_bus[881]) );
  BUFFD12BWP30P140 U1475 ( .I(n1758), .Z(o_data_bus[882]) );
  BUFFD12BWP30P140 U1476 ( .I(n1757), .Z(o_data_bus[883]) );
  BUFFD12BWP30P140 U1477 ( .I(n1756), .Z(o_data_bus[884]) );
  BUFFD12BWP30P140 U1478 ( .I(n1755), .Z(o_data_bus[885]) );
  BUFFD12BWP30P140 U1479 ( .I(n1754), .Z(o_data_bus[886]) );
  BUFFD12BWP30P140 U1480 ( .I(n1753), .Z(o_data_bus[887]) );
  BUFFD12BWP30P140 U1481 ( .I(n1752), .Z(o_data_bus[888]) );
  BUFFD12BWP30P140 U1482 ( .I(n1751), .Z(o_data_bus[889]) );
  BUFFD12BWP30P140 U1483 ( .I(n1750), .Z(o_data_bus[890]) );
  BUFFD12BWP30P140 U1484 ( .I(n1749), .Z(o_data_bus[891]) );
  BUFFD12BWP30P140 U1485 ( .I(n1748), .Z(o_data_bus[892]) );
  BUFFD12BWP30P140 U1486 ( .I(n1747), .Z(o_data_bus[893]) );
  BUFFD12BWP30P140 U1487 ( .I(n1746), .Z(o_data_bus[894]) );
  BUFFD12BWP30P140 U1488 ( .I(n1745), .Z(o_data_bus[895]) );
  BUFFD12BWP30P140 U1489 ( .I(n1712), .Z(o_data_bus[928]) );
  BUFFD12BWP30P140 U1490 ( .I(n1711), .Z(o_data_bus[929]) );
  BUFFD12BWP30P140 U1491 ( .I(n1710), .Z(o_data_bus[930]) );
  BUFFD12BWP30P140 U1492 ( .I(n1709), .Z(o_data_bus[931]) );
  BUFFD12BWP30P140 U1493 ( .I(n1708), .Z(o_data_bus[932]) );
  BUFFD12BWP30P140 U1494 ( .I(n1707), .Z(o_data_bus[933]) );
  BUFFD12BWP30P140 U1495 ( .I(n1706), .Z(o_data_bus[934]) );
  BUFFD12BWP30P140 U1496 ( .I(n1705), .Z(o_data_bus[935]) );
  BUFFD12BWP30P140 U1497 ( .I(n1704), .Z(o_data_bus[936]) );
  BUFFD12BWP30P140 U1498 ( .I(n1703), .Z(o_data_bus[937]) );
  BUFFD12BWP30P140 U1499 ( .I(n1702), .Z(o_data_bus[938]) );
  BUFFD12BWP30P140 U1500 ( .I(n1701), .Z(o_data_bus[939]) );
  BUFFD12BWP30P140 U1501 ( .I(n1700), .Z(o_data_bus[940]) );
  BUFFD12BWP30P140 U1502 ( .I(n1699), .Z(o_data_bus[941]) );
  BUFFD12BWP30P140 U1503 ( .I(n1698), .Z(o_data_bus[942]) );
  BUFFD12BWP30P140 U1504 ( .I(n1697), .Z(o_data_bus[943]) );
  BUFFD12BWP30P140 U1505 ( .I(n1696), .Z(o_data_bus[944]) );
  BUFFD12BWP30P140 U1506 ( .I(n1695), .Z(o_data_bus[945]) );
  BUFFD12BWP30P140 U1507 ( .I(n1694), .Z(o_data_bus[946]) );
  BUFFD12BWP30P140 U1508 ( .I(n1693), .Z(o_data_bus[947]) );
  BUFFD12BWP30P140 U1509 ( .I(n1692), .Z(o_data_bus[948]) );
  BUFFD12BWP30P140 U1510 ( .I(n1691), .Z(o_data_bus[949]) );
  BUFFD12BWP30P140 U1511 ( .I(n1690), .Z(o_data_bus[950]) );
  BUFFD12BWP30P140 U1512 ( .I(n1689), .Z(o_data_bus[951]) );
  BUFFD12BWP30P140 U1513 ( .I(n1688), .Z(o_data_bus[952]) );
  BUFFD12BWP30P140 U1514 ( .I(n1687), .Z(o_data_bus[953]) );
  BUFFD12BWP30P140 U1515 ( .I(n1686), .Z(o_data_bus[954]) );
  BUFFD12BWP30P140 U1516 ( .I(n1685), .Z(o_data_bus[955]) );
  BUFFD12BWP30P140 U1517 ( .I(n1684), .Z(o_data_bus[956]) );
  BUFFD12BWP30P140 U1518 ( .I(n1683), .Z(o_data_bus[957]) );
  BUFFD12BWP30P140 U1519 ( .I(n1682), .Z(o_data_bus[958]) );
  BUFFD12BWP30P140 U1520 ( .I(n1681), .Z(o_data_bus[959]) );
  BUFFD12BWP30P140 U1521 ( .I(n1650), .Z(o_data_bus[990]) );
  BUFFD12BWP30P140 U1522 ( .I(n1649), .Z(o_data_bus[991]) );
  BUFFD12BWP30P140 U1523 ( .I(n1648), .Z(o_data_bus[992]) );
  BUFFD12BWP30P140 U1524 ( .I(n1647), .Z(o_data_bus[993]) );
  BUFFD12BWP30P140 U1525 ( .I(n1646), .Z(o_data_bus[994]) );
  BUFFD12BWP30P140 U1526 ( .I(n1645), .Z(o_data_bus[995]) );
  BUFFD12BWP30P140 U1527 ( .I(n1644), .Z(o_data_bus[996]) );
  BUFFD12BWP30P140 U1528 ( .I(n1643), .Z(o_data_bus[997]) );
  BUFFD12BWP30P140 U1529 ( .I(n1642), .Z(o_data_bus[998]) );
  BUFFD12BWP30P140 U1530 ( .I(n1641), .Z(o_data_bus[999]) );
  BUFFD12BWP30P140 U1531 ( .I(n1640), .Z(o_data_bus[1000]) );
  BUFFD12BWP30P140 U1532 ( .I(n1639), .Z(o_data_bus[1001]) );
  BUFFD12BWP30P140 U1533 ( .I(n1638), .Z(o_data_bus[1002]) );
  BUFFD12BWP30P140 U1534 ( .I(n1637), .Z(o_data_bus[1003]) );
  BUFFD12BWP30P140 U1535 ( .I(n1636), .Z(o_data_bus[1004]) );
  BUFFD12BWP30P140 U1536 ( .I(n1635), .Z(o_data_bus[1005]) );
  BUFFD12BWP30P140 U1537 ( .I(n1634), .Z(o_data_bus[1006]) );
  BUFFD12BWP30P140 U1538 ( .I(n1633), .Z(o_data_bus[1007]) );
  BUFFD12BWP30P140 U1539 ( .I(n1632), .Z(o_data_bus[1008]) );
  BUFFD12BWP30P140 U1540 ( .I(n1631), .Z(o_data_bus[1009]) );
  BUFFD12BWP30P140 U1541 ( .I(n1630), .Z(o_data_bus[1010]) );
  BUFFD12BWP30P140 U1542 ( .I(n1629), .Z(o_data_bus[1011]) );
  BUFFD12BWP30P140 U1543 ( .I(n1628), .Z(o_data_bus[1012]) );
  BUFFD12BWP30P140 U1544 ( .I(n1627), .Z(o_data_bus[1013]) );
  BUFFD12BWP30P140 U1545 ( .I(n1626), .Z(o_data_bus[1014]) );
  BUFFD12BWP30P140 U1546 ( .I(n1625), .Z(o_data_bus[1015]) );
  BUFFD12BWP30P140 U1547 ( .I(n1624), .Z(o_data_bus[1016]) );
  BUFFD12BWP30P140 U1548 ( .I(n1623), .Z(o_data_bus[1017]) );
  BUFFD12BWP30P140 U1549 ( .I(n1622), .Z(o_data_bus[1018]) );
  BUFFD12BWP30P140 U1550 ( .I(n1621), .Z(o_data_bus[1019]) );
  BUFFD12BWP30P140 U1551 ( .I(n1620), .Z(o_data_bus[1020]) );
  BUFFD12BWP30P140 U1552 ( .I(n1619), .Z(o_data_bus[1021]) );
  BUFFD12BWP30P140 U1553 ( .I(n1618), .Z(o_data_bus[1022]) );
  BUFFD12BWP30P140 U1554 ( .I(n1617), .Z(o_data_bus[1023]) );
  BUFFD12BWP30P140 U1555 ( .I(n1616), .Z(o_valid[0]) );
  BUFFD12BWP30P140 U1556 ( .I(n1614), .Z(o_valid[2]) );
  BUFFD12BWP30P140 U1557 ( .I(n1612), .Z(o_valid[4]) );
  BUFFD12BWP30P140 U1558 ( .I(n1610), .Z(o_valid[6]) );
  BUFFD12BWP30P140 U1559 ( .I(n1608), .Z(o_valid[8]) );
  BUFFD12BWP30P140 U1560 ( .I(n1606), .Z(o_valid[10]) );
  BUFFD12BWP30P140 U1561 ( .I(n1604), .Z(o_valid[12]) );
  BUFFD12BWP30P140 U1562 ( .I(n1602), .Z(o_valid[14]) );
  BUFFD12BWP30P140 U1563 ( .I(n1600), .Z(o_valid[16]) );
  BUFFD12BWP30P140 U1564 ( .I(n1598), .Z(o_valid[18]) );
  BUFFD12BWP30P140 U1565 ( .I(n1596), .Z(o_valid[20]) );
  BUFFD12BWP30P140 U1566 ( .I(n1594), .Z(o_valid[22]) );
  BUFFD12BWP30P140 U1567 ( .I(n1592), .Z(o_valid[24]) );
  BUFFD12BWP30P140 U1568 ( .I(n1590), .Z(o_valid[26]) );
  BUFFD12BWP30P140 U1569 ( .I(n1588), .Z(o_valid[28]) );
  BUFFD12BWP30P140 U1570 ( .I(n1586), .Z(o_valid[30]) );
  INVD2BWP30P140 U1571 ( .I(n1609), .ZN(n1547) );
  INVD2BWP30P140 U1572 ( .I(n1615), .ZN(n1538) );
  INVD2BWP30P140 U1573 ( .I(n1605), .ZN(n1553) );
  INVD2BWP30P140 U1574 ( .I(n1607), .ZN(n1550) );
  INVD2BWP30P140 U1575 ( .I(n1587), .ZN(n1580) );
  INVD2BWP30P140 U1576 ( .I(n1589), .ZN(n1577) );
  INVD2BWP30P140 U1577 ( .I(n1591), .ZN(n1574) );
  INVD2BWP30P140 U1578 ( .I(n1611), .ZN(n1544) );
  INVD2BWP30P140 U1579 ( .I(n1613), .ZN(n1541) );
  INVD2BWP30P140 U1580 ( .I(n1595), .ZN(n1568) );
  INVD2BWP30P140 U1581 ( .I(n1597), .ZN(n1565) );
  INVD2BWP30P140 U1582 ( .I(n1599), .ZN(n1562) );
  INVD2BWP30P140 U1583 ( .I(n1601), .ZN(n1559) );
  INVD2BWP30P140 U1584 ( .I(n1603), .ZN(n1556) );
  INVD2BWP30P140 U1585 ( .I(n1593), .ZN(n1571) );
  INVD2BWP30P140 U1586 ( .I(n1585), .ZN(n1583) );
endmodule

