
module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_0 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  INVD6BWP30P140LVT U3 ( .I(n2), .ZN(n7) );
  OR3D2BWP30P140LVT U4 ( .A1(n3), .A2(i_cmd[0]), .A3(rst), .Z(n2) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n4) );
  BUFFD4BWP30P140LVT U6 ( .I(n5), .Z(n1) );
  BUFFD4BWP30P140LVT U7 ( .I(n5), .Z(n6) );
  NR2OPTPAD2BWP30P140LVT U8 ( .A1(n4), .A2(rst), .ZN(n5) );
  ND2OPTIBD1BWP30P140LVT U9 ( .A1(i_en), .A2(i_valid[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U10 ( .A1(n7), .A2(i_data_bus[0]), .B1(n6), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U11 ( .A1(n7), .A2(i_data_bus[1]), .B1(n6), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U12 ( .A1(n7), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U13 ( .A1(n7), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U14 ( .A1(n7), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U15 ( .A1(n7), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U16 ( .A1(n7), .A2(i_data_bus[6]), .B1(n6), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U17 ( .A1(n7), .A2(i_data_bus[7]), .B1(n6), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U18 ( .A1(n7), .A2(i_data_bus[8]), .B1(n6), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U19 ( .A1(n7), .A2(i_data_bus[9]), .B1(n6), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U20 ( .A1(n7), .A2(i_data_bus[10]), .B1(n6), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U21 ( .A1(n7), .A2(i_data_bus[11]), .B1(n6), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U22 ( .A1(n7), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U23 ( .A1(n7), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U24 ( .A1(n7), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U25 ( .A1(n7), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U26 ( .A1(n7), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U27 ( .A1(n7), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U28 ( .A1(n7), .A2(i_data_bus[18]), .B1(n6), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U29 ( .A1(n7), .A2(i_data_bus[19]), .B1(n6), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U30 ( .A1(n7), .A2(i_data_bus[20]), .B1(n6), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U31 ( .A1(n7), .A2(i_data_bus[21]), .B1(n6), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U32 ( .A1(n7), .A2(i_data_bus[22]), .B1(n6), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U33 ( .A1(n7), .A2(i_data_bus[23]), .B1(n6), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U34 ( .A1(n7), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U35 ( .A1(n7), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U36 ( .A1(n7), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U37 ( .A1(n7), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U38 ( .A1(n7), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U39 ( .A1(n7), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U40 ( .A1(n7), .A2(i_data_bus[30]), .B1(n6), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U41 ( .A1(n7), .A2(i_data_bus[31]), .B1(n6), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U42 ( .A1(n7), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_0 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_0 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_283 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND3D1BWP30P140LVT U3 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  INVD8BWP30P140LVT U4 ( .I(n3), .ZN(n4) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  OR2D4BWP30P140LVT U7 ( .A1(n2), .A2(rst), .Z(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_283 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_283 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_284 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2OPTIBD2BWP30P140LVT U3 ( .A1(i_cmd[0]), .A2(n4), .ZN(n5) );
  INR2D1BWP30P140LVT U4 ( .A1(i_en), .B1(n3), .ZN(n4) );
  NR2D2BWP30P140LVT U5 ( .A1(n5), .A2(rst), .ZN(n1) );
  ND2D1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR2D2BWP30P140LVT U7 ( .A1(n5), .A2(rst), .ZN(n6) );
  NR3OPTPAD2BWP30P140LVT U8 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n7) );
  INVD1BWP30P140LVT U9 ( .I(i_valid[1]), .ZN(n3) );
  AO22D1BWP30P140LVT U10 ( .A1(n7), .A2(i_data_bus[0]), .B1(n6), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U11 ( .A1(n7), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U12 ( .A1(n7), .A2(i_data_bus[2]), .B1(n6), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U13 ( .A1(n7), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U14 ( .A1(n7), .A2(i_data_bus[4]), .B1(n6), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U15 ( .A1(n7), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U16 ( .A1(n7), .A2(i_data_bus[6]), .B1(n6), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U17 ( .A1(n7), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U18 ( .A1(n7), .A2(i_data_bus[8]), .B1(n6), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U19 ( .A1(n7), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U20 ( .A1(n7), .A2(i_data_bus[10]), .B1(n6), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U21 ( .A1(n7), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U22 ( .A1(n7), .A2(i_data_bus[12]), .B1(n6), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U23 ( .A1(n7), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U24 ( .A1(n7), .A2(i_data_bus[14]), .B1(n6), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U25 ( .A1(n7), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U26 ( .A1(n7), .A2(i_data_bus[16]), .B1(n6), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U27 ( .A1(n7), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U28 ( .A1(n7), .A2(i_data_bus[18]), .B1(n6), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U29 ( .A1(n7), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U30 ( .A1(n7), .A2(i_data_bus[20]), .B1(n6), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U31 ( .A1(n7), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U32 ( .A1(n7), .A2(i_data_bus[22]), .B1(n6), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U33 ( .A1(n7), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U34 ( .A1(n7), .A2(i_data_bus[24]), .B1(n6), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U35 ( .A1(n7), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U36 ( .A1(n7), .A2(i_data_bus[26]), .B1(n6), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U37 ( .A1(n7), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U38 ( .A1(n7), .A2(i_data_bus[28]), .B1(n6), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U39 ( .A1(n7), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U40 ( .A1(n7), .A2(i_data_bus[30]), .B1(n6), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U41 ( .A1(n7), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U42 ( .A1(n7), .A2(n6), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_284 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_284 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_285 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D2BWP30P140LVT U3 ( .A1(i_cmd[0]), .A2(n3), .ZN(N91) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U36 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  IND2D1BWP30P140LVT U37 ( .A1(n2), .B1(n1), .ZN(n3) );
  INVD1BWP30P140LVT U38 ( .I(rst), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_285 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_285 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_286 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  INVD6BWP30P140LVT U3 ( .I(n3), .ZN(n4) );
  ND3D1BWP30P140LVT U4 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  OR2D4BWP30P140LVT U7 ( .A1(n2), .A2(rst), .Z(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_286 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_286 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_287 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  INR2D4BWP30P140LVT U3 ( .A1(n1), .B1(rst), .ZN(n38) );
  NR3D1P5BWP30P140LVT U4 ( .A1(n4), .A2(i_cmd[0]), .A3(rst), .ZN(n39) );
  INVD1BWP30P140LVT U5 ( .I(i_en), .ZN(n2) );
  INVD3BWP30P140LVT U6 ( .I(n39), .ZN(n37) );
  INVD1BWP30P140LVT U7 ( .I(i_cmd[0]), .ZN(n3) );
  INR3D1BWP30P140LVT U8 ( .A1(i_valid[1]), .B1(n2), .B2(n3), .ZN(n1) );
  ND2OPTIBD1BWP30P140LVT U9 ( .A1(i_en), .A2(i_valid[0]), .ZN(n4) );
  INVD1BWP30P140LVT U10 ( .I(i_data_bus[25]), .ZN(n5) );
  MOAI22D1BWP30P140LVT U11 ( .A1(n37), .A2(n5), .B1(n38), .B2(i_data_bus[57]), 
        .ZN(N117) );
  INVD1BWP30P140LVT U12 ( .I(i_data_bus[9]), .ZN(n6) );
  MOAI22D1BWP30P140LVT U13 ( .A1(n37), .A2(n6), .B1(n38), .B2(i_data_bus[41]), 
        .ZN(N101) );
  INVD1BWP30P140LVT U14 ( .I(i_data_bus[7]), .ZN(n7) );
  MOAI22D1BWP30P140LVT U15 ( .A1(n37), .A2(n7), .B1(n38), .B2(i_data_bus[39]), 
        .ZN(N99) );
  INVD1BWP30P140LVT U16 ( .I(i_data_bus[17]), .ZN(n8) );
  MOAI22D1BWP30P140LVT U17 ( .A1(n37), .A2(n8), .B1(n38), .B2(i_data_bus[49]), 
        .ZN(N109) );
  INVD1BWP30P140LVT U18 ( .I(i_data_bus[3]), .ZN(n9) );
  MOAI22D1BWP30P140LVT U19 ( .A1(n37), .A2(n9), .B1(n38), .B2(i_data_bus[35]), 
        .ZN(N95) );
  INVD1BWP30P140LVT U20 ( .I(i_data_bus[19]), .ZN(n10) );
  MOAI22D1BWP30P140LVT U21 ( .A1(n37), .A2(n10), .B1(n38), .B2(i_data_bus[51]), 
        .ZN(N111) );
  INVD1BWP30P140LVT U22 ( .I(i_data_bus[31]), .ZN(n11) );
  MOAI22D1BWP30P140LVT U23 ( .A1(n37), .A2(n11), .B1(n38), .B2(i_data_bus[63]), 
        .ZN(N123) );
  INVD1BWP30P140LVT U24 ( .I(i_data_bus[5]), .ZN(n12) );
  MOAI22D1BWP30P140LVT U25 ( .A1(n37), .A2(n12), .B1(n38), .B2(i_data_bus[37]), 
        .ZN(N97) );
  INVD1BWP30P140LVT U26 ( .I(i_data_bus[27]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U27 ( .A1(n37), .A2(n13), .B1(n38), .B2(i_data_bus[59]), 
        .ZN(N119) );
  INVD1BWP30P140LVT U28 ( .I(i_data_bus[13]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U29 ( .A1(n37), .A2(n14), .B1(n38), .B2(i_data_bus[45]), 
        .ZN(N105) );
  INVD1BWP30P140LVT U30 ( .I(i_data_bus[1]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U31 ( .A1(n37), .A2(n15), .B1(n38), .B2(i_data_bus[33]), 
        .ZN(N93) );
  INVD1BWP30P140LVT U32 ( .I(i_data_bus[15]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U33 ( .A1(n37), .A2(n16), .B1(n38), .B2(i_data_bus[47]), 
        .ZN(N107) );
  INVD1BWP30P140LVT U34 ( .I(i_data_bus[11]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U35 ( .A1(n37), .A2(n17), .B1(n38), .B2(i_data_bus[43]), 
        .ZN(N103) );
  INVD1BWP30P140LVT U36 ( .I(i_data_bus[29]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U37 ( .A1(n37), .A2(n18), .B1(n38), .B2(i_data_bus[61]), 
        .ZN(N121) );
  INVD1BWP30P140LVT U38 ( .I(i_data_bus[23]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U39 ( .A1(n37), .A2(n19), .B1(n38), .B2(i_data_bus[55]), 
        .ZN(N115) );
  INVD1BWP30P140LVT U40 ( .I(i_data_bus[21]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U41 ( .A1(n37), .A2(n20), .B1(n38), .B2(i_data_bus[53]), 
        .ZN(N113) );
  INVD1BWP30P140LVT U42 ( .I(i_data_bus[20]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U43 ( .A1(n37), .A2(n21), .B1(n38), .B2(i_data_bus[52]), 
        .ZN(N112) );
  INVD1BWP30P140LVT U44 ( .I(i_data_bus[28]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U45 ( .A1(n37), .A2(n22), .B1(n38), .B2(i_data_bus[60]), 
        .ZN(N120) );
  INVD1BWP30P140LVT U46 ( .I(i_data_bus[24]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U47 ( .A1(n37), .A2(n23), .B1(n38), .B2(i_data_bus[56]), 
        .ZN(N116) );
  INVD1BWP30P140LVT U48 ( .I(i_data_bus[18]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U49 ( .A1(n37), .A2(n24), .B1(n38), .B2(i_data_bus[50]), 
        .ZN(N110) );
  INVD1BWP30P140LVT U50 ( .I(i_data_bus[10]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U51 ( .A1(n37), .A2(n25), .B1(n38), .B2(i_data_bus[42]), 
        .ZN(N102) );
  INVD1BWP30P140LVT U52 ( .I(i_data_bus[0]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U53 ( .A1(n37), .A2(n26), .B1(n38), .B2(i_data_bus[32]), 
        .ZN(N92) );
  INVD1BWP30P140LVT U54 ( .I(i_data_bus[8]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U55 ( .A1(n37), .A2(n27), .B1(n38), .B2(i_data_bus[40]), 
        .ZN(N100) );
  INVD1BWP30P140LVT U56 ( .I(i_data_bus[6]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U57 ( .A1(n37), .A2(n28), .B1(n38), .B2(i_data_bus[38]), 
        .ZN(N98) );
  INVD1BWP30P140LVT U58 ( .I(i_data_bus[14]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U59 ( .A1(n37), .A2(n29), .B1(n38), .B2(i_data_bus[46]), 
        .ZN(N106) );
  INVD1BWP30P140LVT U60 ( .I(i_data_bus[22]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U61 ( .A1(n37), .A2(n30), .B1(n38), .B2(i_data_bus[54]), 
        .ZN(N114) );
  INVD1BWP30P140LVT U62 ( .I(i_data_bus[30]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U63 ( .A1(n37), .A2(n31), .B1(n38), .B2(i_data_bus[62]), 
        .ZN(N122) );
  INVD1BWP30P140LVT U64 ( .I(i_data_bus[16]), .ZN(n32) );
  MOAI22D1BWP30P140LVT U65 ( .A1(n37), .A2(n32), .B1(n38), .B2(i_data_bus[48]), 
        .ZN(N108) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[4]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U67 ( .A1(n37), .A2(n33), .B1(n38), .B2(i_data_bus[36]), 
        .ZN(N96) );
  INVD1BWP30P140LVT U68 ( .I(i_data_bus[2]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U69 ( .A1(n37), .A2(n34), .B1(n38), .B2(i_data_bus[34]), 
        .ZN(N94) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[26]), .ZN(n35) );
  MOAI22D1BWP30P140LVT U71 ( .A1(n37), .A2(n35), .B1(n38), .B2(i_data_bus[58]), 
        .ZN(N118) );
  INVD1BWP30P140LVT U72 ( .I(i_data_bus[12]), .ZN(n36) );
  MOAI22D1BWP30P140LVT U73 ( .A1(n37), .A2(n36), .B1(n38), .B2(i_data_bus[44]), 
        .ZN(N104) );
  OR2D1BWP30P140LVT U74 ( .A1(n39), .A2(n38), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_287 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_287 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_0 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_0 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_287 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_286 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_285 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_284 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_283 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_0 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1])
         );
  DFQD1BWP30P140LVT o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0])
         );
  INVD1BWP30P140LVT U3 ( .I(i_valid[1]), .ZN(n9) );
  INR2D1BWP30P140LVT U4 ( .A1(i_en), .B1(rst), .ZN(n7) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(n7), .A2(i_valid[0]), .ZN(n2) );
  NR2D2BWP30P140LVT U6 ( .A1(i_cmd[0]), .A2(n2), .ZN(n5) );
  AOI31D1BWP30P140LVT U7 ( .A1(i_cmd[0]), .A2(n7), .A3(i_valid[1]), .B(n5), 
        .ZN(n1) );
  INVD1BWP30P140LVT U8 ( .I(n1), .ZN(N353) );
  ND3D2BWP30P140LVT U9 ( .A1(n7), .A2(i_cmd[1]), .A3(i_valid[1]), .ZN(n43) );
  OAI21D1BWP30P140LVT U10 ( .A1(i_cmd[1]), .A2(n2), .B(n43), .ZN(N354) );
  INVD1BWP30P140LVT U11 ( .I(i_data_bus[32]), .ZN(n11) );
  INVD1BWP30P140LVT U12 ( .I(n7), .ZN(n3) );
  AOI21D1BWP30P140LVT U13 ( .A1(i_cmd[1]), .A2(n9), .B(n3), .ZN(n4) );
  OAI211OPTREPBD2BWP30P140LVT U14 ( .A1(i_cmd[1]), .A2(i_valid[0]), .B(
        i_cmd[0]), .C(n4), .ZN(n6) );
  MOAI22D1BWP30P140LVT U15 ( .A1(n11), .A2(n6), .B1(i_data_bus[0]), .B2(n5), 
        .ZN(N287) );
  INVD1BWP30P140LVT U16 ( .I(i_data_bus[33]), .ZN(n12) );
  MOAI22D1BWP30P140LVT U17 ( .A1(n6), .A2(n12), .B1(n5), .B2(i_data_bus[1]), 
        .ZN(N288) );
  INVD1BWP30P140LVT U18 ( .I(i_data_bus[34]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U19 ( .A1(n6), .A2(n13), .B1(n5), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140LVT U20 ( .I(i_data_bus[35]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U21 ( .A1(n6), .A2(n14), .B1(n5), .B2(i_data_bus[3]), 
        .ZN(N290) );
  INVD1BWP30P140LVT U22 ( .I(i_data_bus[36]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U23 ( .A1(n6), .A2(n15), .B1(n5), .B2(i_data_bus[4]), 
        .ZN(N291) );
  INVD1BWP30P140LVT U24 ( .I(i_data_bus[37]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U25 ( .A1(n6), .A2(n16), .B1(n5), .B2(i_data_bus[5]), 
        .ZN(N292) );
  INVD1BWP30P140LVT U26 ( .I(i_data_bus[38]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U27 ( .A1(n6), .A2(n17), .B1(n5), .B2(i_data_bus[6]), 
        .ZN(N293) );
  INVD1BWP30P140LVT U28 ( .I(i_data_bus[39]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U29 ( .A1(n6), .A2(n18), .B1(n5), .B2(i_data_bus[7]), 
        .ZN(N294) );
  INVD1BWP30P140LVT U30 ( .I(i_data_bus[40]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U31 ( .A1(n6), .A2(n19), .B1(n5), .B2(i_data_bus[8]), 
        .ZN(N295) );
  INVD1BWP30P140LVT U32 ( .I(i_data_bus[41]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U33 ( .A1(n6), .A2(n20), .B1(n5), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140LVT U34 ( .I(i_data_bus[42]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U35 ( .A1(n6), .A2(n21), .B1(n5), .B2(i_data_bus[10]), 
        .ZN(N297) );
  INVD1BWP30P140LVT U36 ( .I(i_data_bus[43]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U37 ( .A1(n6), .A2(n22), .B1(n5), .B2(i_data_bus[11]), 
        .ZN(N298) );
  INVD1BWP30P140LVT U38 ( .I(i_data_bus[44]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U39 ( .A1(n6), .A2(n23), .B1(n5), .B2(i_data_bus[12]), 
        .ZN(N299) );
  INVD1BWP30P140LVT U40 ( .I(i_data_bus[45]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U41 ( .A1(n6), .A2(n24), .B1(n5), .B2(i_data_bus[13]), 
        .ZN(N300) );
  INVD1BWP30P140LVT U42 ( .I(i_data_bus[46]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U43 ( .A1(n6), .A2(n25), .B1(n5), .B2(i_data_bus[14]), 
        .ZN(N301) );
  INVD1BWP30P140LVT U44 ( .I(i_data_bus[47]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U45 ( .A1(n6), .A2(n26), .B1(n5), .B2(i_data_bus[15]), 
        .ZN(N302) );
  INVD1BWP30P140LVT U46 ( .I(i_data_bus[48]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U47 ( .A1(n6), .A2(n27), .B1(n5), .B2(i_data_bus[16]), 
        .ZN(N303) );
  INVD1BWP30P140LVT U48 ( .I(i_data_bus[49]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U49 ( .A1(n6), .A2(n28), .B1(n5), .B2(i_data_bus[17]), 
        .ZN(N304) );
  INVD1BWP30P140LVT U50 ( .I(i_data_bus[50]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U51 ( .A1(n6), .A2(n29), .B1(n5), .B2(i_data_bus[18]), 
        .ZN(N305) );
  INVD1BWP30P140LVT U52 ( .I(i_data_bus[51]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U53 ( .A1(n6), .A2(n30), .B1(n5), .B2(i_data_bus[19]), 
        .ZN(N306) );
  INVD1BWP30P140LVT U54 ( .I(i_data_bus[52]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U55 ( .A1(n6), .A2(n31), .B1(n5), .B2(i_data_bus[20]), 
        .ZN(N307) );
  INVD1BWP30P140LVT U56 ( .I(i_data_bus[53]), .ZN(n32) );
  MOAI22D1BWP30P140LVT U57 ( .A1(n6), .A2(n32), .B1(n5), .B2(i_data_bus[21]), 
        .ZN(N308) );
  INVD1BWP30P140LVT U58 ( .I(i_data_bus[54]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U59 ( .A1(n6), .A2(n33), .B1(n5), .B2(i_data_bus[22]), 
        .ZN(N309) );
  INVD1BWP30P140LVT U60 ( .I(i_data_bus[55]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U61 ( .A1(n6), .A2(n34), .B1(n5), .B2(i_data_bus[23]), 
        .ZN(N310) );
  INVD1BWP30P140LVT U62 ( .I(i_data_bus[56]), .ZN(n35) );
  MOAI22D1BWP30P140LVT U63 ( .A1(n6), .A2(n35), .B1(n5), .B2(i_data_bus[24]), 
        .ZN(N311) );
  INVD1BWP30P140LVT U64 ( .I(i_data_bus[57]), .ZN(n36) );
  MOAI22D1BWP30P140LVT U65 ( .A1(n6), .A2(n36), .B1(n5), .B2(i_data_bus[25]), 
        .ZN(N312) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[58]), .ZN(n37) );
  MOAI22D1BWP30P140LVT U67 ( .A1(n6), .A2(n37), .B1(n5), .B2(i_data_bus[26]), 
        .ZN(N313) );
  INVD1BWP30P140LVT U68 ( .I(i_data_bus[59]), .ZN(n38) );
  MOAI22D1BWP30P140LVT U69 ( .A1(n6), .A2(n38), .B1(n5), .B2(i_data_bus[27]), 
        .ZN(N314) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[60]), .ZN(n39) );
  MOAI22D1BWP30P140LVT U71 ( .A1(n6), .A2(n39), .B1(n5), .B2(i_data_bus[28]), 
        .ZN(N315) );
  INVD1BWP30P140LVT U72 ( .I(i_data_bus[61]), .ZN(n40) );
  MOAI22D1BWP30P140LVT U73 ( .A1(n6), .A2(n40), .B1(n5), .B2(i_data_bus[29]), 
        .ZN(N316) );
  INVD1BWP30P140LVT U74 ( .I(i_data_bus[62]), .ZN(n41) );
  MOAI22D1BWP30P140LVT U75 ( .A1(n6), .A2(n41), .B1(n5), .B2(i_data_bus[30]), 
        .ZN(N317) );
  INVD1BWP30P140LVT U76 ( .I(i_data_bus[63]), .ZN(n44) );
  MOAI22D1BWP30P140LVT U77 ( .A1(n6), .A2(n44), .B1(n5), .B2(i_data_bus[31]), 
        .ZN(N318) );
  OAI21D1BWP30P140LVT U78 ( .A1(i_cmd[0]), .A2(i_valid[0]), .B(n7), .ZN(n8) );
  AO211D1BWP30P140LVT U79 ( .A1(i_cmd[0]), .A2(n9), .B(i_cmd[1]), .C(n8), .Z(
        n10) );
  INVD2BWP30P140LVT U80 ( .I(n10), .ZN(n42) );
  MOAI22D1BWP30P140LVT U81 ( .A1(n11), .A2(n43), .B1(i_data_bus[0]), .B2(n42), 
        .ZN(N319) );
  MOAI22D1BWP30P140LVT U82 ( .A1(n12), .A2(n43), .B1(i_data_bus[1]), .B2(n42), 
        .ZN(N320) );
  MOAI22D1BWP30P140LVT U83 ( .A1(n13), .A2(n43), .B1(i_data_bus[2]), .B2(n42), 
        .ZN(N321) );
  MOAI22D1BWP30P140LVT U84 ( .A1(n14), .A2(n43), .B1(i_data_bus[3]), .B2(n42), 
        .ZN(N322) );
  MOAI22D1BWP30P140LVT U85 ( .A1(n15), .A2(n43), .B1(i_data_bus[4]), .B2(n42), 
        .ZN(N323) );
  MOAI22D1BWP30P140LVT U86 ( .A1(n16), .A2(n43), .B1(i_data_bus[5]), .B2(n42), 
        .ZN(N324) );
  MOAI22D1BWP30P140LVT U87 ( .A1(n17), .A2(n43), .B1(i_data_bus[6]), .B2(n42), 
        .ZN(N325) );
  MOAI22D1BWP30P140LVT U88 ( .A1(n18), .A2(n43), .B1(i_data_bus[7]), .B2(n42), 
        .ZN(N326) );
  MOAI22D1BWP30P140LVT U89 ( .A1(n19), .A2(n43), .B1(i_data_bus[8]), .B2(n42), 
        .ZN(N327) );
  MOAI22D1BWP30P140LVT U90 ( .A1(n20), .A2(n43), .B1(i_data_bus[9]), .B2(n42), 
        .ZN(N328) );
  MOAI22D1BWP30P140LVT U91 ( .A1(n21), .A2(n43), .B1(i_data_bus[10]), .B2(n42), 
        .ZN(N329) );
  MOAI22D1BWP30P140LVT U92 ( .A1(n22), .A2(n43), .B1(i_data_bus[11]), .B2(n42), 
        .ZN(N330) );
  MOAI22D1BWP30P140LVT U93 ( .A1(n23), .A2(n43), .B1(i_data_bus[12]), .B2(n42), 
        .ZN(N331) );
  MOAI22D1BWP30P140LVT U94 ( .A1(n24), .A2(n43), .B1(i_data_bus[13]), .B2(n42), 
        .ZN(N332) );
  MOAI22D1BWP30P140LVT U95 ( .A1(n25), .A2(n43), .B1(i_data_bus[14]), .B2(n42), 
        .ZN(N333) );
  MOAI22D1BWP30P140LVT U96 ( .A1(n26), .A2(n43), .B1(i_data_bus[15]), .B2(n42), 
        .ZN(N334) );
  MOAI22D1BWP30P140LVT U97 ( .A1(n27), .A2(n43), .B1(i_data_bus[16]), .B2(n42), 
        .ZN(N335) );
  MOAI22D1BWP30P140LVT U98 ( .A1(n28), .A2(n43), .B1(i_data_bus[17]), .B2(n42), 
        .ZN(N336) );
  MOAI22D1BWP30P140LVT U99 ( .A1(n29), .A2(n43), .B1(i_data_bus[18]), .B2(n42), 
        .ZN(N337) );
  MOAI22D1BWP30P140LVT U100 ( .A1(n30), .A2(n43), .B1(i_data_bus[19]), .B2(n42), .ZN(N338) );
  MOAI22D1BWP30P140LVT U101 ( .A1(n31), .A2(n43), .B1(i_data_bus[20]), .B2(n42), .ZN(N339) );
  MOAI22D1BWP30P140LVT U102 ( .A1(n32), .A2(n43), .B1(i_data_bus[21]), .B2(n42), .ZN(N340) );
  MOAI22D1BWP30P140LVT U103 ( .A1(n33), .A2(n43), .B1(i_data_bus[22]), .B2(n42), .ZN(N341) );
  MOAI22D1BWP30P140LVT U104 ( .A1(n34), .A2(n43), .B1(i_data_bus[23]), .B2(n42), .ZN(N342) );
  MOAI22D1BWP30P140LVT U105 ( .A1(n35), .A2(n43), .B1(i_data_bus[24]), .B2(n42), .ZN(N343) );
  MOAI22D1BWP30P140LVT U106 ( .A1(n36), .A2(n43), .B1(i_data_bus[25]), .B2(n42), .ZN(N344) );
  MOAI22D1BWP30P140LVT U107 ( .A1(n37), .A2(n43), .B1(i_data_bus[26]), .B2(n42), .ZN(N345) );
  MOAI22D1BWP30P140LVT U108 ( .A1(n38), .A2(n43), .B1(i_data_bus[27]), .B2(n42), .ZN(N346) );
  MOAI22D1BWP30P140LVT U109 ( .A1(n39), .A2(n43), .B1(i_data_bus[28]), .B2(n42), .ZN(N347) );
  MOAI22D1BWP30P140LVT U110 ( .A1(n40), .A2(n43), .B1(i_data_bus[29]), .B2(n42), .ZN(N348) );
  MOAI22D1BWP30P140LVT U111 ( .A1(n41), .A2(n43), .B1(i_data_bus[30]), .B2(n42), .ZN(N349) );
  MOAI22D1BWP30P140LVT U112 ( .A1(n44), .A2(n43), .B1(i_data_bus[31]), .B2(n42), .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_1 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1])
         );
  DFQD1BWP30P140LVT o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0])
         );
  INVD1BWP30P140LVT U3 ( .I(i_valid[1]), .ZN(n9) );
  INR2D1BWP30P140LVT U4 ( .A1(i_en), .B1(rst), .ZN(n7) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(n7), .A2(i_valid[0]), .ZN(n2) );
  NR2D2BWP30P140LVT U6 ( .A1(i_cmd[0]), .A2(n2), .ZN(n5) );
  AOI31D1BWP30P140LVT U7 ( .A1(i_cmd[0]), .A2(n7), .A3(i_valid[1]), .B(n5), 
        .ZN(n1) );
  INVD1BWP30P140LVT U8 ( .I(n1), .ZN(N353) );
  ND3D2BWP30P140LVT U9 ( .A1(n7), .A2(i_cmd[1]), .A3(i_valid[1]), .ZN(n43) );
  OAI21D1BWP30P140LVT U10 ( .A1(i_cmd[1]), .A2(n2), .B(n43), .ZN(N354) );
  INVD1BWP30P140LVT U11 ( .I(i_data_bus[32]), .ZN(n11) );
  INVD1BWP30P140LVT U12 ( .I(n7), .ZN(n3) );
  AOI21D1BWP30P140LVT U13 ( .A1(i_cmd[1]), .A2(n9), .B(n3), .ZN(n4) );
  OAI211OPTREPBD2BWP30P140LVT U14 ( .A1(i_cmd[1]), .A2(i_valid[0]), .B(
        i_cmd[0]), .C(n4), .ZN(n6) );
  MOAI22D1BWP30P140LVT U15 ( .A1(n11), .A2(n6), .B1(i_data_bus[0]), .B2(n5), 
        .ZN(N287) );
  INVD1BWP30P140LVT U16 ( .I(i_data_bus[33]), .ZN(n12) );
  MOAI22D1BWP30P140LVT U17 ( .A1(n6), .A2(n12), .B1(n5), .B2(i_data_bus[1]), 
        .ZN(N288) );
  INVD1BWP30P140LVT U18 ( .I(i_data_bus[34]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U19 ( .A1(n6), .A2(n13), .B1(n5), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140LVT U20 ( .I(i_data_bus[35]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U21 ( .A1(n6), .A2(n14), .B1(n5), .B2(i_data_bus[3]), 
        .ZN(N290) );
  INVD1BWP30P140LVT U22 ( .I(i_data_bus[36]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U23 ( .A1(n6), .A2(n15), .B1(n5), .B2(i_data_bus[4]), 
        .ZN(N291) );
  INVD1BWP30P140LVT U24 ( .I(i_data_bus[37]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U25 ( .A1(n6), .A2(n16), .B1(n5), .B2(i_data_bus[5]), 
        .ZN(N292) );
  INVD1BWP30P140LVT U26 ( .I(i_data_bus[38]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U27 ( .A1(n6), .A2(n17), .B1(n5), .B2(i_data_bus[6]), 
        .ZN(N293) );
  INVD1BWP30P140LVT U28 ( .I(i_data_bus[39]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U29 ( .A1(n6), .A2(n18), .B1(n5), .B2(i_data_bus[7]), 
        .ZN(N294) );
  INVD1BWP30P140LVT U30 ( .I(i_data_bus[40]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U31 ( .A1(n6), .A2(n19), .B1(n5), .B2(i_data_bus[8]), 
        .ZN(N295) );
  INVD1BWP30P140LVT U32 ( .I(i_data_bus[41]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U33 ( .A1(n6), .A2(n20), .B1(n5), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140LVT U34 ( .I(i_data_bus[42]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U35 ( .A1(n6), .A2(n21), .B1(n5), .B2(i_data_bus[10]), 
        .ZN(N297) );
  INVD1BWP30P140LVT U36 ( .I(i_data_bus[43]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U37 ( .A1(n6), .A2(n22), .B1(n5), .B2(i_data_bus[11]), 
        .ZN(N298) );
  INVD1BWP30P140LVT U38 ( .I(i_data_bus[44]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U39 ( .A1(n6), .A2(n23), .B1(n5), .B2(i_data_bus[12]), 
        .ZN(N299) );
  INVD1BWP30P140LVT U40 ( .I(i_data_bus[45]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U41 ( .A1(n6), .A2(n24), .B1(n5), .B2(i_data_bus[13]), 
        .ZN(N300) );
  INVD1BWP30P140LVT U42 ( .I(i_data_bus[46]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U43 ( .A1(n6), .A2(n25), .B1(n5), .B2(i_data_bus[14]), 
        .ZN(N301) );
  INVD1BWP30P140LVT U44 ( .I(i_data_bus[47]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U45 ( .A1(n6), .A2(n26), .B1(n5), .B2(i_data_bus[15]), 
        .ZN(N302) );
  INVD1BWP30P140LVT U46 ( .I(i_data_bus[48]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U47 ( .A1(n6), .A2(n27), .B1(n5), .B2(i_data_bus[16]), 
        .ZN(N303) );
  INVD1BWP30P140LVT U48 ( .I(i_data_bus[49]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U49 ( .A1(n6), .A2(n28), .B1(n5), .B2(i_data_bus[17]), 
        .ZN(N304) );
  INVD1BWP30P140LVT U50 ( .I(i_data_bus[50]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U51 ( .A1(n6), .A2(n29), .B1(n5), .B2(i_data_bus[18]), 
        .ZN(N305) );
  INVD1BWP30P140LVT U52 ( .I(i_data_bus[51]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U53 ( .A1(n6), .A2(n30), .B1(n5), .B2(i_data_bus[19]), 
        .ZN(N306) );
  INVD1BWP30P140LVT U54 ( .I(i_data_bus[52]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U55 ( .A1(n6), .A2(n31), .B1(n5), .B2(i_data_bus[20]), 
        .ZN(N307) );
  INVD1BWP30P140LVT U56 ( .I(i_data_bus[53]), .ZN(n32) );
  MOAI22D1BWP30P140LVT U57 ( .A1(n6), .A2(n32), .B1(n5), .B2(i_data_bus[21]), 
        .ZN(N308) );
  INVD1BWP30P140LVT U58 ( .I(i_data_bus[54]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U59 ( .A1(n6), .A2(n33), .B1(n5), .B2(i_data_bus[22]), 
        .ZN(N309) );
  INVD1BWP30P140LVT U60 ( .I(i_data_bus[55]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U61 ( .A1(n6), .A2(n34), .B1(n5), .B2(i_data_bus[23]), 
        .ZN(N310) );
  INVD1BWP30P140LVT U62 ( .I(i_data_bus[56]), .ZN(n35) );
  MOAI22D1BWP30P140LVT U63 ( .A1(n6), .A2(n35), .B1(n5), .B2(i_data_bus[24]), 
        .ZN(N311) );
  INVD1BWP30P140LVT U64 ( .I(i_data_bus[57]), .ZN(n36) );
  MOAI22D1BWP30P140LVT U65 ( .A1(n6), .A2(n36), .B1(n5), .B2(i_data_bus[25]), 
        .ZN(N312) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[58]), .ZN(n37) );
  MOAI22D1BWP30P140LVT U67 ( .A1(n6), .A2(n37), .B1(n5), .B2(i_data_bus[26]), 
        .ZN(N313) );
  INVD1BWP30P140LVT U68 ( .I(i_data_bus[59]), .ZN(n38) );
  MOAI22D1BWP30P140LVT U69 ( .A1(n6), .A2(n38), .B1(n5), .B2(i_data_bus[27]), 
        .ZN(N314) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[60]), .ZN(n39) );
  MOAI22D1BWP30P140LVT U71 ( .A1(n6), .A2(n39), .B1(n5), .B2(i_data_bus[28]), 
        .ZN(N315) );
  INVD1BWP30P140LVT U72 ( .I(i_data_bus[61]), .ZN(n40) );
  MOAI22D1BWP30P140LVT U73 ( .A1(n6), .A2(n40), .B1(n5), .B2(i_data_bus[29]), 
        .ZN(N316) );
  INVD1BWP30P140LVT U74 ( .I(i_data_bus[62]), .ZN(n41) );
  MOAI22D1BWP30P140LVT U75 ( .A1(n6), .A2(n41), .B1(n5), .B2(i_data_bus[30]), 
        .ZN(N317) );
  INVD1BWP30P140LVT U76 ( .I(i_data_bus[63]), .ZN(n44) );
  MOAI22D1BWP30P140LVT U77 ( .A1(n6), .A2(n44), .B1(n5), .B2(i_data_bus[31]), 
        .ZN(N318) );
  OAI21D1BWP30P140LVT U78 ( .A1(i_cmd[0]), .A2(i_valid[0]), .B(n7), .ZN(n8) );
  AO211D1BWP30P140LVT U79 ( .A1(i_cmd[0]), .A2(n9), .B(i_cmd[1]), .C(n8), .Z(
        n10) );
  INVD2BWP30P140LVT U80 ( .I(n10), .ZN(n42) );
  MOAI22D1BWP30P140LVT U81 ( .A1(n11), .A2(n43), .B1(i_data_bus[0]), .B2(n42), 
        .ZN(N319) );
  MOAI22D1BWP30P140LVT U82 ( .A1(n12), .A2(n43), .B1(i_data_bus[1]), .B2(n42), 
        .ZN(N320) );
  MOAI22D1BWP30P140LVT U83 ( .A1(n13), .A2(n43), .B1(i_data_bus[2]), .B2(n42), 
        .ZN(N321) );
  MOAI22D1BWP30P140LVT U84 ( .A1(n14), .A2(n43), .B1(i_data_bus[3]), .B2(n42), 
        .ZN(N322) );
  MOAI22D1BWP30P140LVT U85 ( .A1(n15), .A2(n43), .B1(i_data_bus[4]), .B2(n42), 
        .ZN(N323) );
  MOAI22D1BWP30P140LVT U86 ( .A1(n16), .A2(n43), .B1(i_data_bus[5]), .B2(n42), 
        .ZN(N324) );
  MOAI22D1BWP30P140LVT U87 ( .A1(n17), .A2(n43), .B1(i_data_bus[6]), .B2(n42), 
        .ZN(N325) );
  MOAI22D1BWP30P140LVT U88 ( .A1(n18), .A2(n43), .B1(i_data_bus[7]), .B2(n42), 
        .ZN(N326) );
  MOAI22D1BWP30P140LVT U89 ( .A1(n19), .A2(n43), .B1(i_data_bus[8]), .B2(n42), 
        .ZN(N327) );
  MOAI22D1BWP30P140LVT U90 ( .A1(n20), .A2(n43), .B1(i_data_bus[9]), .B2(n42), 
        .ZN(N328) );
  MOAI22D1BWP30P140LVT U91 ( .A1(n21), .A2(n43), .B1(i_data_bus[10]), .B2(n42), 
        .ZN(N329) );
  MOAI22D1BWP30P140LVT U92 ( .A1(n22), .A2(n43), .B1(i_data_bus[11]), .B2(n42), 
        .ZN(N330) );
  MOAI22D1BWP30P140LVT U93 ( .A1(n23), .A2(n43), .B1(i_data_bus[12]), .B2(n42), 
        .ZN(N331) );
  MOAI22D1BWP30P140LVT U94 ( .A1(n24), .A2(n43), .B1(i_data_bus[13]), .B2(n42), 
        .ZN(N332) );
  MOAI22D1BWP30P140LVT U95 ( .A1(n25), .A2(n43), .B1(i_data_bus[14]), .B2(n42), 
        .ZN(N333) );
  MOAI22D1BWP30P140LVT U96 ( .A1(n26), .A2(n43), .B1(i_data_bus[15]), .B2(n42), 
        .ZN(N334) );
  MOAI22D1BWP30P140LVT U97 ( .A1(n27), .A2(n43), .B1(i_data_bus[16]), .B2(n42), 
        .ZN(N335) );
  MOAI22D1BWP30P140LVT U98 ( .A1(n28), .A2(n43), .B1(i_data_bus[17]), .B2(n42), 
        .ZN(N336) );
  MOAI22D1BWP30P140LVT U99 ( .A1(n29), .A2(n43), .B1(i_data_bus[18]), .B2(n42), 
        .ZN(N337) );
  MOAI22D1BWP30P140LVT U100 ( .A1(n30), .A2(n43), .B1(i_data_bus[19]), .B2(n42), .ZN(N338) );
  MOAI22D1BWP30P140LVT U101 ( .A1(n31), .A2(n43), .B1(i_data_bus[20]), .B2(n42), .ZN(N339) );
  MOAI22D1BWP30P140LVT U102 ( .A1(n32), .A2(n43), .B1(i_data_bus[21]), .B2(n42), .ZN(N340) );
  MOAI22D1BWP30P140LVT U103 ( .A1(n33), .A2(n43), .B1(i_data_bus[22]), .B2(n42), .ZN(N341) );
  MOAI22D1BWP30P140LVT U104 ( .A1(n34), .A2(n43), .B1(i_data_bus[23]), .B2(n42), .ZN(N342) );
  MOAI22D1BWP30P140LVT U105 ( .A1(n35), .A2(n43), .B1(i_data_bus[24]), .B2(n42), .ZN(N343) );
  MOAI22D1BWP30P140LVT U106 ( .A1(n36), .A2(n43), .B1(i_data_bus[25]), .B2(n42), .ZN(N344) );
  MOAI22D1BWP30P140LVT U107 ( .A1(n37), .A2(n43), .B1(i_data_bus[26]), .B2(n42), .ZN(N345) );
  MOAI22D1BWP30P140LVT U108 ( .A1(n38), .A2(n43), .B1(i_data_bus[27]), .B2(n42), .ZN(N346) );
  MOAI22D1BWP30P140LVT U109 ( .A1(n39), .A2(n43), .B1(i_data_bus[28]), .B2(n42), .ZN(N347) );
  MOAI22D1BWP30P140LVT U110 ( .A1(n40), .A2(n43), .B1(i_data_bus[29]), .B2(n42), .ZN(N348) );
  MOAI22D1BWP30P140LVT U111 ( .A1(n41), .A2(n43), .B1(i_data_bus[30]), .B2(n42), .ZN(N349) );
  MOAI22D1BWP30P140LVT U112 ( .A1(n44), .A2(n43), .B1(i_data_bus[31]), .B2(n42), .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_2 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1])
         );
  DFQD1BWP30P140LVT o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0])
         );
  INVD1BWP30P140LVT U3 ( .I(i_valid[1]), .ZN(n9) );
  INR2D1BWP30P140LVT U4 ( .A1(i_en), .B1(rst), .ZN(n7) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(n7), .A2(i_valid[0]), .ZN(n2) );
  NR2D2BWP30P140LVT U6 ( .A1(i_cmd[0]), .A2(n2), .ZN(n5) );
  AOI31D1BWP30P140LVT U7 ( .A1(i_cmd[0]), .A2(n7), .A3(i_valid[1]), .B(n5), 
        .ZN(n1) );
  INVD1BWP30P140LVT U8 ( .I(n1), .ZN(N353) );
  ND3D2BWP30P140LVT U9 ( .A1(n7), .A2(i_cmd[1]), .A3(i_valid[1]), .ZN(n43) );
  OAI21D1BWP30P140LVT U10 ( .A1(i_cmd[1]), .A2(n2), .B(n43), .ZN(N354) );
  INVD1BWP30P140LVT U11 ( .I(i_data_bus[32]), .ZN(n11) );
  INVD1BWP30P140LVT U12 ( .I(n7), .ZN(n3) );
  AOI21D1BWP30P140LVT U13 ( .A1(i_cmd[1]), .A2(n9), .B(n3), .ZN(n4) );
  OAI211OPTREPBD2BWP30P140LVT U14 ( .A1(i_cmd[1]), .A2(i_valid[0]), .B(
        i_cmd[0]), .C(n4), .ZN(n6) );
  MOAI22D1BWP30P140LVT U15 ( .A1(n11), .A2(n6), .B1(i_data_bus[0]), .B2(n5), 
        .ZN(N287) );
  INVD1BWP30P140LVT U16 ( .I(i_data_bus[33]), .ZN(n12) );
  MOAI22D1BWP30P140LVT U17 ( .A1(n6), .A2(n12), .B1(n5), .B2(i_data_bus[1]), 
        .ZN(N288) );
  INVD1BWP30P140LVT U18 ( .I(i_data_bus[34]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U19 ( .A1(n6), .A2(n13), .B1(n5), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140LVT U20 ( .I(i_data_bus[35]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U21 ( .A1(n6), .A2(n14), .B1(n5), .B2(i_data_bus[3]), 
        .ZN(N290) );
  INVD1BWP30P140LVT U22 ( .I(i_data_bus[36]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U23 ( .A1(n6), .A2(n15), .B1(n5), .B2(i_data_bus[4]), 
        .ZN(N291) );
  INVD1BWP30P140LVT U24 ( .I(i_data_bus[37]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U25 ( .A1(n6), .A2(n16), .B1(n5), .B2(i_data_bus[5]), 
        .ZN(N292) );
  INVD1BWP30P140LVT U26 ( .I(i_data_bus[38]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U27 ( .A1(n6), .A2(n17), .B1(n5), .B2(i_data_bus[6]), 
        .ZN(N293) );
  INVD1BWP30P140LVT U28 ( .I(i_data_bus[39]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U29 ( .A1(n6), .A2(n18), .B1(n5), .B2(i_data_bus[7]), 
        .ZN(N294) );
  INVD1BWP30P140LVT U30 ( .I(i_data_bus[40]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U31 ( .A1(n6), .A2(n19), .B1(n5), .B2(i_data_bus[8]), 
        .ZN(N295) );
  INVD1BWP30P140LVT U32 ( .I(i_data_bus[41]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U33 ( .A1(n6), .A2(n20), .B1(n5), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140LVT U34 ( .I(i_data_bus[42]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U35 ( .A1(n6), .A2(n21), .B1(n5), .B2(i_data_bus[10]), 
        .ZN(N297) );
  INVD1BWP30P140LVT U36 ( .I(i_data_bus[43]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U37 ( .A1(n6), .A2(n22), .B1(n5), .B2(i_data_bus[11]), 
        .ZN(N298) );
  INVD1BWP30P140LVT U38 ( .I(i_data_bus[44]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U39 ( .A1(n6), .A2(n23), .B1(n5), .B2(i_data_bus[12]), 
        .ZN(N299) );
  INVD1BWP30P140LVT U40 ( .I(i_data_bus[45]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U41 ( .A1(n6), .A2(n24), .B1(n5), .B2(i_data_bus[13]), 
        .ZN(N300) );
  INVD1BWP30P140LVT U42 ( .I(i_data_bus[46]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U43 ( .A1(n6), .A2(n25), .B1(n5), .B2(i_data_bus[14]), 
        .ZN(N301) );
  INVD1BWP30P140LVT U44 ( .I(i_data_bus[47]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U45 ( .A1(n6), .A2(n26), .B1(n5), .B2(i_data_bus[15]), 
        .ZN(N302) );
  INVD1BWP30P140LVT U46 ( .I(i_data_bus[48]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U47 ( .A1(n6), .A2(n27), .B1(n5), .B2(i_data_bus[16]), 
        .ZN(N303) );
  INVD1BWP30P140LVT U48 ( .I(i_data_bus[49]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U49 ( .A1(n6), .A2(n28), .B1(n5), .B2(i_data_bus[17]), 
        .ZN(N304) );
  INVD1BWP30P140LVT U50 ( .I(i_data_bus[50]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U51 ( .A1(n6), .A2(n29), .B1(n5), .B2(i_data_bus[18]), 
        .ZN(N305) );
  INVD1BWP30P140LVT U52 ( .I(i_data_bus[51]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U53 ( .A1(n6), .A2(n30), .B1(n5), .B2(i_data_bus[19]), 
        .ZN(N306) );
  INVD1BWP30P140LVT U54 ( .I(i_data_bus[52]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U55 ( .A1(n6), .A2(n31), .B1(n5), .B2(i_data_bus[20]), 
        .ZN(N307) );
  INVD1BWP30P140LVT U56 ( .I(i_data_bus[53]), .ZN(n32) );
  MOAI22D1BWP30P140LVT U57 ( .A1(n6), .A2(n32), .B1(n5), .B2(i_data_bus[21]), 
        .ZN(N308) );
  INVD1BWP30P140LVT U58 ( .I(i_data_bus[54]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U59 ( .A1(n6), .A2(n33), .B1(n5), .B2(i_data_bus[22]), 
        .ZN(N309) );
  INVD1BWP30P140LVT U60 ( .I(i_data_bus[55]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U61 ( .A1(n6), .A2(n34), .B1(n5), .B2(i_data_bus[23]), 
        .ZN(N310) );
  INVD1BWP30P140LVT U62 ( .I(i_data_bus[56]), .ZN(n35) );
  MOAI22D1BWP30P140LVT U63 ( .A1(n6), .A2(n35), .B1(n5), .B2(i_data_bus[24]), 
        .ZN(N311) );
  INVD1BWP30P140LVT U64 ( .I(i_data_bus[57]), .ZN(n36) );
  MOAI22D1BWP30P140LVT U65 ( .A1(n6), .A2(n36), .B1(n5), .B2(i_data_bus[25]), 
        .ZN(N312) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[58]), .ZN(n37) );
  MOAI22D1BWP30P140LVT U67 ( .A1(n6), .A2(n37), .B1(n5), .B2(i_data_bus[26]), 
        .ZN(N313) );
  INVD1BWP30P140LVT U68 ( .I(i_data_bus[59]), .ZN(n38) );
  MOAI22D1BWP30P140LVT U69 ( .A1(n6), .A2(n38), .B1(n5), .B2(i_data_bus[27]), 
        .ZN(N314) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[60]), .ZN(n39) );
  MOAI22D1BWP30P140LVT U71 ( .A1(n6), .A2(n39), .B1(n5), .B2(i_data_bus[28]), 
        .ZN(N315) );
  INVD1BWP30P140LVT U72 ( .I(i_data_bus[61]), .ZN(n40) );
  MOAI22D1BWP30P140LVT U73 ( .A1(n6), .A2(n40), .B1(n5), .B2(i_data_bus[29]), 
        .ZN(N316) );
  INVD1BWP30P140LVT U74 ( .I(i_data_bus[62]), .ZN(n41) );
  MOAI22D1BWP30P140LVT U75 ( .A1(n6), .A2(n41), .B1(n5), .B2(i_data_bus[30]), 
        .ZN(N317) );
  INVD1BWP30P140LVT U76 ( .I(i_data_bus[63]), .ZN(n44) );
  MOAI22D1BWP30P140LVT U77 ( .A1(n6), .A2(n44), .B1(n5), .B2(i_data_bus[31]), 
        .ZN(N318) );
  OAI21D1BWP30P140LVT U78 ( .A1(i_cmd[0]), .A2(i_valid[0]), .B(n7), .ZN(n8) );
  AO211D1BWP30P140LVT U79 ( .A1(i_cmd[0]), .A2(n9), .B(i_cmd[1]), .C(n8), .Z(
        n10) );
  INVD2BWP30P140LVT U80 ( .I(n10), .ZN(n42) );
  MOAI22D1BWP30P140LVT U81 ( .A1(n11), .A2(n43), .B1(i_data_bus[0]), .B2(n42), 
        .ZN(N319) );
  MOAI22D1BWP30P140LVT U82 ( .A1(n12), .A2(n43), .B1(i_data_bus[1]), .B2(n42), 
        .ZN(N320) );
  MOAI22D1BWP30P140LVT U83 ( .A1(n13), .A2(n43), .B1(i_data_bus[2]), .B2(n42), 
        .ZN(N321) );
  MOAI22D1BWP30P140LVT U84 ( .A1(n14), .A2(n43), .B1(i_data_bus[3]), .B2(n42), 
        .ZN(N322) );
  MOAI22D1BWP30P140LVT U85 ( .A1(n15), .A2(n43), .B1(i_data_bus[4]), .B2(n42), 
        .ZN(N323) );
  MOAI22D1BWP30P140LVT U86 ( .A1(n16), .A2(n43), .B1(i_data_bus[5]), .B2(n42), 
        .ZN(N324) );
  MOAI22D1BWP30P140LVT U87 ( .A1(n17), .A2(n43), .B1(i_data_bus[6]), .B2(n42), 
        .ZN(N325) );
  MOAI22D1BWP30P140LVT U88 ( .A1(n18), .A2(n43), .B1(i_data_bus[7]), .B2(n42), 
        .ZN(N326) );
  MOAI22D1BWP30P140LVT U89 ( .A1(n19), .A2(n43), .B1(i_data_bus[8]), .B2(n42), 
        .ZN(N327) );
  MOAI22D1BWP30P140LVT U90 ( .A1(n20), .A2(n43), .B1(i_data_bus[9]), .B2(n42), 
        .ZN(N328) );
  MOAI22D1BWP30P140LVT U91 ( .A1(n21), .A2(n43), .B1(i_data_bus[10]), .B2(n42), 
        .ZN(N329) );
  MOAI22D1BWP30P140LVT U92 ( .A1(n22), .A2(n43), .B1(i_data_bus[11]), .B2(n42), 
        .ZN(N330) );
  MOAI22D1BWP30P140LVT U93 ( .A1(n23), .A2(n43), .B1(i_data_bus[12]), .B2(n42), 
        .ZN(N331) );
  MOAI22D1BWP30P140LVT U94 ( .A1(n24), .A2(n43), .B1(i_data_bus[13]), .B2(n42), 
        .ZN(N332) );
  MOAI22D1BWP30P140LVT U95 ( .A1(n25), .A2(n43), .B1(i_data_bus[14]), .B2(n42), 
        .ZN(N333) );
  MOAI22D1BWP30P140LVT U96 ( .A1(n26), .A2(n43), .B1(i_data_bus[15]), .B2(n42), 
        .ZN(N334) );
  MOAI22D1BWP30P140LVT U97 ( .A1(n27), .A2(n43), .B1(i_data_bus[16]), .B2(n42), 
        .ZN(N335) );
  MOAI22D1BWP30P140LVT U98 ( .A1(n28), .A2(n43), .B1(i_data_bus[17]), .B2(n42), 
        .ZN(N336) );
  MOAI22D1BWP30P140LVT U99 ( .A1(n29), .A2(n43), .B1(i_data_bus[18]), .B2(n42), 
        .ZN(N337) );
  MOAI22D1BWP30P140LVT U100 ( .A1(n30), .A2(n43), .B1(i_data_bus[19]), .B2(n42), .ZN(N338) );
  MOAI22D1BWP30P140LVT U101 ( .A1(n31), .A2(n43), .B1(i_data_bus[20]), .B2(n42), .ZN(N339) );
  MOAI22D1BWP30P140LVT U102 ( .A1(n32), .A2(n43), .B1(i_data_bus[21]), .B2(n42), .ZN(N340) );
  MOAI22D1BWP30P140LVT U103 ( .A1(n33), .A2(n43), .B1(i_data_bus[22]), .B2(n42), .ZN(N341) );
  MOAI22D1BWP30P140LVT U104 ( .A1(n34), .A2(n43), .B1(i_data_bus[23]), .B2(n42), .ZN(N342) );
  MOAI22D1BWP30P140LVT U105 ( .A1(n35), .A2(n43), .B1(i_data_bus[24]), .B2(n42), .ZN(N343) );
  MOAI22D1BWP30P140LVT U106 ( .A1(n36), .A2(n43), .B1(i_data_bus[25]), .B2(n42), .ZN(N344) );
  MOAI22D1BWP30P140LVT U107 ( .A1(n37), .A2(n43), .B1(i_data_bus[26]), .B2(n42), .ZN(N345) );
  MOAI22D1BWP30P140LVT U108 ( .A1(n38), .A2(n43), .B1(i_data_bus[27]), .B2(n42), .ZN(N346) );
  MOAI22D1BWP30P140LVT U109 ( .A1(n39), .A2(n43), .B1(i_data_bus[28]), .B2(n42), .ZN(N347) );
  MOAI22D1BWP30P140LVT U110 ( .A1(n40), .A2(n43), .B1(i_data_bus[29]), .B2(n42), .ZN(N348) );
  MOAI22D1BWP30P140LVT U111 ( .A1(n41), .A2(n43), .B1(i_data_bus[30]), .B2(n42), .ZN(N349) );
  MOAI22D1BWP30P140LVT U112 ( .A1(n44), .A2(n43), .B1(i_data_bus[31]), .B2(n42), .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_3 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1])
         );
  DFQD1BWP30P140LVT o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0])
         );
  INVD1BWP30P140LVT U3 ( .I(i_valid[1]), .ZN(n9) );
  INR2D1BWP30P140LVT U4 ( .A1(i_en), .B1(rst), .ZN(n7) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(n7), .A2(i_valid[0]), .ZN(n2) );
  NR2D2BWP30P140LVT U6 ( .A1(i_cmd[0]), .A2(n2), .ZN(n5) );
  AOI31D1BWP30P140LVT U7 ( .A1(i_cmd[0]), .A2(n7), .A3(i_valid[1]), .B(n5), 
        .ZN(n1) );
  INVD1BWP30P140LVT U8 ( .I(n1), .ZN(N353) );
  ND3D2BWP30P140LVT U9 ( .A1(n7), .A2(i_cmd[1]), .A3(i_valid[1]), .ZN(n43) );
  OAI21D1BWP30P140LVT U10 ( .A1(i_cmd[1]), .A2(n2), .B(n43), .ZN(N354) );
  INVD1BWP30P140LVT U11 ( .I(i_data_bus[32]), .ZN(n11) );
  INVD1BWP30P140LVT U12 ( .I(n7), .ZN(n3) );
  AOI21D1BWP30P140LVT U13 ( .A1(i_cmd[1]), .A2(n9), .B(n3), .ZN(n4) );
  OAI211OPTREPBD2BWP30P140LVT U14 ( .A1(i_cmd[1]), .A2(i_valid[0]), .B(
        i_cmd[0]), .C(n4), .ZN(n6) );
  MOAI22D1BWP30P140LVT U15 ( .A1(n11), .A2(n6), .B1(i_data_bus[0]), .B2(n5), 
        .ZN(N287) );
  INVD1BWP30P140LVT U16 ( .I(i_data_bus[33]), .ZN(n12) );
  MOAI22D1BWP30P140LVT U17 ( .A1(n6), .A2(n12), .B1(n5), .B2(i_data_bus[1]), 
        .ZN(N288) );
  INVD1BWP30P140LVT U18 ( .I(i_data_bus[34]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U19 ( .A1(n6), .A2(n13), .B1(n5), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140LVT U20 ( .I(i_data_bus[35]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U21 ( .A1(n6), .A2(n14), .B1(n5), .B2(i_data_bus[3]), 
        .ZN(N290) );
  INVD1BWP30P140LVT U22 ( .I(i_data_bus[36]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U23 ( .A1(n6), .A2(n15), .B1(n5), .B2(i_data_bus[4]), 
        .ZN(N291) );
  INVD1BWP30P140LVT U24 ( .I(i_data_bus[37]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U25 ( .A1(n6), .A2(n16), .B1(n5), .B2(i_data_bus[5]), 
        .ZN(N292) );
  INVD1BWP30P140LVT U26 ( .I(i_data_bus[38]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U27 ( .A1(n6), .A2(n17), .B1(n5), .B2(i_data_bus[6]), 
        .ZN(N293) );
  INVD1BWP30P140LVT U28 ( .I(i_data_bus[39]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U29 ( .A1(n6), .A2(n18), .B1(n5), .B2(i_data_bus[7]), 
        .ZN(N294) );
  INVD1BWP30P140LVT U30 ( .I(i_data_bus[40]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U31 ( .A1(n6), .A2(n19), .B1(n5), .B2(i_data_bus[8]), 
        .ZN(N295) );
  INVD1BWP30P140LVT U32 ( .I(i_data_bus[41]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U33 ( .A1(n6), .A2(n20), .B1(n5), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140LVT U34 ( .I(i_data_bus[42]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U35 ( .A1(n6), .A2(n21), .B1(n5), .B2(i_data_bus[10]), 
        .ZN(N297) );
  INVD1BWP30P140LVT U36 ( .I(i_data_bus[43]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U37 ( .A1(n6), .A2(n22), .B1(n5), .B2(i_data_bus[11]), 
        .ZN(N298) );
  INVD1BWP30P140LVT U38 ( .I(i_data_bus[44]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U39 ( .A1(n6), .A2(n23), .B1(n5), .B2(i_data_bus[12]), 
        .ZN(N299) );
  INVD1BWP30P140LVT U40 ( .I(i_data_bus[45]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U41 ( .A1(n6), .A2(n24), .B1(n5), .B2(i_data_bus[13]), 
        .ZN(N300) );
  INVD1BWP30P140LVT U42 ( .I(i_data_bus[46]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U43 ( .A1(n6), .A2(n25), .B1(n5), .B2(i_data_bus[14]), 
        .ZN(N301) );
  INVD1BWP30P140LVT U44 ( .I(i_data_bus[47]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U45 ( .A1(n6), .A2(n26), .B1(n5), .B2(i_data_bus[15]), 
        .ZN(N302) );
  INVD1BWP30P140LVT U46 ( .I(i_data_bus[48]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U47 ( .A1(n6), .A2(n27), .B1(n5), .B2(i_data_bus[16]), 
        .ZN(N303) );
  INVD1BWP30P140LVT U48 ( .I(i_data_bus[49]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U49 ( .A1(n6), .A2(n28), .B1(n5), .B2(i_data_bus[17]), 
        .ZN(N304) );
  INVD1BWP30P140LVT U50 ( .I(i_data_bus[50]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U51 ( .A1(n6), .A2(n29), .B1(n5), .B2(i_data_bus[18]), 
        .ZN(N305) );
  INVD1BWP30P140LVT U52 ( .I(i_data_bus[51]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U53 ( .A1(n6), .A2(n30), .B1(n5), .B2(i_data_bus[19]), 
        .ZN(N306) );
  INVD1BWP30P140LVT U54 ( .I(i_data_bus[52]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U55 ( .A1(n6), .A2(n31), .B1(n5), .B2(i_data_bus[20]), 
        .ZN(N307) );
  INVD1BWP30P140LVT U56 ( .I(i_data_bus[53]), .ZN(n32) );
  MOAI22D1BWP30P140LVT U57 ( .A1(n6), .A2(n32), .B1(n5), .B2(i_data_bus[21]), 
        .ZN(N308) );
  INVD1BWP30P140LVT U58 ( .I(i_data_bus[54]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U59 ( .A1(n6), .A2(n33), .B1(n5), .B2(i_data_bus[22]), 
        .ZN(N309) );
  INVD1BWP30P140LVT U60 ( .I(i_data_bus[55]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U61 ( .A1(n6), .A2(n34), .B1(n5), .B2(i_data_bus[23]), 
        .ZN(N310) );
  INVD1BWP30P140LVT U62 ( .I(i_data_bus[56]), .ZN(n35) );
  MOAI22D1BWP30P140LVT U63 ( .A1(n6), .A2(n35), .B1(n5), .B2(i_data_bus[24]), 
        .ZN(N311) );
  INVD1BWP30P140LVT U64 ( .I(i_data_bus[57]), .ZN(n36) );
  MOAI22D1BWP30P140LVT U65 ( .A1(n6), .A2(n36), .B1(n5), .B2(i_data_bus[25]), 
        .ZN(N312) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[58]), .ZN(n37) );
  MOAI22D1BWP30P140LVT U67 ( .A1(n6), .A2(n37), .B1(n5), .B2(i_data_bus[26]), 
        .ZN(N313) );
  INVD1BWP30P140LVT U68 ( .I(i_data_bus[59]), .ZN(n38) );
  MOAI22D1BWP30P140LVT U69 ( .A1(n6), .A2(n38), .B1(n5), .B2(i_data_bus[27]), 
        .ZN(N314) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[60]), .ZN(n39) );
  MOAI22D1BWP30P140LVT U71 ( .A1(n6), .A2(n39), .B1(n5), .B2(i_data_bus[28]), 
        .ZN(N315) );
  INVD1BWP30P140LVT U72 ( .I(i_data_bus[61]), .ZN(n40) );
  MOAI22D1BWP30P140LVT U73 ( .A1(n6), .A2(n40), .B1(n5), .B2(i_data_bus[29]), 
        .ZN(N316) );
  INVD1BWP30P140LVT U74 ( .I(i_data_bus[62]), .ZN(n41) );
  MOAI22D1BWP30P140LVT U75 ( .A1(n6), .A2(n41), .B1(n5), .B2(i_data_bus[30]), 
        .ZN(N317) );
  INVD1BWP30P140LVT U76 ( .I(i_data_bus[63]), .ZN(n44) );
  MOAI22D1BWP30P140LVT U77 ( .A1(n6), .A2(n44), .B1(n5), .B2(i_data_bus[31]), 
        .ZN(N318) );
  OAI21D1BWP30P140LVT U78 ( .A1(i_cmd[0]), .A2(i_valid[0]), .B(n7), .ZN(n8) );
  AO211D1BWP30P140LVT U79 ( .A1(i_cmd[0]), .A2(n9), .B(i_cmd[1]), .C(n8), .Z(
        n10) );
  INVD2BWP30P140LVT U80 ( .I(n10), .ZN(n42) );
  MOAI22D1BWP30P140LVT U81 ( .A1(n11), .A2(n43), .B1(i_data_bus[0]), .B2(n42), 
        .ZN(N319) );
  MOAI22D1BWP30P140LVT U82 ( .A1(n12), .A2(n43), .B1(i_data_bus[1]), .B2(n42), 
        .ZN(N320) );
  MOAI22D1BWP30P140LVT U83 ( .A1(n13), .A2(n43), .B1(i_data_bus[2]), .B2(n42), 
        .ZN(N321) );
  MOAI22D1BWP30P140LVT U84 ( .A1(n14), .A2(n43), .B1(i_data_bus[3]), .B2(n42), 
        .ZN(N322) );
  MOAI22D1BWP30P140LVT U85 ( .A1(n15), .A2(n43), .B1(i_data_bus[4]), .B2(n42), 
        .ZN(N323) );
  MOAI22D1BWP30P140LVT U86 ( .A1(n16), .A2(n43), .B1(i_data_bus[5]), .B2(n42), 
        .ZN(N324) );
  MOAI22D1BWP30P140LVT U87 ( .A1(n17), .A2(n43), .B1(i_data_bus[6]), .B2(n42), 
        .ZN(N325) );
  MOAI22D1BWP30P140LVT U88 ( .A1(n18), .A2(n43), .B1(i_data_bus[7]), .B2(n42), 
        .ZN(N326) );
  MOAI22D1BWP30P140LVT U89 ( .A1(n19), .A2(n43), .B1(i_data_bus[8]), .B2(n42), 
        .ZN(N327) );
  MOAI22D1BWP30P140LVT U90 ( .A1(n20), .A2(n43), .B1(i_data_bus[9]), .B2(n42), 
        .ZN(N328) );
  MOAI22D1BWP30P140LVT U91 ( .A1(n21), .A2(n43), .B1(i_data_bus[10]), .B2(n42), 
        .ZN(N329) );
  MOAI22D1BWP30P140LVT U92 ( .A1(n22), .A2(n43), .B1(i_data_bus[11]), .B2(n42), 
        .ZN(N330) );
  MOAI22D1BWP30P140LVT U93 ( .A1(n23), .A2(n43), .B1(i_data_bus[12]), .B2(n42), 
        .ZN(N331) );
  MOAI22D1BWP30P140LVT U94 ( .A1(n24), .A2(n43), .B1(i_data_bus[13]), .B2(n42), 
        .ZN(N332) );
  MOAI22D1BWP30P140LVT U95 ( .A1(n25), .A2(n43), .B1(i_data_bus[14]), .B2(n42), 
        .ZN(N333) );
  MOAI22D1BWP30P140LVT U96 ( .A1(n26), .A2(n43), .B1(i_data_bus[15]), .B2(n42), 
        .ZN(N334) );
  MOAI22D1BWP30P140LVT U97 ( .A1(n27), .A2(n43), .B1(i_data_bus[16]), .B2(n42), 
        .ZN(N335) );
  MOAI22D1BWP30P140LVT U98 ( .A1(n28), .A2(n43), .B1(i_data_bus[17]), .B2(n42), 
        .ZN(N336) );
  MOAI22D1BWP30P140LVT U99 ( .A1(n29), .A2(n43), .B1(i_data_bus[18]), .B2(n42), 
        .ZN(N337) );
  MOAI22D1BWP30P140LVT U100 ( .A1(n30), .A2(n43), .B1(i_data_bus[19]), .B2(n42), .ZN(N338) );
  MOAI22D1BWP30P140LVT U101 ( .A1(n31), .A2(n43), .B1(i_data_bus[20]), .B2(n42), .ZN(N339) );
  MOAI22D1BWP30P140LVT U102 ( .A1(n32), .A2(n43), .B1(i_data_bus[21]), .B2(n42), .ZN(N340) );
  MOAI22D1BWP30P140LVT U103 ( .A1(n33), .A2(n43), .B1(i_data_bus[22]), .B2(n42), .ZN(N341) );
  MOAI22D1BWP30P140LVT U104 ( .A1(n34), .A2(n43), .B1(i_data_bus[23]), .B2(n42), .ZN(N342) );
  MOAI22D1BWP30P140LVT U105 ( .A1(n35), .A2(n43), .B1(i_data_bus[24]), .B2(n42), .ZN(N343) );
  MOAI22D1BWP30P140LVT U106 ( .A1(n36), .A2(n43), .B1(i_data_bus[25]), .B2(n42), .ZN(N344) );
  MOAI22D1BWP30P140LVT U107 ( .A1(n37), .A2(n43), .B1(i_data_bus[26]), .B2(n42), .ZN(N345) );
  MOAI22D1BWP30P140LVT U108 ( .A1(n38), .A2(n43), .B1(i_data_bus[27]), .B2(n42), .ZN(N346) );
  MOAI22D1BWP30P140LVT U109 ( .A1(n39), .A2(n43), .B1(i_data_bus[28]), .B2(n42), .ZN(N347) );
  MOAI22D1BWP30P140LVT U110 ( .A1(n40), .A2(n43), .B1(i_data_bus[29]), .B2(n42), .ZN(N348) );
  MOAI22D1BWP30P140LVT U111 ( .A1(n41), .A2(n43), .B1(i_data_bus[30]), .B2(n42), .ZN(N349) );
  MOAI22D1BWP30P140LVT U112 ( .A1(n44), .A2(n43), .B1(i_data_bus[31]), .B2(n42), .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_4 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1])
         );
  DFQD1BWP30P140LVT o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0])
         );
  INVD1BWP30P140LVT U3 ( .I(i_valid[1]), .ZN(n9) );
  INR2D1BWP30P140LVT U4 ( .A1(i_en), .B1(rst), .ZN(n7) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(n7), .A2(i_valid[0]), .ZN(n2) );
  NR2D2BWP30P140LVT U6 ( .A1(i_cmd[0]), .A2(n2), .ZN(n5) );
  AOI31D1BWP30P140LVT U7 ( .A1(i_cmd[0]), .A2(n7), .A3(i_valid[1]), .B(n5), 
        .ZN(n1) );
  INVD1BWP30P140LVT U8 ( .I(n1), .ZN(N353) );
  ND3D2BWP30P140LVT U9 ( .A1(n7), .A2(i_cmd[1]), .A3(i_valid[1]), .ZN(n43) );
  OAI21D1BWP30P140LVT U10 ( .A1(i_cmd[1]), .A2(n2), .B(n43), .ZN(N354) );
  INVD1BWP30P140LVT U11 ( .I(i_data_bus[32]), .ZN(n11) );
  INVD1BWP30P140LVT U12 ( .I(n7), .ZN(n3) );
  AOI21D1BWP30P140LVT U13 ( .A1(i_cmd[1]), .A2(n9), .B(n3), .ZN(n4) );
  OAI211OPTREPBD2BWP30P140LVT U14 ( .A1(i_cmd[1]), .A2(i_valid[0]), .B(
        i_cmd[0]), .C(n4), .ZN(n6) );
  MOAI22D1BWP30P140LVT U15 ( .A1(n11), .A2(n6), .B1(i_data_bus[0]), .B2(n5), 
        .ZN(N287) );
  INVD1BWP30P140LVT U16 ( .I(i_data_bus[33]), .ZN(n12) );
  MOAI22D1BWP30P140LVT U17 ( .A1(n6), .A2(n12), .B1(n5), .B2(i_data_bus[1]), 
        .ZN(N288) );
  INVD1BWP30P140LVT U18 ( .I(i_data_bus[34]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U19 ( .A1(n6), .A2(n13), .B1(n5), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140LVT U20 ( .I(i_data_bus[35]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U21 ( .A1(n6), .A2(n14), .B1(n5), .B2(i_data_bus[3]), 
        .ZN(N290) );
  INVD1BWP30P140LVT U22 ( .I(i_data_bus[36]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U23 ( .A1(n6), .A2(n15), .B1(n5), .B2(i_data_bus[4]), 
        .ZN(N291) );
  INVD1BWP30P140LVT U24 ( .I(i_data_bus[37]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U25 ( .A1(n6), .A2(n16), .B1(n5), .B2(i_data_bus[5]), 
        .ZN(N292) );
  INVD1BWP30P140LVT U26 ( .I(i_data_bus[38]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U27 ( .A1(n6), .A2(n17), .B1(n5), .B2(i_data_bus[6]), 
        .ZN(N293) );
  INVD1BWP30P140LVT U28 ( .I(i_data_bus[39]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U29 ( .A1(n6), .A2(n18), .B1(n5), .B2(i_data_bus[7]), 
        .ZN(N294) );
  INVD1BWP30P140LVT U30 ( .I(i_data_bus[40]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U31 ( .A1(n6), .A2(n19), .B1(n5), .B2(i_data_bus[8]), 
        .ZN(N295) );
  INVD1BWP30P140LVT U32 ( .I(i_data_bus[41]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U33 ( .A1(n6), .A2(n20), .B1(n5), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140LVT U34 ( .I(i_data_bus[42]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U35 ( .A1(n6), .A2(n21), .B1(n5), .B2(i_data_bus[10]), 
        .ZN(N297) );
  INVD1BWP30P140LVT U36 ( .I(i_data_bus[43]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U37 ( .A1(n6), .A2(n22), .B1(n5), .B2(i_data_bus[11]), 
        .ZN(N298) );
  INVD1BWP30P140LVT U38 ( .I(i_data_bus[44]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U39 ( .A1(n6), .A2(n23), .B1(n5), .B2(i_data_bus[12]), 
        .ZN(N299) );
  INVD1BWP30P140LVT U40 ( .I(i_data_bus[45]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U41 ( .A1(n6), .A2(n24), .B1(n5), .B2(i_data_bus[13]), 
        .ZN(N300) );
  INVD1BWP30P140LVT U42 ( .I(i_data_bus[46]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U43 ( .A1(n6), .A2(n25), .B1(n5), .B2(i_data_bus[14]), 
        .ZN(N301) );
  INVD1BWP30P140LVT U44 ( .I(i_data_bus[47]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U45 ( .A1(n6), .A2(n26), .B1(n5), .B2(i_data_bus[15]), 
        .ZN(N302) );
  INVD1BWP30P140LVT U46 ( .I(i_data_bus[48]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U47 ( .A1(n6), .A2(n27), .B1(n5), .B2(i_data_bus[16]), 
        .ZN(N303) );
  INVD1BWP30P140LVT U48 ( .I(i_data_bus[49]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U49 ( .A1(n6), .A2(n28), .B1(n5), .B2(i_data_bus[17]), 
        .ZN(N304) );
  INVD1BWP30P140LVT U50 ( .I(i_data_bus[50]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U51 ( .A1(n6), .A2(n29), .B1(n5), .B2(i_data_bus[18]), 
        .ZN(N305) );
  INVD1BWP30P140LVT U52 ( .I(i_data_bus[51]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U53 ( .A1(n6), .A2(n30), .B1(n5), .B2(i_data_bus[19]), 
        .ZN(N306) );
  INVD1BWP30P140LVT U54 ( .I(i_data_bus[52]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U55 ( .A1(n6), .A2(n31), .B1(n5), .B2(i_data_bus[20]), 
        .ZN(N307) );
  INVD1BWP30P140LVT U56 ( .I(i_data_bus[53]), .ZN(n32) );
  MOAI22D1BWP30P140LVT U57 ( .A1(n6), .A2(n32), .B1(n5), .B2(i_data_bus[21]), 
        .ZN(N308) );
  INVD1BWP30P140LVT U58 ( .I(i_data_bus[54]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U59 ( .A1(n6), .A2(n33), .B1(n5), .B2(i_data_bus[22]), 
        .ZN(N309) );
  INVD1BWP30P140LVT U60 ( .I(i_data_bus[55]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U61 ( .A1(n6), .A2(n34), .B1(n5), .B2(i_data_bus[23]), 
        .ZN(N310) );
  INVD1BWP30P140LVT U62 ( .I(i_data_bus[56]), .ZN(n35) );
  MOAI22D1BWP30P140LVT U63 ( .A1(n6), .A2(n35), .B1(n5), .B2(i_data_bus[24]), 
        .ZN(N311) );
  INVD1BWP30P140LVT U64 ( .I(i_data_bus[57]), .ZN(n36) );
  MOAI22D1BWP30P140LVT U65 ( .A1(n6), .A2(n36), .B1(n5), .B2(i_data_bus[25]), 
        .ZN(N312) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[58]), .ZN(n37) );
  MOAI22D1BWP30P140LVT U67 ( .A1(n6), .A2(n37), .B1(n5), .B2(i_data_bus[26]), 
        .ZN(N313) );
  INVD1BWP30P140LVT U68 ( .I(i_data_bus[59]), .ZN(n38) );
  MOAI22D1BWP30P140LVT U69 ( .A1(n6), .A2(n38), .B1(n5), .B2(i_data_bus[27]), 
        .ZN(N314) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[60]), .ZN(n39) );
  MOAI22D1BWP30P140LVT U71 ( .A1(n6), .A2(n39), .B1(n5), .B2(i_data_bus[28]), 
        .ZN(N315) );
  INVD1BWP30P140LVT U72 ( .I(i_data_bus[61]), .ZN(n40) );
  MOAI22D1BWP30P140LVT U73 ( .A1(n6), .A2(n40), .B1(n5), .B2(i_data_bus[29]), 
        .ZN(N316) );
  INVD1BWP30P140LVT U74 ( .I(i_data_bus[62]), .ZN(n41) );
  MOAI22D1BWP30P140LVT U75 ( .A1(n6), .A2(n41), .B1(n5), .B2(i_data_bus[30]), 
        .ZN(N317) );
  INVD1BWP30P140LVT U76 ( .I(i_data_bus[63]), .ZN(n44) );
  MOAI22D1BWP30P140LVT U77 ( .A1(n6), .A2(n44), .B1(n5), .B2(i_data_bus[31]), 
        .ZN(N318) );
  OAI21D1BWP30P140LVT U78 ( .A1(i_cmd[0]), .A2(i_valid[0]), .B(n7), .ZN(n8) );
  AO211D1BWP30P140LVT U79 ( .A1(i_cmd[0]), .A2(n9), .B(i_cmd[1]), .C(n8), .Z(
        n10) );
  INVD2BWP30P140LVT U80 ( .I(n10), .ZN(n42) );
  MOAI22D1BWP30P140LVT U81 ( .A1(n11), .A2(n43), .B1(i_data_bus[0]), .B2(n42), 
        .ZN(N319) );
  MOAI22D1BWP30P140LVT U82 ( .A1(n12), .A2(n43), .B1(i_data_bus[1]), .B2(n42), 
        .ZN(N320) );
  MOAI22D1BWP30P140LVT U83 ( .A1(n13), .A2(n43), .B1(i_data_bus[2]), .B2(n42), 
        .ZN(N321) );
  MOAI22D1BWP30P140LVT U84 ( .A1(n14), .A2(n43), .B1(i_data_bus[3]), .B2(n42), 
        .ZN(N322) );
  MOAI22D1BWP30P140LVT U85 ( .A1(n15), .A2(n43), .B1(i_data_bus[4]), .B2(n42), 
        .ZN(N323) );
  MOAI22D1BWP30P140LVT U86 ( .A1(n16), .A2(n43), .B1(i_data_bus[5]), .B2(n42), 
        .ZN(N324) );
  MOAI22D1BWP30P140LVT U87 ( .A1(n17), .A2(n43), .B1(i_data_bus[6]), .B2(n42), 
        .ZN(N325) );
  MOAI22D1BWP30P140LVT U88 ( .A1(n18), .A2(n43), .B1(i_data_bus[7]), .B2(n42), 
        .ZN(N326) );
  MOAI22D1BWP30P140LVT U89 ( .A1(n19), .A2(n43), .B1(i_data_bus[8]), .B2(n42), 
        .ZN(N327) );
  MOAI22D1BWP30P140LVT U90 ( .A1(n20), .A2(n43), .B1(i_data_bus[9]), .B2(n42), 
        .ZN(N328) );
  MOAI22D1BWP30P140LVT U91 ( .A1(n21), .A2(n43), .B1(i_data_bus[10]), .B2(n42), 
        .ZN(N329) );
  MOAI22D1BWP30P140LVT U92 ( .A1(n22), .A2(n43), .B1(i_data_bus[11]), .B2(n42), 
        .ZN(N330) );
  MOAI22D1BWP30P140LVT U93 ( .A1(n23), .A2(n43), .B1(i_data_bus[12]), .B2(n42), 
        .ZN(N331) );
  MOAI22D1BWP30P140LVT U94 ( .A1(n24), .A2(n43), .B1(i_data_bus[13]), .B2(n42), 
        .ZN(N332) );
  MOAI22D1BWP30P140LVT U95 ( .A1(n25), .A2(n43), .B1(i_data_bus[14]), .B2(n42), 
        .ZN(N333) );
  MOAI22D1BWP30P140LVT U96 ( .A1(n26), .A2(n43), .B1(i_data_bus[15]), .B2(n42), 
        .ZN(N334) );
  MOAI22D1BWP30P140LVT U97 ( .A1(n27), .A2(n43), .B1(i_data_bus[16]), .B2(n42), 
        .ZN(N335) );
  MOAI22D1BWP30P140LVT U98 ( .A1(n28), .A2(n43), .B1(i_data_bus[17]), .B2(n42), 
        .ZN(N336) );
  MOAI22D1BWP30P140LVT U99 ( .A1(n29), .A2(n43), .B1(i_data_bus[18]), .B2(n42), 
        .ZN(N337) );
  MOAI22D1BWP30P140LVT U100 ( .A1(n30), .A2(n43), .B1(i_data_bus[19]), .B2(n42), .ZN(N338) );
  MOAI22D1BWP30P140LVT U101 ( .A1(n31), .A2(n43), .B1(i_data_bus[20]), .B2(n42), .ZN(N339) );
  MOAI22D1BWP30P140LVT U102 ( .A1(n32), .A2(n43), .B1(i_data_bus[21]), .B2(n42), .ZN(N340) );
  MOAI22D1BWP30P140LVT U103 ( .A1(n33), .A2(n43), .B1(i_data_bus[22]), .B2(n42), .ZN(N341) );
  MOAI22D1BWP30P140LVT U104 ( .A1(n34), .A2(n43), .B1(i_data_bus[23]), .B2(n42), .ZN(N342) );
  MOAI22D1BWP30P140LVT U105 ( .A1(n35), .A2(n43), .B1(i_data_bus[24]), .B2(n42), .ZN(N343) );
  MOAI22D1BWP30P140LVT U106 ( .A1(n36), .A2(n43), .B1(i_data_bus[25]), .B2(n42), .ZN(N344) );
  MOAI22D1BWP30P140LVT U107 ( .A1(n37), .A2(n43), .B1(i_data_bus[26]), .B2(n42), .ZN(N345) );
  MOAI22D1BWP30P140LVT U108 ( .A1(n38), .A2(n43), .B1(i_data_bus[27]), .B2(n42), .ZN(N346) );
  MOAI22D1BWP30P140LVT U109 ( .A1(n39), .A2(n43), .B1(i_data_bus[28]), .B2(n42), .ZN(N347) );
  MOAI22D1BWP30P140LVT U110 ( .A1(n40), .A2(n43), .B1(i_data_bus[29]), .B2(n42), .ZN(N348) );
  MOAI22D1BWP30P140LVT U111 ( .A1(n41), .A2(n43), .B1(i_data_bus[30]), .B2(n42), .ZN(N349) );
  MOAI22D1BWP30P140LVT U112 ( .A1(n44), .A2(n43), .B1(i_data_bus[31]), .B2(n42), .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_5 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0])
         );
  DFQD1BWP30P140LVT o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1])
         );
  INVD1BWP30P140LVT U3 ( .I(i_valid[1]), .ZN(n9) );
  INR2D1BWP30P140LVT U4 ( .A1(i_en), .B1(rst), .ZN(n7) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(n7), .A2(i_valid[0]), .ZN(n2) );
  NR2D2BWP30P140LVT U6 ( .A1(i_cmd[0]), .A2(n2), .ZN(n5) );
  AOI31D1BWP30P140LVT U7 ( .A1(i_cmd[0]), .A2(n7), .A3(i_valid[1]), .B(n5), 
        .ZN(n1) );
  INVD1BWP30P140LVT U8 ( .I(n1), .ZN(N353) );
  ND3D2BWP30P140LVT U9 ( .A1(n7), .A2(i_cmd[1]), .A3(i_valid[1]), .ZN(n43) );
  OAI21D1BWP30P140LVT U10 ( .A1(i_cmd[1]), .A2(n2), .B(n43), .ZN(N354) );
  INVD1BWP30P140LVT U11 ( .I(i_data_bus[32]), .ZN(n11) );
  INVD1BWP30P140LVT U12 ( .I(n7), .ZN(n3) );
  AOI21D1BWP30P140LVT U13 ( .A1(i_cmd[1]), .A2(n9), .B(n3), .ZN(n4) );
  OAI211OPTREPBD2BWP30P140LVT U14 ( .A1(i_cmd[1]), .A2(i_valid[0]), .B(
        i_cmd[0]), .C(n4), .ZN(n6) );
  MOAI22D1BWP30P140LVT U15 ( .A1(n11), .A2(n6), .B1(i_data_bus[0]), .B2(n5), 
        .ZN(N287) );
  INVD1BWP30P140LVT U16 ( .I(i_data_bus[33]), .ZN(n12) );
  MOAI22D1BWP30P140LVT U17 ( .A1(n6), .A2(n12), .B1(n5), .B2(i_data_bus[1]), 
        .ZN(N288) );
  INVD1BWP30P140LVT U18 ( .I(i_data_bus[34]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U19 ( .A1(n6), .A2(n13), .B1(n5), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140LVT U20 ( .I(i_data_bus[35]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U21 ( .A1(n6), .A2(n14), .B1(n5), .B2(i_data_bus[3]), 
        .ZN(N290) );
  INVD1BWP30P140LVT U22 ( .I(i_data_bus[36]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U23 ( .A1(n6), .A2(n15), .B1(n5), .B2(i_data_bus[4]), 
        .ZN(N291) );
  INVD1BWP30P140LVT U24 ( .I(i_data_bus[37]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U25 ( .A1(n6), .A2(n16), .B1(n5), .B2(i_data_bus[5]), 
        .ZN(N292) );
  INVD1BWP30P140LVT U26 ( .I(i_data_bus[38]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U27 ( .A1(n6), .A2(n17), .B1(n5), .B2(i_data_bus[6]), 
        .ZN(N293) );
  INVD1BWP30P140LVT U28 ( .I(i_data_bus[39]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U29 ( .A1(n6), .A2(n18), .B1(n5), .B2(i_data_bus[7]), 
        .ZN(N294) );
  INVD1BWP30P140LVT U30 ( .I(i_data_bus[40]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U31 ( .A1(n6), .A2(n19), .B1(n5), .B2(i_data_bus[8]), 
        .ZN(N295) );
  INVD1BWP30P140LVT U32 ( .I(i_data_bus[41]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U33 ( .A1(n6), .A2(n20), .B1(n5), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140LVT U34 ( .I(i_data_bus[42]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U35 ( .A1(n6), .A2(n21), .B1(n5), .B2(i_data_bus[10]), 
        .ZN(N297) );
  INVD1BWP30P140LVT U36 ( .I(i_data_bus[43]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U37 ( .A1(n6), .A2(n22), .B1(n5), .B2(i_data_bus[11]), 
        .ZN(N298) );
  INVD1BWP30P140LVT U38 ( .I(i_data_bus[44]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U39 ( .A1(n6), .A2(n23), .B1(n5), .B2(i_data_bus[12]), 
        .ZN(N299) );
  INVD1BWP30P140LVT U40 ( .I(i_data_bus[45]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U41 ( .A1(n6), .A2(n24), .B1(n5), .B2(i_data_bus[13]), 
        .ZN(N300) );
  INVD1BWP30P140LVT U42 ( .I(i_data_bus[46]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U43 ( .A1(n6), .A2(n25), .B1(n5), .B2(i_data_bus[14]), 
        .ZN(N301) );
  INVD1BWP30P140LVT U44 ( .I(i_data_bus[47]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U45 ( .A1(n6), .A2(n26), .B1(n5), .B2(i_data_bus[15]), 
        .ZN(N302) );
  INVD1BWP30P140LVT U46 ( .I(i_data_bus[48]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U47 ( .A1(n6), .A2(n27), .B1(n5), .B2(i_data_bus[16]), 
        .ZN(N303) );
  INVD1BWP30P140LVT U48 ( .I(i_data_bus[49]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U49 ( .A1(n6), .A2(n28), .B1(n5), .B2(i_data_bus[17]), 
        .ZN(N304) );
  INVD1BWP30P140LVT U50 ( .I(i_data_bus[50]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U51 ( .A1(n6), .A2(n29), .B1(n5), .B2(i_data_bus[18]), 
        .ZN(N305) );
  INVD1BWP30P140LVT U52 ( .I(i_data_bus[51]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U53 ( .A1(n6), .A2(n30), .B1(n5), .B2(i_data_bus[19]), 
        .ZN(N306) );
  INVD1BWP30P140LVT U54 ( .I(i_data_bus[52]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U55 ( .A1(n6), .A2(n31), .B1(n5), .B2(i_data_bus[20]), 
        .ZN(N307) );
  INVD1BWP30P140LVT U56 ( .I(i_data_bus[53]), .ZN(n32) );
  MOAI22D1BWP30P140LVT U57 ( .A1(n6), .A2(n32), .B1(n5), .B2(i_data_bus[21]), 
        .ZN(N308) );
  INVD1BWP30P140LVT U58 ( .I(i_data_bus[54]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U59 ( .A1(n6), .A2(n33), .B1(n5), .B2(i_data_bus[22]), 
        .ZN(N309) );
  INVD1BWP30P140LVT U60 ( .I(i_data_bus[55]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U61 ( .A1(n6), .A2(n34), .B1(n5), .B2(i_data_bus[23]), 
        .ZN(N310) );
  INVD1BWP30P140LVT U62 ( .I(i_data_bus[56]), .ZN(n35) );
  MOAI22D1BWP30P140LVT U63 ( .A1(n6), .A2(n35), .B1(n5), .B2(i_data_bus[24]), 
        .ZN(N311) );
  INVD1BWP30P140LVT U64 ( .I(i_data_bus[57]), .ZN(n36) );
  MOAI22D1BWP30P140LVT U65 ( .A1(n6), .A2(n36), .B1(n5), .B2(i_data_bus[25]), 
        .ZN(N312) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[58]), .ZN(n37) );
  MOAI22D1BWP30P140LVT U67 ( .A1(n6), .A2(n37), .B1(n5), .B2(i_data_bus[26]), 
        .ZN(N313) );
  INVD1BWP30P140LVT U68 ( .I(i_data_bus[59]), .ZN(n38) );
  MOAI22D1BWP30P140LVT U69 ( .A1(n6), .A2(n38), .B1(n5), .B2(i_data_bus[27]), 
        .ZN(N314) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[60]), .ZN(n39) );
  MOAI22D1BWP30P140LVT U71 ( .A1(n6), .A2(n39), .B1(n5), .B2(i_data_bus[28]), 
        .ZN(N315) );
  INVD1BWP30P140LVT U72 ( .I(i_data_bus[61]), .ZN(n40) );
  MOAI22D1BWP30P140LVT U73 ( .A1(n6), .A2(n40), .B1(n5), .B2(i_data_bus[29]), 
        .ZN(N316) );
  INVD1BWP30P140LVT U74 ( .I(i_data_bus[62]), .ZN(n41) );
  MOAI22D1BWP30P140LVT U75 ( .A1(n6), .A2(n41), .B1(n5), .B2(i_data_bus[30]), 
        .ZN(N317) );
  INVD1BWP30P140LVT U76 ( .I(i_data_bus[63]), .ZN(n44) );
  MOAI22D1BWP30P140LVT U77 ( .A1(n6), .A2(n44), .B1(n5), .B2(i_data_bus[31]), 
        .ZN(N318) );
  OAI21D1BWP30P140LVT U78 ( .A1(i_cmd[0]), .A2(i_valid[0]), .B(n7), .ZN(n8) );
  AO211D1BWP30P140LVT U79 ( .A1(i_cmd[0]), .A2(n9), .B(i_cmd[1]), .C(n8), .Z(
        n10) );
  INVD2BWP30P140LVT U80 ( .I(n10), .ZN(n42) );
  MOAI22D1BWP30P140LVT U81 ( .A1(n11), .A2(n43), .B1(i_data_bus[0]), .B2(n42), 
        .ZN(N319) );
  MOAI22D1BWP30P140LVT U82 ( .A1(n12), .A2(n43), .B1(i_data_bus[1]), .B2(n42), 
        .ZN(N320) );
  MOAI22D1BWP30P140LVT U83 ( .A1(n13), .A2(n43), .B1(i_data_bus[2]), .B2(n42), 
        .ZN(N321) );
  MOAI22D1BWP30P140LVT U84 ( .A1(n14), .A2(n43), .B1(i_data_bus[3]), .B2(n42), 
        .ZN(N322) );
  MOAI22D1BWP30P140LVT U85 ( .A1(n15), .A2(n43), .B1(i_data_bus[4]), .B2(n42), 
        .ZN(N323) );
  MOAI22D1BWP30P140LVT U86 ( .A1(n16), .A2(n43), .B1(i_data_bus[5]), .B2(n42), 
        .ZN(N324) );
  MOAI22D1BWP30P140LVT U87 ( .A1(n17), .A2(n43), .B1(i_data_bus[6]), .B2(n42), 
        .ZN(N325) );
  MOAI22D1BWP30P140LVT U88 ( .A1(n18), .A2(n43), .B1(i_data_bus[7]), .B2(n42), 
        .ZN(N326) );
  MOAI22D1BWP30P140LVT U89 ( .A1(n19), .A2(n43), .B1(i_data_bus[8]), .B2(n42), 
        .ZN(N327) );
  MOAI22D1BWP30P140LVT U90 ( .A1(n20), .A2(n43), .B1(i_data_bus[9]), .B2(n42), 
        .ZN(N328) );
  MOAI22D1BWP30P140LVT U91 ( .A1(n21), .A2(n43), .B1(i_data_bus[10]), .B2(n42), 
        .ZN(N329) );
  MOAI22D1BWP30P140LVT U92 ( .A1(n22), .A2(n43), .B1(i_data_bus[11]), .B2(n42), 
        .ZN(N330) );
  MOAI22D1BWP30P140LVT U93 ( .A1(n23), .A2(n43), .B1(i_data_bus[12]), .B2(n42), 
        .ZN(N331) );
  MOAI22D1BWP30P140LVT U94 ( .A1(n24), .A2(n43), .B1(i_data_bus[13]), .B2(n42), 
        .ZN(N332) );
  MOAI22D1BWP30P140LVT U95 ( .A1(n25), .A2(n43), .B1(i_data_bus[14]), .B2(n42), 
        .ZN(N333) );
  MOAI22D1BWP30P140LVT U96 ( .A1(n26), .A2(n43), .B1(i_data_bus[15]), .B2(n42), 
        .ZN(N334) );
  MOAI22D1BWP30P140LVT U97 ( .A1(n27), .A2(n43), .B1(i_data_bus[16]), .B2(n42), 
        .ZN(N335) );
  MOAI22D1BWP30P140LVT U98 ( .A1(n28), .A2(n43), .B1(i_data_bus[17]), .B2(n42), 
        .ZN(N336) );
  MOAI22D1BWP30P140LVT U99 ( .A1(n29), .A2(n43), .B1(i_data_bus[18]), .B2(n42), 
        .ZN(N337) );
  MOAI22D1BWP30P140LVT U100 ( .A1(n30), .A2(n43), .B1(i_data_bus[19]), .B2(n42), .ZN(N338) );
  MOAI22D1BWP30P140LVT U101 ( .A1(n31), .A2(n43), .B1(i_data_bus[20]), .B2(n42), .ZN(N339) );
  MOAI22D1BWP30P140LVT U102 ( .A1(n32), .A2(n43), .B1(i_data_bus[21]), .B2(n42), .ZN(N340) );
  MOAI22D1BWP30P140LVT U103 ( .A1(n33), .A2(n43), .B1(i_data_bus[22]), .B2(n42), .ZN(N341) );
  MOAI22D1BWP30P140LVT U104 ( .A1(n34), .A2(n43), .B1(i_data_bus[23]), .B2(n42), .ZN(N342) );
  MOAI22D1BWP30P140LVT U105 ( .A1(n35), .A2(n43), .B1(i_data_bus[24]), .B2(n42), .ZN(N343) );
  MOAI22D1BWP30P140LVT U106 ( .A1(n36), .A2(n43), .B1(i_data_bus[25]), .B2(n42), .ZN(N344) );
  MOAI22D1BWP30P140LVT U107 ( .A1(n37), .A2(n43), .B1(i_data_bus[26]), .B2(n42), .ZN(N345) );
  MOAI22D1BWP30P140LVT U108 ( .A1(n38), .A2(n43), .B1(i_data_bus[27]), .B2(n42), .ZN(N346) );
  MOAI22D1BWP30P140LVT U109 ( .A1(n39), .A2(n43), .B1(i_data_bus[28]), .B2(n42), .ZN(N347) );
  MOAI22D1BWP30P140LVT U110 ( .A1(n40), .A2(n43), .B1(i_data_bus[29]), .B2(n42), .ZN(N348) );
  MOAI22D1BWP30P140LVT U111 ( .A1(n41), .A2(n43), .B1(i_data_bus[30]), .B2(n42), .ZN(N349) );
  MOAI22D1BWP30P140LVT U112 ( .A1(n44), .A2(n43), .B1(i_data_bus[31]), .B2(n42), .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_6 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1])
         );
  DFQD1BWP30P140LVT o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0])
         );
  INVD1BWP30P140LVT U3 ( .I(i_valid[1]), .ZN(n9) );
  INR2D1BWP30P140LVT U4 ( .A1(i_en), .B1(rst), .ZN(n7) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(n7), .A2(i_valid[0]), .ZN(n2) );
  NR2D2BWP30P140LVT U6 ( .A1(i_cmd[0]), .A2(n2), .ZN(n5) );
  AOI31D1BWP30P140LVT U7 ( .A1(i_cmd[0]), .A2(n7), .A3(i_valid[1]), .B(n5), 
        .ZN(n1) );
  INVD1BWP30P140LVT U8 ( .I(n1), .ZN(N353) );
  ND3D2BWP30P140LVT U9 ( .A1(n7), .A2(i_cmd[1]), .A3(i_valid[1]), .ZN(n43) );
  OAI21D1BWP30P140LVT U10 ( .A1(i_cmd[1]), .A2(n2), .B(n43), .ZN(N354) );
  INVD1BWP30P140LVT U11 ( .I(i_data_bus[32]), .ZN(n11) );
  INVD1BWP30P140LVT U12 ( .I(n7), .ZN(n3) );
  AOI21D1BWP30P140LVT U13 ( .A1(i_cmd[1]), .A2(n9), .B(n3), .ZN(n4) );
  OAI211OPTREPBD2BWP30P140LVT U14 ( .A1(i_cmd[1]), .A2(i_valid[0]), .B(
        i_cmd[0]), .C(n4), .ZN(n6) );
  MOAI22D1BWP30P140LVT U15 ( .A1(n11), .A2(n6), .B1(i_data_bus[0]), .B2(n5), 
        .ZN(N287) );
  INVD1BWP30P140LVT U16 ( .I(i_data_bus[33]), .ZN(n12) );
  MOAI22D1BWP30P140LVT U17 ( .A1(n6), .A2(n12), .B1(n5), .B2(i_data_bus[1]), 
        .ZN(N288) );
  INVD1BWP30P140LVT U18 ( .I(i_data_bus[34]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U19 ( .A1(n6), .A2(n13), .B1(n5), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140LVT U20 ( .I(i_data_bus[35]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U21 ( .A1(n6), .A2(n14), .B1(n5), .B2(i_data_bus[3]), 
        .ZN(N290) );
  INVD1BWP30P140LVT U22 ( .I(i_data_bus[36]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U23 ( .A1(n6), .A2(n15), .B1(n5), .B2(i_data_bus[4]), 
        .ZN(N291) );
  INVD1BWP30P140LVT U24 ( .I(i_data_bus[37]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U25 ( .A1(n6), .A2(n16), .B1(n5), .B2(i_data_bus[5]), 
        .ZN(N292) );
  INVD1BWP30P140LVT U26 ( .I(i_data_bus[38]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U27 ( .A1(n6), .A2(n17), .B1(n5), .B2(i_data_bus[6]), 
        .ZN(N293) );
  INVD1BWP30P140LVT U28 ( .I(i_data_bus[39]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U29 ( .A1(n6), .A2(n18), .B1(n5), .B2(i_data_bus[7]), 
        .ZN(N294) );
  INVD1BWP30P140LVT U30 ( .I(i_data_bus[40]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U31 ( .A1(n6), .A2(n19), .B1(n5), .B2(i_data_bus[8]), 
        .ZN(N295) );
  INVD1BWP30P140LVT U32 ( .I(i_data_bus[41]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U33 ( .A1(n6), .A2(n20), .B1(n5), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140LVT U34 ( .I(i_data_bus[42]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U35 ( .A1(n6), .A2(n21), .B1(n5), .B2(i_data_bus[10]), 
        .ZN(N297) );
  INVD1BWP30P140LVT U36 ( .I(i_data_bus[43]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U37 ( .A1(n6), .A2(n22), .B1(n5), .B2(i_data_bus[11]), 
        .ZN(N298) );
  INVD1BWP30P140LVT U38 ( .I(i_data_bus[44]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U39 ( .A1(n6), .A2(n23), .B1(n5), .B2(i_data_bus[12]), 
        .ZN(N299) );
  INVD1BWP30P140LVT U40 ( .I(i_data_bus[45]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U41 ( .A1(n6), .A2(n24), .B1(n5), .B2(i_data_bus[13]), 
        .ZN(N300) );
  INVD1BWP30P140LVT U42 ( .I(i_data_bus[46]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U43 ( .A1(n6), .A2(n25), .B1(n5), .B2(i_data_bus[14]), 
        .ZN(N301) );
  INVD1BWP30P140LVT U44 ( .I(i_data_bus[47]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U45 ( .A1(n6), .A2(n26), .B1(n5), .B2(i_data_bus[15]), 
        .ZN(N302) );
  INVD1BWP30P140LVT U46 ( .I(i_data_bus[48]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U47 ( .A1(n6), .A2(n27), .B1(n5), .B2(i_data_bus[16]), 
        .ZN(N303) );
  INVD1BWP30P140LVT U48 ( .I(i_data_bus[49]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U49 ( .A1(n6), .A2(n28), .B1(n5), .B2(i_data_bus[17]), 
        .ZN(N304) );
  INVD1BWP30P140LVT U50 ( .I(i_data_bus[50]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U51 ( .A1(n6), .A2(n29), .B1(n5), .B2(i_data_bus[18]), 
        .ZN(N305) );
  INVD1BWP30P140LVT U52 ( .I(i_data_bus[51]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U53 ( .A1(n6), .A2(n30), .B1(n5), .B2(i_data_bus[19]), 
        .ZN(N306) );
  INVD1BWP30P140LVT U54 ( .I(i_data_bus[52]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U55 ( .A1(n6), .A2(n31), .B1(n5), .B2(i_data_bus[20]), 
        .ZN(N307) );
  INVD1BWP30P140LVT U56 ( .I(i_data_bus[53]), .ZN(n32) );
  MOAI22D1BWP30P140LVT U57 ( .A1(n6), .A2(n32), .B1(n5), .B2(i_data_bus[21]), 
        .ZN(N308) );
  INVD1BWP30P140LVT U58 ( .I(i_data_bus[54]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U59 ( .A1(n6), .A2(n33), .B1(n5), .B2(i_data_bus[22]), 
        .ZN(N309) );
  INVD1BWP30P140LVT U60 ( .I(i_data_bus[55]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U61 ( .A1(n6), .A2(n34), .B1(n5), .B2(i_data_bus[23]), 
        .ZN(N310) );
  INVD1BWP30P140LVT U62 ( .I(i_data_bus[56]), .ZN(n35) );
  MOAI22D1BWP30P140LVT U63 ( .A1(n6), .A2(n35), .B1(n5), .B2(i_data_bus[24]), 
        .ZN(N311) );
  INVD1BWP30P140LVT U64 ( .I(i_data_bus[57]), .ZN(n36) );
  MOAI22D1BWP30P140LVT U65 ( .A1(n6), .A2(n36), .B1(n5), .B2(i_data_bus[25]), 
        .ZN(N312) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[58]), .ZN(n37) );
  MOAI22D1BWP30P140LVT U67 ( .A1(n6), .A2(n37), .B1(n5), .B2(i_data_bus[26]), 
        .ZN(N313) );
  INVD1BWP30P140LVT U68 ( .I(i_data_bus[59]), .ZN(n38) );
  MOAI22D1BWP30P140LVT U69 ( .A1(n6), .A2(n38), .B1(n5), .B2(i_data_bus[27]), 
        .ZN(N314) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[60]), .ZN(n39) );
  MOAI22D1BWP30P140LVT U71 ( .A1(n6), .A2(n39), .B1(n5), .B2(i_data_bus[28]), 
        .ZN(N315) );
  INVD1BWP30P140LVT U72 ( .I(i_data_bus[61]), .ZN(n40) );
  MOAI22D1BWP30P140LVT U73 ( .A1(n6), .A2(n40), .B1(n5), .B2(i_data_bus[29]), 
        .ZN(N316) );
  INVD1BWP30P140LVT U74 ( .I(i_data_bus[62]), .ZN(n41) );
  MOAI22D1BWP30P140LVT U75 ( .A1(n6), .A2(n41), .B1(n5), .B2(i_data_bus[30]), 
        .ZN(N317) );
  INVD1BWP30P140LVT U76 ( .I(i_data_bus[63]), .ZN(n44) );
  MOAI22D1BWP30P140LVT U77 ( .A1(n6), .A2(n44), .B1(n5), .B2(i_data_bus[31]), 
        .ZN(N318) );
  OAI21D1BWP30P140LVT U78 ( .A1(i_cmd[0]), .A2(i_valid[0]), .B(n7), .ZN(n8) );
  AO211D1BWP30P140LVT U79 ( .A1(i_cmd[0]), .A2(n9), .B(i_cmd[1]), .C(n8), .Z(
        n10) );
  INVD2BWP30P140LVT U80 ( .I(n10), .ZN(n42) );
  MOAI22D1BWP30P140LVT U81 ( .A1(n11), .A2(n43), .B1(i_data_bus[0]), .B2(n42), 
        .ZN(N319) );
  MOAI22D1BWP30P140LVT U82 ( .A1(n12), .A2(n43), .B1(i_data_bus[1]), .B2(n42), 
        .ZN(N320) );
  MOAI22D1BWP30P140LVT U83 ( .A1(n13), .A2(n43), .B1(i_data_bus[2]), .B2(n42), 
        .ZN(N321) );
  MOAI22D1BWP30P140LVT U84 ( .A1(n14), .A2(n43), .B1(i_data_bus[3]), .B2(n42), 
        .ZN(N322) );
  MOAI22D1BWP30P140LVT U85 ( .A1(n15), .A2(n43), .B1(i_data_bus[4]), .B2(n42), 
        .ZN(N323) );
  MOAI22D1BWP30P140LVT U86 ( .A1(n16), .A2(n43), .B1(i_data_bus[5]), .B2(n42), 
        .ZN(N324) );
  MOAI22D1BWP30P140LVT U87 ( .A1(n17), .A2(n43), .B1(i_data_bus[6]), .B2(n42), 
        .ZN(N325) );
  MOAI22D1BWP30P140LVT U88 ( .A1(n18), .A2(n43), .B1(i_data_bus[7]), .B2(n42), 
        .ZN(N326) );
  MOAI22D1BWP30P140LVT U89 ( .A1(n19), .A2(n43), .B1(i_data_bus[8]), .B2(n42), 
        .ZN(N327) );
  MOAI22D1BWP30P140LVT U90 ( .A1(n20), .A2(n43), .B1(i_data_bus[9]), .B2(n42), 
        .ZN(N328) );
  MOAI22D1BWP30P140LVT U91 ( .A1(n21), .A2(n43), .B1(i_data_bus[10]), .B2(n42), 
        .ZN(N329) );
  MOAI22D1BWP30P140LVT U92 ( .A1(n22), .A2(n43), .B1(i_data_bus[11]), .B2(n42), 
        .ZN(N330) );
  MOAI22D1BWP30P140LVT U93 ( .A1(n23), .A2(n43), .B1(i_data_bus[12]), .B2(n42), 
        .ZN(N331) );
  MOAI22D1BWP30P140LVT U94 ( .A1(n24), .A2(n43), .B1(i_data_bus[13]), .B2(n42), 
        .ZN(N332) );
  MOAI22D1BWP30P140LVT U95 ( .A1(n25), .A2(n43), .B1(i_data_bus[14]), .B2(n42), 
        .ZN(N333) );
  MOAI22D1BWP30P140LVT U96 ( .A1(n26), .A2(n43), .B1(i_data_bus[15]), .B2(n42), 
        .ZN(N334) );
  MOAI22D1BWP30P140LVT U97 ( .A1(n27), .A2(n43), .B1(i_data_bus[16]), .B2(n42), 
        .ZN(N335) );
  MOAI22D1BWP30P140LVT U98 ( .A1(n28), .A2(n43), .B1(i_data_bus[17]), .B2(n42), 
        .ZN(N336) );
  MOAI22D1BWP30P140LVT U99 ( .A1(n29), .A2(n43), .B1(i_data_bus[18]), .B2(n42), 
        .ZN(N337) );
  MOAI22D1BWP30P140LVT U100 ( .A1(n30), .A2(n43), .B1(i_data_bus[19]), .B2(n42), .ZN(N338) );
  MOAI22D1BWP30P140LVT U101 ( .A1(n31), .A2(n43), .B1(i_data_bus[20]), .B2(n42), .ZN(N339) );
  MOAI22D1BWP30P140LVT U102 ( .A1(n32), .A2(n43), .B1(i_data_bus[21]), .B2(n42), .ZN(N340) );
  MOAI22D1BWP30P140LVT U103 ( .A1(n33), .A2(n43), .B1(i_data_bus[22]), .B2(n42), .ZN(N341) );
  MOAI22D1BWP30P140LVT U104 ( .A1(n34), .A2(n43), .B1(i_data_bus[23]), .B2(n42), .ZN(N342) );
  MOAI22D1BWP30P140LVT U105 ( .A1(n35), .A2(n43), .B1(i_data_bus[24]), .B2(n42), .ZN(N343) );
  MOAI22D1BWP30P140LVT U106 ( .A1(n36), .A2(n43), .B1(i_data_bus[25]), .B2(n42), .ZN(N344) );
  MOAI22D1BWP30P140LVT U107 ( .A1(n37), .A2(n43), .B1(i_data_bus[26]), .B2(n42), .ZN(N345) );
  MOAI22D1BWP30P140LVT U108 ( .A1(n38), .A2(n43), .B1(i_data_bus[27]), .B2(n42), .ZN(N346) );
  MOAI22D1BWP30P140LVT U109 ( .A1(n39), .A2(n43), .B1(i_data_bus[28]), .B2(n42), .ZN(N347) );
  MOAI22D1BWP30P140LVT U110 ( .A1(n40), .A2(n43), .B1(i_data_bus[29]), .B2(n42), .ZN(N348) );
  MOAI22D1BWP30P140LVT U111 ( .A1(n41), .A2(n43), .B1(i_data_bus[30]), .B2(n42), .ZN(N349) );
  MOAI22D1BWP30P140LVT U112 ( .A1(n44), .A2(n43), .B1(i_data_bus[31]), .B2(n42), .ZN(N350) );
endmodule


module distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_7 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_en;
  wire   N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N353, N354, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_63_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_62_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_61_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_60_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_59_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_58_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_57_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_56_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_55_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_54_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_53_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_52_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_51_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_50_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_49_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_48_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_47_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_46_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_45_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_44_ ( .D(N331), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_43_ ( .D(N330), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_42_ ( .D(N329), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_41_ ( .D(N328), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_40_ ( .D(N327), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_39_ ( .D(N326), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_38_ ( .D(N325), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_37_ ( .D(N324), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_36_ ( .D(N323), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_35_ ( .D(N322), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_34_ ( .D(N321), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_33_ ( .D(N320), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_32_ ( .D(N319), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N318), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N317), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N316), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N315), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N314), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N313), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N312), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N311), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N310), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N309), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N308), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N307), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N306), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N305), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N304), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N303), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N302), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N301), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N300), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N299), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N298), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg_1_ ( .D(N354), .CP(clk), .Q(o_valid[1])
         );
  DFQD1BWP30P140LVT o_valid_inner_reg_0_ ( .D(N353), .CP(clk), .Q(o_valid[0])
         );
  INVD1BWP30P140LVT U3 ( .I(i_valid[1]), .ZN(n9) );
  INR2D1BWP30P140LVT U4 ( .A1(i_en), .B1(rst), .ZN(n7) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(n7), .A2(i_valid[0]), .ZN(n2) );
  NR2D2BWP30P140LVT U6 ( .A1(i_cmd[0]), .A2(n2), .ZN(n5) );
  AOI31D1BWP30P140LVT U7 ( .A1(i_cmd[0]), .A2(n7), .A3(i_valid[1]), .B(n5), 
        .ZN(n1) );
  INVD1BWP30P140LVT U8 ( .I(n1), .ZN(N353) );
  ND3D2BWP30P140LVT U9 ( .A1(n7), .A2(i_cmd[1]), .A3(i_valid[1]), .ZN(n43) );
  OAI21D1BWP30P140LVT U10 ( .A1(i_cmd[1]), .A2(n2), .B(n43), .ZN(N354) );
  INVD1BWP30P140LVT U11 ( .I(i_data_bus[32]), .ZN(n11) );
  INVD1BWP30P140LVT U12 ( .I(n7), .ZN(n3) );
  AOI21D1BWP30P140LVT U13 ( .A1(i_cmd[1]), .A2(n9), .B(n3), .ZN(n4) );
  OAI211OPTREPBD2BWP30P140LVT U14 ( .A1(i_cmd[1]), .A2(i_valid[0]), .B(
        i_cmd[0]), .C(n4), .ZN(n6) );
  MOAI22D1BWP30P140LVT U15 ( .A1(n11), .A2(n6), .B1(i_data_bus[0]), .B2(n5), 
        .ZN(N287) );
  INVD1BWP30P140LVT U16 ( .I(i_data_bus[33]), .ZN(n12) );
  MOAI22D1BWP30P140LVT U17 ( .A1(n6), .A2(n12), .B1(n5), .B2(i_data_bus[1]), 
        .ZN(N288) );
  INVD1BWP30P140LVT U18 ( .I(i_data_bus[34]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U19 ( .A1(n6), .A2(n13), .B1(n5), .B2(i_data_bus[2]), 
        .ZN(N289) );
  INVD1BWP30P140LVT U20 ( .I(i_data_bus[35]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U21 ( .A1(n6), .A2(n14), .B1(n5), .B2(i_data_bus[3]), 
        .ZN(N290) );
  INVD1BWP30P140LVT U22 ( .I(i_data_bus[36]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U23 ( .A1(n6), .A2(n15), .B1(n5), .B2(i_data_bus[4]), 
        .ZN(N291) );
  INVD1BWP30P140LVT U24 ( .I(i_data_bus[37]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U25 ( .A1(n6), .A2(n16), .B1(n5), .B2(i_data_bus[5]), 
        .ZN(N292) );
  INVD1BWP30P140LVT U26 ( .I(i_data_bus[38]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U27 ( .A1(n6), .A2(n17), .B1(n5), .B2(i_data_bus[6]), 
        .ZN(N293) );
  INVD1BWP30P140LVT U28 ( .I(i_data_bus[39]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U29 ( .A1(n6), .A2(n18), .B1(n5), .B2(i_data_bus[7]), 
        .ZN(N294) );
  INVD1BWP30P140LVT U30 ( .I(i_data_bus[40]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U31 ( .A1(n6), .A2(n19), .B1(n5), .B2(i_data_bus[8]), 
        .ZN(N295) );
  INVD1BWP30P140LVT U32 ( .I(i_data_bus[41]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U33 ( .A1(n6), .A2(n20), .B1(n5), .B2(i_data_bus[9]), 
        .ZN(N296) );
  INVD1BWP30P140LVT U34 ( .I(i_data_bus[42]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U35 ( .A1(n6), .A2(n21), .B1(n5), .B2(i_data_bus[10]), 
        .ZN(N297) );
  INVD1BWP30P140LVT U36 ( .I(i_data_bus[43]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U37 ( .A1(n6), .A2(n22), .B1(n5), .B2(i_data_bus[11]), 
        .ZN(N298) );
  INVD1BWP30P140LVT U38 ( .I(i_data_bus[44]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U39 ( .A1(n6), .A2(n23), .B1(n5), .B2(i_data_bus[12]), 
        .ZN(N299) );
  INVD1BWP30P140LVT U40 ( .I(i_data_bus[45]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U41 ( .A1(n6), .A2(n24), .B1(n5), .B2(i_data_bus[13]), 
        .ZN(N300) );
  INVD1BWP30P140LVT U42 ( .I(i_data_bus[46]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U43 ( .A1(n6), .A2(n25), .B1(n5), .B2(i_data_bus[14]), 
        .ZN(N301) );
  INVD1BWP30P140LVT U44 ( .I(i_data_bus[47]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U45 ( .A1(n6), .A2(n26), .B1(n5), .B2(i_data_bus[15]), 
        .ZN(N302) );
  INVD1BWP30P140LVT U46 ( .I(i_data_bus[48]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U47 ( .A1(n6), .A2(n27), .B1(n5), .B2(i_data_bus[16]), 
        .ZN(N303) );
  INVD1BWP30P140LVT U48 ( .I(i_data_bus[49]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U49 ( .A1(n6), .A2(n28), .B1(n5), .B2(i_data_bus[17]), 
        .ZN(N304) );
  INVD1BWP30P140LVT U50 ( .I(i_data_bus[50]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U51 ( .A1(n6), .A2(n29), .B1(n5), .B2(i_data_bus[18]), 
        .ZN(N305) );
  INVD1BWP30P140LVT U52 ( .I(i_data_bus[51]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U53 ( .A1(n6), .A2(n30), .B1(n5), .B2(i_data_bus[19]), 
        .ZN(N306) );
  INVD1BWP30P140LVT U54 ( .I(i_data_bus[52]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U55 ( .A1(n6), .A2(n31), .B1(n5), .B2(i_data_bus[20]), 
        .ZN(N307) );
  INVD1BWP30P140LVT U56 ( .I(i_data_bus[53]), .ZN(n32) );
  MOAI22D1BWP30P140LVT U57 ( .A1(n6), .A2(n32), .B1(n5), .B2(i_data_bus[21]), 
        .ZN(N308) );
  INVD1BWP30P140LVT U58 ( .I(i_data_bus[54]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U59 ( .A1(n6), .A2(n33), .B1(n5), .B2(i_data_bus[22]), 
        .ZN(N309) );
  INVD1BWP30P140LVT U60 ( .I(i_data_bus[55]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U61 ( .A1(n6), .A2(n34), .B1(n5), .B2(i_data_bus[23]), 
        .ZN(N310) );
  INVD1BWP30P140LVT U62 ( .I(i_data_bus[56]), .ZN(n35) );
  MOAI22D1BWP30P140LVT U63 ( .A1(n6), .A2(n35), .B1(n5), .B2(i_data_bus[24]), 
        .ZN(N311) );
  INVD1BWP30P140LVT U64 ( .I(i_data_bus[57]), .ZN(n36) );
  MOAI22D1BWP30P140LVT U65 ( .A1(n6), .A2(n36), .B1(n5), .B2(i_data_bus[25]), 
        .ZN(N312) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[58]), .ZN(n37) );
  MOAI22D1BWP30P140LVT U67 ( .A1(n6), .A2(n37), .B1(n5), .B2(i_data_bus[26]), 
        .ZN(N313) );
  INVD1BWP30P140LVT U68 ( .I(i_data_bus[59]), .ZN(n38) );
  MOAI22D1BWP30P140LVT U69 ( .A1(n6), .A2(n38), .B1(n5), .B2(i_data_bus[27]), 
        .ZN(N314) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[60]), .ZN(n39) );
  MOAI22D1BWP30P140LVT U71 ( .A1(n6), .A2(n39), .B1(n5), .B2(i_data_bus[28]), 
        .ZN(N315) );
  INVD1BWP30P140LVT U72 ( .I(i_data_bus[61]), .ZN(n40) );
  MOAI22D1BWP30P140LVT U73 ( .A1(n6), .A2(n40), .B1(n5), .B2(i_data_bus[29]), 
        .ZN(N316) );
  INVD1BWP30P140LVT U74 ( .I(i_data_bus[62]), .ZN(n41) );
  MOAI22D1BWP30P140LVT U75 ( .A1(n6), .A2(n41), .B1(n5), .B2(i_data_bus[30]), 
        .ZN(N317) );
  INVD1BWP30P140LVT U76 ( .I(i_data_bus[63]), .ZN(n44) );
  MOAI22D1BWP30P140LVT U77 ( .A1(n6), .A2(n44), .B1(n5), .B2(i_data_bus[31]), 
        .ZN(N318) );
  OAI21D1BWP30P140LVT U78 ( .A1(i_cmd[0]), .A2(i_valid[0]), .B(n7), .ZN(n8) );
  AO211D1BWP30P140LVT U79 ( .A1(i_cmd[0]), .A2(n9), .B(i_cmd[1]), .C(n8), .Z(
        n10) );
  INVD2BWP30P140LVT U80 ( .I(n10), .ZN(n42) );
  MOAI22D1BWP30P140LVT U81 ( .A1(n11), .A2(n43), .B1(i_data_bus[0]), .B2(n42), 
        .ZN(N319) );
  MOAI22D1BWP30P140LVT U82 ( .A1(n12), .A2(n43), .B1(i_data_bus[1]), .B2(n42), 
        .ZN(N320) );
  MOAI22D1BWP30P140LVT U83 ( .A1(n13), .A2(n43), .B1(i_data_bus[2]), .B2(n42), 
        .ZN(N321) );
  MOAI22D1BWP30P140LVT U84 ( .A1(n14), .A2(n43), .B1(i_data_bus[3]), .B2(n42), 
        .ZN(N322) );
  MOAI22D1BWP30P140LVT U85 ( .A1(n15), .A2(n43), .B1(i_data_bus[4]), .B2(n42), 
        .ZN(N323) );
  MOAI22D1BWP30P140LVT U86 ( .A1(n16), .A2(n43), .B1(i_data_bus[5]), .B2(n42), 
        .ZN(N324) );
  MOAI22D1BWP30P140LVT U87 ( .A1(n17), .A2(n43), .B1(i_data_bus[6]), .B2(n42), 
        .ZN(N325) );
  MOAI22D1BWP30P140LVT U88 ( .A1(n18), .A2(n43), .B1(i_data_bus[7]), .B2(n42), 
        .ZN(N326) );
  MOAI22D1BWP30P140LVT U89 ( .A1(n19), .A2(n43), .B1(i_data_bus[8]), .B2(n42), 
        .ZN(N327) );
  MOAI22D1BWP30P140LVT U90 ( .A1(n20), .A2(n43), .B1(i_data_bus[9]), .B2(n42), 
        .ZN(N328) );
  MOAI22D1BWP30P140LVT U91 ( .A1(n21), .A2(n43), .B1(i_data_bus[10]), .B2(n42), 
        .ZN(N329) );
  MOAI22D1BWP30P140LVT U92 ( .A1(n22), .A2(n43), .B1(i_data_bus[11]), .B2(n42), 
        .ZN(N330) );
  MOAI22D1BWP30P140LVT U93 ( .A1(n23), .A2(n43), .B1(i_data_bus[12]), .B2(n42), 
        .ZN(N331) );
  MOAI22D1BWP30P140LVT U94 ( .A1(n24), .A2(n43), .B1(i_data_bus[13]), .B2(n42), 
        .ZN(N332) );
  MOAI22D1BWP30P140LVT U95 ( .A1(n25), .A2(n43), .B1(i_data_bus[14]), .B2(n42), 
        .ZN(N333) );
  MOAI22D1BWP30P140LVT U96 ( .A1(n26), .A2(n43), .B1(i_data_bus[15]), .B2(n42), 
        .ZN(N334) );
  MOAI22D1BWP30P140LVT U97 ( .A1(n27), .A2(n43), .B1(i_data_bus[16]), .B2(n42), 
        .ZN(N335) );
  MOAI22D1BWP30P140LVT U98 ( .A1(n28), .A2(n43), .B1(i_data_bus[17]), .B2(n42), 
        .ZN(N336) );
  MOAI22D1BWP30P140LVT U99 ( .A1(n29), .A2(n43), .B1(i_data_bus[18]), .B2(n42), 
        .ZN(N337) );
  MOAI22D1BWP30P140LVT U100 ( .A1(n30), .A2(n43), .B1(i_data_bus[19]), .B2(n42), .ZN(N338) );
  MOAI22D1BWP30P140LVT U101 ( .A1(n31), .A2(n43), .B1(i_data_bus[20]), .B2(n42), .ZN(N339) );
  MOAI22D1BWP30P140LVT U102 ( .A1(n32), .A2(n43), .B1(i_data_bus[21]), .B2(n42), .ZN(N340) );
  MOAI22D1BWP30P140LVT U103 ( .A1(n33), .A2(n43), .B1(i_data_bus[22]), .B2(n42), .ZN(N341) );
  MOAI22D1BWP30P140LVT U104 ( .A1(n34), .A2(n43), .B1(i_data_bus[23]), .B2(n42), .ZN(N342) );
  MOAI22D1BWP30P140LVT U105 ( .A1(n35), .A2(n43), .B1(i_data_bus[24]), .B2(n42), .ZN(N343) );
  MOAI22D1BWP30P140LVT U106 ( .A1(n36), .A2(n43), .B1(i_data_bus[25]), .B2(n42), .ZN(N344) );
  MOAI22D1BWP30P140LVT U107 ( .A1(n37), .A2(n43), .B1(i_data_bus[26]), .B2(n42), .ZN(N345) );
  MOAI22D1BWP30P140LVT U108 ( .A1(n38), .A2(n43), .B1(i_data_bus[27]), .B2(n42), .ZN(N346) );
  MOAI22D1BWP30P140LVT U109 ( .A1(n39), .A2(n43), .B1(i_data_bus[28]), .B2(n42), .ZN(N347) );
  MOAI22D1BWP30P140LVT U110 ( .A1(n40), .A2(n43), .B1(i_data_bus[29]), .B2(n42), .ZN(N348) );
  MOAI22D1BWP30P140LVT U111 ( .A1(n41), .A2(n43), .B1(i_data_bus[30]), .B2(n42), .ZN(N349) );
  MOAI22D1BWP30P140LVT U112 ( .A1(n44), .A2(n43), .B1(i_data_bus[31]), .B2(n42), .ZN(N350) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_1 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  INVD1BWP30P140LVT U3 ( .I(n6), .ZN(n7) );
  IND2D1BWP30P140LVT U4 ( .A1(n5), .B1(n4), .ZN(n6) );
  INVD1BWP30P140LVT U5 ( .I(n7), .ZN(n35) );
  ND2D1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n3) );
  INVD1BWP30P140LVT U7 ( .I(n7), .ZN(n40) );
  NR2D3BWP30P140LVT U8 ( .A1(n3), .A2(n2), .ZN(n1) );
  OR2D1BWP30P140LVT U9 ( .A1(rst), .A2(i_cmd[0]), .Z(n2) );
  ND3D1BWP30P140LVT U10 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n5)
         );
  INVD1BWP30P140LVT U11 ( .I(rst), .ZN(n4) );
  IND2D1BWP30P140LVT U12 ( .A1(n1), .B1(n40), .ZN(N91) );
  INVD1BWP30P140LVT U13 ( .I(i_data_bus[54]), .ZN(n8) );
  MOAI22D1BWP30P140LVT U14 ( .A1(n8), .A2(n35), .B1(i_data_bus[22]), .B2(n1), 
        .ZN(N114) );
  INVD1BWP30P140LVT U15 ( .I(i_data_bus[52]), .ZN(n9) );
  MOAI22D1BWP30P140LVT U16 ( .A1(n9), .A2(n35), .B1(i_data_bus[20]), .B2(n1), 
        .ZN(N112) );
  INVD1BWP30P140LVT U17 ( .I(i_data_bus[50]), .ZN(n10) );
  MOAI22D1BWP30P140LVT U18 ( .A1(n10), .A2(n35), .B1(i_data_bus[18]), .B2(n1), 
        .ZN(N110) );
  INVD1BWP30P140LVT U19 ( .I(i_data_bus[48]), .ZN(n11) );
  MOAI22D1BWP30P140LVT U20 ( .A1(n11), .A2(n35), .B1(i_data_bus[16]), .B2(n1), 
        .ZN(N108) );
  INVD1BWP30P140LVT U21 ( .I(i_data_bus[37]), .ZN(n12) );
  MOAI22D1BWP30P140LVT U22 ( .A1(n12), .A2(n40), .B1(i_data_bus[5]), .B2(n1), 
        .ZN(N97) );
  INVD1BWP30P140LVT U23 ( .I(i_data_bus[38]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U24 ( .A1(n13), .A2(n40), .B1(i_data_bus[6]), .B2(n1), 
        .ZN(N98) );
  INVD1BWP30P140LVT U25 ( .I(i_data_bus[39]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U26 ( .A1(n14), .A2(n40), .B1(i_data_bus[7]), .B2(n1), 
        .ZN(N99) );
  INVD1BWP30P140LVT U27 ( .I(i_data_bus[40]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U28 ( .A1(n15), .A2(n40), .B1(i_data_bus[8]), .B2(n1), 
        .ZN(N100) );
  INVD1BWP30P140LVT U29 ( .I(i_data_bus[41]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U30 ( .A1(n16), .A2(n40), .B1(i_data_bus[9]), .B2(n1), 
        .ZN(N101) );
  INVD1BWP30P140LVT U31 ( .I(i_data_bus[42]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U32 ( .A1(n17), .A2(n40), .B1(i_data_bus[10]), .B2(n1), 
        .ZN(N102) );
  INVD1BWP30P140LVT U33 ( .I(i_data_bus[43]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U34 ( .A1(n18), .A2(n40), .B1(i_data_bus[11]), .B2(n1), 
        .ZN(N103) );
  INVD1BWP30P140LVT U35 ( .I(i_data_bus[36]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U36 ( .A1(n19), .A2(n40), .B1(i_data_bus[4]), .B2(n1), 
        .ZN(N96) );
  INVD1BWP30P140LVT U37 ( .I(i_data_bus[35]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U38 ( .A1(n20), .A2(n40), .B1(i_data_bus[3]), .B2(n1), 
        .ZN(N95) );
  INVD1BWP30P140LVT U39 ( .I(i_data_bus[34]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U40 ( .A1(n21), .A2(n40), .B1(i_data_bus[2]), .B2(n1), 
        .ZN(N94) );
  INVD1BWP30P140LVT U41 ( .I(i_data_bus[33]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U42 ( .A1(n22), .A2(n40), .B1(i_data_bus[1]), .B2(n1), 
        .ZN(N93) );
  INVD1BWP30P140LVT U43 ( .I(i_data_bus[32]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U44 ( .A1(n23), .A2(n40), .B1(i_data_bus[0]), .B2(n1), 
        .ZN(N92) );
  INVD1BWP30P140LVT U45 ( .I(i_data_bus[57]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U46 ( .A1(n24), .A2(n35), .B1(i_data_bus[25]), .B2(n1), 
        .ZN(N117) );
  INVD1BWP30P140LVT U47 ( .I(i_data_bus[47]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U48 ( .A1(n25), .A2(n35), .B1(i_data_bus[15]), .B2(n1), 
        .ZN(N107) );
  INVD1BWP30P140LVT U49 ( .I(i_data_bus[44]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U50 ( .A1(n26), .A2(n35), .B1(i_data_bus[12]), .B2(n1), 
        .ZN(N104) );
  INVD1BWP30P140LVT U51 ( .I(i_data_bus[45]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U52 ( .A1(n27), .A2(n35), .B1(i_data_bus[13]), .B2(n1), 
        .ZN(N105) );
  INVD1BWP30P140LVT U53 ( .I(i_data_bus[46]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U54 ( .A1(n28), .A2(n35), .B1(i_data_bus[14]), .B2(n1), 
        .ZN(N106) );
  INVD1BWP30P140LVT U55 ( .I(i_data_bus[61]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U56 ( .A1(n29), .A2(n35), .B1(i_data_bus[29]), .B2(n1), 
        .ZN(N121) );
  INVD1BWP30P140LVT U57 ( .I(i_data_bus[59]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U58 ( .A1(n30), .A2(n35), .B1(i_data_bus[27]), .B2(n1), 
        .ZN(N119) );
  INVD1BWP30P140LVT U59 ( .I(i_data_bus[63]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U60 ( .A1(n31), .A2(n35), .B1(i_data_bus[31]), .B2(n1), 
        .ZN(N123) );
  INVD1BWP30P140LVT U61 ( .I(i_data_bus[55]), .ZN(n32) );
  MOAI22D1BWP30P140LVT U62 ( .A1(n32), .A2(n35), .B1(i_data_bus[23]), .B2(n1), 
        .ZN(N115) );
  INVD1BWP30P140LVT U63 ( .I(i_data_bus[49]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U64 ( .A1(n33), .A2(n35), .B1(i_data_bus[17]), .B2(n1), 
        .ZN(N109) );
  INVD1BWP30P140LVT U65 ( .I(i_data_bus[53]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U66 ( .A1(n34), .A2(n35), .B1(i_data_bus[21]), .B2(n1), 
        .ZN(N113) );
  INVD1BWP30P140LVT U67 ( .I(i_data_bus[51]), .ZN(n36) );
  MOAI22D1BWP30P140LVT U68 ( .A1(n36), .A2(n35), .B1(i_data_bus[19]), .B2(n1), 
        .ZN(N111) );
  INVD1BWP30P140LVT U69 ( .I(i_data_bus[56]), .ZN(n37) );
  MOAI22D1BWP30P140LVT U70 ( .A1(n37), .A2(n40), .B1(i_data_bus[24]), .B2(n1), 
        .ZN(N116) );
  INVD1BWP30P140LVT U71 ( .I(i_data_bus[58]), .ZN(n38) );
  MOAI22D1BWP30P140LVT U72 ( .A1(n38), .A2(n40), .B1(i_data_bus[26]), .B2(n1), 
        .ZN(N118) );
  INVD1BWP30P140LVT U73 ( .I(i_data_bus[60]), .ZN(n39) );
  MOAI22D1BWP30P140LVT U74 ( .A1(n39), .A2(n40), .B1(i_data_bus[28]), .B2(n1), 
        .ZN(N120) );
  INVD1BWP30P140LVT U75 ( .I(i_data_bus[62]), .ZN(n41) );
  MOAI22D1BWP30P140LVT U76 ( .A1(n41), .A2(n40), .B1(i_data_bus[30]), .B2(n1), 
        .ZN(N122) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_1 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_1 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_2 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  INVD1BWP30P140LVT U3 ( .I(n6), .ZN(n7) );
  IND2D1BWP30P140LVT U4 ( .A1(n5), .B1(n4), .ZN(n6) );
  INVD1BWP30P140LVT U5 ( .I(n7), .ZN(n35) );
  ND2D1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n3) );
  INVD1BWP30P140LVT U7 ( .I(n7), .ZN(n40) );
  NR2D3BWP30P140LVT U8 ( .A1(n3), .A2(n2), .ZN(n1) );
  OR2D1BWP30P140LVT U9 ( .A1(rst), .A2(i_cmd[0]), .Z(n2) );
  ND3D1BWP30P140LVT U10 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n5)
         );
  INVD1BWP30P140LVT U11 ( .I(rst), .ZN(n4) );
  IND2D1BWP30P140LVT U12 ( .A1(n1), .B1(n40), .ZN(N91) );
  INVD1BWP30P140LVT U13 ( .I(i_data_bus[54]), .ZN(n8) );
  MOAI22D1BWP30P140LVT U14 ( .A1(n8), .A2(n35), .B1(i_data_bus[22]), .B2(n1), 
        .ZN(N114) );
  INVD1BWP30P140LVT U15 ( .I(i_data_bus[50]), .ZN(n9) );
  MOAI22D1BWP30P140LVT U16 ( .A1(n9), .A2(n35), .B1(i_data_bus[18]), .B2(n1), 
        .ZN(N110) );
  INVD1BWP30P140LVT U17 ( .I(i_data_bus[52]), .ZN(n10) );
  MOAI22D1BWP30P140LVT U18 ( .A1(n10), .A2(n35), .B1(i_data_bus[20]), .B2(n1), 
        .ZN(N112) );
  INVD1BWP30P140LVT U19 ( .I(i_data_bus[48]), .ZN(n11) );
  MOAI22D1BWP30P140LVT U20 ( .A1(n11), .A2(n35), .B1(i_data_bus[16]), .B2(n1), 
        .ZN(N108) );
  INVD1BWP30P140LVT U21 ( .I(i_data_bus[37]), .ZN(n12) );
  MOAI22D1BWP30P140LVT U22 ( .A1(n12), .A2(n40), .B1(i_data_bus[5]), .B2(n1), 
        .ZN(N97) );
  INVD1BWP30P140LVT U23 ( .I(i_data_bus[33]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U24 ( .A1(n13), .A2(n40), .B1(i_data_bus[1]), .B2(n1), 
        .ZN(N93) );
  INVD1BWP30P140LVT U25 ( .I(i_data_bus[36]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U26 ( .A1(n14), .A2(n40), .B1(i_data_bus[4]), .B2(n1), 
        .ZN(N96) );
  INVD1BWP30P140LVT U27 ( .I(i_data_bus[35]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U28 ( .A1(n15), .A2(n40), .B1(i_data_bus[3]), .B2(n1), 
        .ZN(N95) );
  INVD1BWP30P140LVT U29 ( .I(i_data_bus[43]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U30 ( .A1(n16), .A2(n40), .B1(i_data_bus[11]), .B2(n1), 
        .ZN(N103) );
  INVD1BWP30P140LVT U31 ( .I(i_data_bus[39]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U32 ( .A1(n17), .A2(n40), .B1(i_data_bus[7]), .B2(n1), 
        .ZN(N99) );
  INVD1BWP30P140LVT U33 ( .I(i_data_bus[42]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U34 ( .A1(n18), .A2(n40), .B1(i_data_bus[10]), .B2(n1), 
        .ZN(N102) );
  INVD1BWP30P140LVT U35 ( .I(i_data_bus[41]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U36 ( .A1(n19), .A2(n40), .B1(i_data_bus[9]), .B2(n1), 
        .ZN(N101) );
  INVD1BWP30P140LVT U37 ( .I(i_data_bus[40]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U38 ( .A1(n20), .A2(n40), .B1(i_data_bus[8]), .B2(n1), 
        .ZN(N100) );
  INVD1BWP30P140LVT U39 ( .I(i_data_bus[38]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U40 ( .A1(n21), .A2(n40), .B1(i_data_bus[6]), .B2(n1), 
        .ZN(N98) );
  INVD1BWP30P140LVT U41 ( .I(i_data_bus[32]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U42 ( .A1(n22), .A2(n40), .B1(i_data_bus[0]), .B2(n1), 
        .ZN(N92) );
  INVD1BWP30P140LVT U43 ( .I(i_data_bus[34]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U44 ( .A1(n23), .A2(n40), .B1(i_data_bus[2]), .B2(n1), 
        .ZN(N94) );
  INVD1BWP30P140LVT U45 ( .I(i_data_bus[45]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U46 ( .A1(n24), .A2(n35), .B1(i_data_bus[13]), .B2(n1), 
        .ZN(N105) );
  INVD1BWP30P140LVT U47 ( .I(i_data_bus[47]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U48 ( .A1(n25), .A2(n35), .B1(i_data_bus[15]), .B2(n1), 
        .ZN(N107) );
  INVD1BWP30P140LVT U49 ( .I(i_data_bus[46]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U50 ( .A1(n26), .A2(n35), .B1(i_data_bus[14]), .B2(n1), 
        .ZN(N106) );
  INVD1BWP30P140LVT U51 ( .I(i_data_bus[55]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U52 ( .A1(n27), .A2(n35), .B1(i_data_bus[23]), .B2(n1), 
        .ZN(N115) );
  INVD1BWP30P140LVT U53 ( .I(i_data_bus[49]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U54 ( .A1(n28), .A2(n35), .B1(i_data_bus[17]), .B2(n1), 
        .ZN(N109) );
  INVD1BWP30P140LVT U55 ( .I(i_data_bus[59]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U56 ( .A1(n29), .A2(n35), .B1(i_data_bus[27]), .B2(n1), 
        .ZN(N119) );
  INVD1BWP30P140LVT U57 ( .I(i_data_bus[61]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U58 ( .A1(n30), .A2(n35), .B1(i_data_bus[29]), .B2(n1), 
        .ZN(N121) );
  INVD1BWP30P140LVT U59 ( .I(i_data_bus[63]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U60 ( .A1(n31), .A2(n35), .B1(i_data_bus[31]), .B2(n1), 
        .ZN(N123) );
  INVD1BWP30P140LVT U61 ( .I(i_data_bus[44]), .ZN(n32) );
  MOAI22D1BWP30P140LVT U62 ( .A1(n32), .A2(n35), .B1(i_data_bus[12]), .B2(n1), 
        .ZN(N104) );
  INVD1BWP30P140LVT U63 ( .I(i_data_bus[53]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U64 ( .A1(n33), .A2(n35), .B1(i_data_bus[21]), .B2(n1), 
        .ZN(N113) );
  INVD1BWP30P140LVT U65 ( .I(i_data_bus[57]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U66 ( .A1(n34), .A2(n35), .B1(i_data_bus[25]), .B2(n1), 
        .ZN(N117) );
  INVD1BWP30P140LVT U67 ( .I(i_data_bus[51]), .ZN(n36) );
  MOAI22D1BWP30P140LVT U68 ( .A1(n36), .A2(n35), .B1(i_data_bus[19]), .B2(n1), 
        .ZN(N111) );
  INVD1BWP30P140LVT U69 ( .I(i_data_bus[58]), .ZN(n37) );
  MOAI22D1BWP30P140LVT U70 ( .A1(n37), .A2(n40), .B1(i_data_bus[26]), .B2(n1), 
        .ZN(N118) );
  INVD1BWP30P140LVT U71 ( .I(i_data_bus[56]), .ZN(n38) );
  MOAI22D1BWP30P140LVT U72 ( .A1(n38), .A2(n40), .B1(i_data_bus[24]), .B2(n1), 
        .ZN(N116) );
  INVD1BWP30P140LVT U73 ( .I(i_data_bus[60]), .ZN(n39) );
  MOAI22D1BWP30P140LVT U74 ( .A1(n39), .A2(n40), .B1(i_data_bus[28]), .B2(n1), 
        .ZN(N120) );
  INVD1BWP30P140LVT U75 ( .I(i_data_bus[62]), .ZN(n41) );
  MOAI22D1BWP30P140LVT U76 ( .A1(n41), .A2(n40), .B1(i_data_bus[30]), .B2(n1), 
        .ZN(N122) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_2 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_2 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_3 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U36 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_3 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_3 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_4 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2D1BWP30P140LVT U3 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n2), .A2(rst), .ZN(n3) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_4 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_4 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_5 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_5 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_5 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_6 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_6 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_6 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_1 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_6 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_5 merge_i_data_low ( .clk(
        clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(i_en), 
        .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_4 o_fwd ( .clk(clk), .rst(
        rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), .o_valid(
        inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), 
        .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_3 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_2 o_data_high ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_1 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_7 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D3BWP30P140LVT U3 ( .A1(n3), .A2(n2), .ZN(n1) );
  INVD1BWP30P140LVT U4 ( .I(n6), .ZN(n7) );
  IND2D1BWP30P140LVT U5 ( .A1(n5), .B1(n4), .ZN(n6) );
  INVD1BWP30P140LVT U6 ( .I(n7), .ZN(n35) );
  ND2D1BWP30P140LVT U7 ( .A1(i_en), .A2(i_valid[0]), .ZN(n3) );
  INVD1BWP30P140LVT U8 ( .I(n7), .ZN(n40) );
  OR2D1BWP30P140LVT U9 ( .A1(rst), .A2(i_cmd[0]), .Z(n2) );
  ND3D1BWP30P140LVT U10 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n5)
         );
  INVD1BWP30P140LVT U11 ( .I(rst), .ZN(n4) );
  IND2D1BWP30P140LVT U12 ( .A1(n1), .B1(n40), .ZN(N91) );
  INVD1BWP30P140LVT U13 ( .I(i_data_bus[48]), .ZN(n8) );
  MOAI22D1BWP30P140LVT U14 ( .A1(n8), .A2(n35), .B1(i_data_bus[16]), .B2(n1), 
        .ZN(N108) );
  INVD1BWP30P140LVT U15 ( .I(i_data_bus[54]), .ZN(n9) );
  MOAI22D1BWP30P140LVT U16 ( .A1(n9), .A2(n35), .B1(i_data_bus[22]), .B2(n1), 
        .ZN(N114) );
  INVD1BWP30P140LVT U17 ( .I(i_data_bus[50]), .ZN(n10) );
  MOAI22D1BWP30P140LVT U18 ( .A1(n10), .A2(n35), .B1(i_data_bus[18]), .B2(n1), 
        .ZN(N110) );
  INVD1BWP30P140LVT U19 ( .I(i_data_bus[52]), .ZN(n11) );
  MOAI22D1BWP30P140LVT U20 ( .A1(n11), .A2(n35), .B1(i_data_bus[20]), .B2(n1), 
        .ZN(N112) );
  INVD1BWP30P140LVT U21 ( .I(i_data_bus[36]), .ZN(n12) );
  MOAI22D1BWP30P140LVT U22 ( .A1(n12), .A2(n40), .B1(i_data_bus[4]), .B2(n1), 
        .ZN(N96) );
  INVD1BWP30P140LVT U23 ( .I(i_data_bus[38]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U24 ( .A1(n13), .A2(n40), .B1(i_data_bus[6]), .B2(n1), 
        .ZN(N98) );
  INVD1BWP30P140LVT U25 ( .I(i_data_bus[39]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U26 ( .A1(n14), .A2(n40), .B1(i_data_bus[7]), .B2(n1), 
        .ZN(N99) );
  INVD1BWP30P140LVT U27 ( .I(i_data_bus[32]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U28 ( .A1(n15), .A2(n40), .B1(i_data_bus[0]), .B2(n1), 
        .ZN(N92) );
  INVD1BWP30P140LVT U29 ( .I(i_data_bus[37]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U30 ( .A1(n16), .A2(n40), .B1(i_data_bus[5]), .B2(n1), 
        .ZN(N97) );
  INVD1BWP30P140LVT U31 ( .I(i_data_bus[34]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U32 ( .A1(n17), .A2(n40), .B1(i_data_bus[2]), .B2(n1), 
        .ZN(N94) );
  INVD1BWP30P140LVT U33 ( .I(i_data_bus[35]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U34 ( .A1(n18), .A2(n40), .B1(i_data_bus[3]), .B2(n1), 
        .ZN(N95) );
  INVD1BWP30P140LVT U35 ( .I(i_data_bus[40]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U36 ( .A1(n19), .A2(n40), .B1(i_data_bus[8]), .B2(n1), 
        .ZN(N100) );
  INVD1BWP30P140LVT U37 ( .I(i_data_bus[41]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U38 ( .A1(n20), .A2(n40), .B1(i_data_bus[9]), .B2(n1), 
        .ZN(N101) );
  INVD1BWP30P140LVT U39 ( .I(i_data_bus[42]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U40 ( .A1(n21), .A2(n40), .B1(i_data_bus[10]), .B2(n1), 
        .ZN(N102) );
  INVD1BWP30P140LVT U41 ( .I(i_data_bus[43]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U42 ( .A1(n22), .A2(n40), .B1(i_data_bus[11]), .B2(n1), 
        .ZN(N103) );
  INVD1BWP30P140LVT U43 ( .I(i_data_bus[33]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U44 ( .A1(n23), .A2(n40), .B1(i_data_bus[1]), .B2(n1), 
        .ZN(N93) );
  INVD1BWP30P140LVT U45 ( .I(i_data_bus[61]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U46 ( .A1(n24), .A2(n35), .B1(i_data_bus[29]), .B2(n1), 
        .ZN(N121) );
  INVD1BWP30P140LVT U47 ( .I(i_data_bus[59]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U48 ( .A1(n25), .A2(n35), .B1(i_data_bus[27]), .B2(n1), 
        .ZN(N119) );
  INVD1BWP30P140LVT U49 ( .I(i_data_bus[53]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U50 ( .A1(n26), .A2(n35), .B1(i_data_bus[21]), .B2(n1), 
        .ZN(N113) );
  INVD1BWP30P140LVT U51 ( .I(i_data_bus[49]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U52 ( .A1(n27), .A2(n35), .B1(i_data_bus[17]), .B2(n1), 
        .ZN(N109) );
  INVD1BWP30P140LVT U53 ( .I(i_data_bus[63]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U54 ( .A1(n28), .A2(n35), .B1(i_data_bus[31]), .B2(n1), 
        .ZN(N123) );
  INVD1BWP30P140LVT U55 ( .I(i_data_bus[51]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U56 ( .A1(n29), .A2(n35), .B1(i_data_bus[19]), .B2(n1), 
        .ZN(N111) );
  INVD1BWP30P140LVT U57 ( .I(i_data_bus[47]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U58 ( .A1(n30), .A2(n35), .B1(i_data_bus[15]), .B2(n1), 
        .ZN(N107) );
  INVD1BWP30P140LVT U59 ( .I(i_data_bus[44]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U60 ( .A1(n31), .A2(n35), .B1(i_data_bus[12]), .B2(n1), 
        .ZN(N104) );
  INVD1BWP30P140LVT U61 ( .I(i_data_bus[45]), .ZN(n32) );
  MOAI22D1BWP30P140LVT U62 ( .A1(n32), .A2(n35), .B1(i_data_bus[13]), .B2(n1), 
        .ZN(N105) );
  INVD1BWP30P140LVT U63 ( .I(i_data_bus[46]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U64 ( .A1(n33), .A2(n35), .B1(i_data_bus[14]), .B2(n1), 
        .ZN(N106) );
  INVD1BWP30P140LVT U65 ( .I(i_data_bus[55]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U66 ( .A1(n34), .A2(n35), .B1(i_data_bus[23]), .B2(n1), 
        .ZN(N115) );
  INVD1BWP30P140LVT U67 ( .I(i_data_bus[57]), .ZN(n36) );
  MOAI22D1BWP30P140LVT U68 ( .A1(n36), .A2(n35), .B1(i_data_bus[25]), .B2(n1), 
        .ZN(N117) );
  INVD1BWP30P140LVT U69 ( .I(i_data_bus[58]), .ZN(n37) );
  MOAI22D1BWP30P140LVT U70 ( .A1(n37), .A2(n40), .B1(i_data_bus[26]), .B2(n1), 
        .ZN(N118) );
  INVD1BWP30P140LVT U71 ( .I(i_data_bus[62]), .ZN(n38) );
  MOAI22D1BWP30P140LVT U72 ( .A1(n38), .A2(n40), .B1(i_data_bus[30]), .B2(n1), 
        .ZN(N122) );
  INVD1BWP30P140LVT U73 ( .I(i_data_bus[56]), .ZN(n39) );
  MOAI22D1BWP30P140LVT U74 ( .A1(n39), .A2(n40), .B1(i_data_bus[24]), .B2(n1), 
        .ZN(N116) );
  INVD1BWP30P140LVT U75 ( .I(i_data_bus[60]), .ZN(n41) );
  MOAI22D1BWP30P140LVT U76 ( .A1(n41), .A2(n40), .B1(i_data_bus[28]), .B2(n1), 
        .ZN(N120) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_7 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_7 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_8 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  INVD1BWP30P140LVT U3 ( .I(n5), .ZN(n6) );
  IND2D1BWP30P140LVT U4 ( .A1(n4), .B1(n3), .ZN(n5) );
  INVD1BWP30P140LVT U5 ( .I(n6), .ZN(n35) );
  ND2D1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  INVD1BWP30P140LVT U7 ( .I(n6), .ZN(n41) );
  OR2D1BWP30P140LVT U8 ( .A1(rst), .A2(i_cmd[0]), .Z(n1) );
  OR2D1BWP30P140LVT U9 ( .A1(n2), .A2(n1), .Z(n7) );
  INVD2BWP30P140LVT U10 ( .I(n7), .ZN(n40) );
  ND3D1BWP30P140LVT U11 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n4)
         );
  INVD1BWP30P140LVT U12 ( .I(rst), .ZN(n3) );
  IND2D1BWP30P140LVT U13 ( .A1(n40), .B1(n41), .ZN(N91) );
  INVD1BWP30P140LVT U14 ( .I(i_data_bus[52]), .ZN(n8) );
  MOAI22D1BWP30P140LVT U15 ( .A1(n8), .A2(n35), .B1(i_data_bus[20]), .B2(n40), 
        .ZN(N112) );
  INVD1BWP30P140LVT U16 ( .I(i_data_bus[54]), .ZN(n9) );
  MOAI22D1BWP30P140LVT U17 ( .A1(n9), .A2(n35), .B1(i_data_bus[22]), .B2(n40), 
        .ZN(N114) );
  INVD1BWP30P140LVT U18 ( .I(i_data_bus[48]), .ZN(n10) );
  MOAI22D1BWP30P140LVT U19 ( .A1(n10), .A2(n35), .B1(i_data_bus[16]), .B2(n40), 
        .ZN(N108) );
  INVD1BWP30P140LVT U20 ( .I(i_data_bus[50]), .ZN(n11) );
  MOAI22D1BWP30P140LVT U21 ( .A1(n11), .A2(n35), .B1(i_data_bus[18]), .B2(n40), 
        .ZN(N110) );
  INVD1BWP30P140LVT U22 ( .I(i_data_bus[38]), .ZN(n12) );
  MOAI22D1BWP30P140LVT U23 ( .A1(n12), .A2(n41), .B1(i_data_bus[6]), .B2(n40), 
        .ZN(N98) );
  INVD1BWP30P140LVT U24 ( .I(i_data_bus[43]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U25 ( .A1(n13), .A2(n41), .B1(i_data_bus[11]), .B2(n40), 
        .ZN(N103) );
  INVD1BWP30P140LVT U26 ( .I(i_data_bus[36]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U27 ( .A1(n14), .A2(n41), .B1(i_data_bus[4]), .B2(n40), 
        .ZN(N96) );
  INVD1BWP30P140LVT U28 ( .I(i_data_bus[39]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U29 ( .A1(n15), .A2(n41), .B1(i_data_bus[7]), .B2(n40), 
        .ZN(N99) );
  INVD1BWP30P140LVT U30 ( .I(i_data_bus[40]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U31 ( .A1(n16), .A2(n41), .B1(i_data_bus[8]), .B2(n40), 
        .ZN(N100) );
  INVD1BWP30P140LVT U32 ( .I(i_data_bus[41]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U33 ( .A1(n17), .A2(n41), .B1(i_data_bus[9]), .B2(n40), 
        .ZN(N101) );
  INVD1BWP30P140LVT U34 ( .I(i_data_bus[42]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U35 ( .A1(n18), .A2(n41), .B1(i_data_bus[10]), .B2(n40), 
        .ZN(N102) );
  INVD1BWP30P140LVT U36 ( .I(i_data_bus[35]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U37 ( .A1(n19), .A2(n41), .B1(i_data_bus[3]), .B2(n40), 
        .ZN(N95) );
  INVD1BWP30P140LVT U38 ( .I(i_data_bus[37]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U39 ( .A1(n20), .A2(n41), .B1(i_data_bus[5]), .B2(n40), 
        .ZN(N97) );
  INVD1BWP30P140LVT U40 ( .I(i_data_bus[34]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U41 ( .A1(n21), .A2(n41), .B1(i_data_bus[2]), .B2(n40), 
        .ZN(N94) );
  INVD1BWP30P140LVT U42 ( .I(i_data_bus[33]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U43 ( .A1(n22), .A2(n41), .B1(i_data_bus[1]), .B2(n40), 
        .ZN(N93) );
  INVD1BWP30P140LVT U44 ( .I(i_data_bus[32]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U45 ( .A1(n23), .A2(n41), .B1(i_data_bus[0]), .B2(n40), 
        .ZN(N92) );
  INVD1BWP30P140LVT U46 ( .I(i_data_bus[45]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U47 ( .A1(n24), .A2(n35), .B1(i_data_bus[13]), .B2(n40), 
        .ZN(N105) );
  INVD1BWP30P140LVT U48 ( .I(i_data_bus[61]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U49 ( .A1(n25), .A2(n35), .B1(i_data_bus[29]), .B2(n40), 
        .ZN(N121) );
  INVD1BWP30P140LVT U50 ( .I(i_data_bus[63]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U51 ( .A1(n26), .A2(n35), .B1(i_data_bus[31]), .B2(n40), 
        .ZN(N123) );
  INVD1BWP30P140LVT U52 ( .I(i_data_bus[57]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U53 ( .A1(n27), .A2(n35), .B1(i_data_bus[25]), .B2(n40), 
        .ZN(N117) );
  INVD1BWP30P140LVT U54 ( .I(i_data_bus[55]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U55 ( .A1(n28), .A2(n35), .B1(i_data_bus[23]), .B2(n40), 
        .ZN(N115) );
  INVD1BWP30P140LVT U56 ( .I(i_data_bus[53]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U57 ( .A1(n29), .A2(n35), .B1(i_data_bus[21]), .B2(n40), 
        .ZN(N113) );
  INVD1BWP30P140LVT U58 ( .I(i_data_bus[51]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U59 ( .A1(n30), .A2(n35), .B1(i_data_bus[19]), .B2(n40), 
        .ZN(N111) );
  INVD1BWP30P140LVT U60 ( .I(i_data_bus[49]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U61 ( .A1(n31), .A2(n35), .B1(i_data_bus[17]), .B2(n40), 
        .ZN(N109) );
  INVD1BWP30P140LVT U62 ( .I(i_data_bus[47]), .ZN(n32) );
  MOAI22D1BWP30P140LVT U63 ( .A1(n32), .A2(n35), .B1(i_data_bus[15]), .B2(n40), 
        .ZN(N107) );
  INVD1BWP30P140LVT U64 ( .I(i_data_bus[46]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U65 ( .A1(n33), .A2(n35), .B1(i_data_bus[14]), .B2(n40), 
        .ZN(N106) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[59]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U67 ( .A1(n34), .A2(n35), .B1(i_data_bus[27]), .B2(n40), 
        .ZN(N119) );
  INVD1BWP30P140LVT U68 ( .I(i_data_bus[44]), .ZN(n36) );
  MOAI22D1BWP30P140LVT U69 ( .A1(n36), .A2(n35), .B1(i_data_bus[12]), .B2(n40), 
        .ZN(N104) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[58]), .ZN(n37) );
  MOAI22D1BWP30P140LVT U71 ( .A1(n37), .A2(n41), .B1(i_data_bus[26]), .B2(n40), 
        .ZN(N118) );
  INVD1BWP30P140LVT U72 ( .I(i_data_bus[56]), .ZN(n38) );
  MOAI22D1BWP30P140LVT U73 ( .A1(n38), .A2(n41), .B1(i_data_bus[24]), .B2(n40), 
        .ZN(N116) );
  INVD1BWP30P140LVT U74 ( .I(i_data_bus[62]), .ZN(n39) );
  MOAI22D1BWP30P140LVT U75 ( .A1(n39), .A2(n41), .B1(i_data_bus[30]), .B2(n40), 
        .ZN(N122) );
  INVD1BWP30P140LVT U76 ( .I(i_data_bus[60]), .ZN(n42) );
  MOAI22D1BWP30P140LVT U77 ( .A1(n42), .A2(n41), .B1(i_data_bus[28]), .B2(n40), 
        .ZN(N120) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_8 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_8 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_9 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(i_cmd[0]), .A2(n2), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2OPTIBD1BWP30P140LVT U24 ( .A1(i_valid[0]), .A2(n1), .ZN(n2) );
  INR2D1BWP30P140LVT U25 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U36 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U37 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_9 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_9 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_10 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2OPTIBD1BWP30P140LVT U3 ( .A1(i_en), .A2(i_valid[0]), .ZN(n3) );
  NR3D0P7BWP30P140LVT U4 ( .A1(n3), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n1) );
  NR2D1BWP30P140LVT U6 ( .A1(n1), .A2(rst), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n2), .Z(n5) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[0]), .B1(n5), .B2(
        i_data_bus[32]), .Z(N92) );
  NR3D1P5BWP30P140LVT U9 ( .A1(n3), .A2(i_cmd[0]), .A3(rst), .ZN(n6) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n5), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n5), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[3]), .B1(n5), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n5), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n5), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[6]), .B1(n5), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n5), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n5), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[9]), .B1(n5), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n5), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n5), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[12]), .B1(n5), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n5), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n5), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[15]), .B1(n5), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n5), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n5), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[18]), .B1(n5), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n5), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n5), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[21]), .B1(n5), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n5), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n5), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[24]), .B1(n5), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n5), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n5), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[27]), .B1(n5), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n5), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n5), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n4), .A2(i_data_bus[30]), .B1(n5), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n5), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n5), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_10 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_10 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_11 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2OPTPAD1BWP30P140LVT U3 ( .A1(i_cmd[0]), .A2(n2), .ZN(n6) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_valid[0]), .A2(n1), .ZN(n2) );
  INR2D1BWP30P140LVT U5 ( .A1(i_en), .B1(rst), .ZN(n1) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  NR2D1BWP30P140LVT U7 ( .A1(n3), .A2(rst), .ZN(n4) );
  BUFFD2BWP30P140LVT U8 ( .I(n4), .Z(n5) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n5), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n5), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n5), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n5), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n5), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n5), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n5), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n5), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n5), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n5), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n5), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n5), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n5), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n5), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n5), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n5), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n5), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n5), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n5), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n5), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n5), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n5), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n5), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n5), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n5), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n5), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n5), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n5), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n5), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n5), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n5), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n5), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n5), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_11 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_11 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_12 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n3), .A2(rst), .A3(i_cmd[0]), .ZN(n68) );
  CKBD1BWP30P140LVT U4 ( .I(n2), .Z(n67) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n3) );
  ND2D1BWP30P140LVT U6 ( .A1(n54), .A2(n53), .ZN(N92) );
  ND2OPTIBD1BWP30P140LVT U7 ( .A1(n67), .A2(i_data_bus[32]), .ZN(n54) );
  ND2D1BWP30P140LVT U8 ( .A1(n68), .A2(i_data_bus[0]), .ZN(n53) );
  ND2D1BWP30P140LVT U9 ( .A1(n56), .A2(n55), .ZN(N93) );
  ND2OPTIBD1BWP30P140LVT U10 ( .A1(n67), .A2(i_data_bus[33]), .ZN(n56) );
  ND2D1BWP30P140LVT U11 ( .A1(n68), .A2(i_data_bus[1]), .ZN(n55) );
  ND2D1BWP30P140LVT U12 ( .A1(n58), .A2(n57), .ZN(N94) );
  ND2OPTIBD1BWP30P140LVT U13 ( .A1(n67), .A2(i_data_bus[34]), .ZN(n58) );
  ND2D1BWP30P140LVT U14 ( .A1(n68), .A2(i_data_bus[2]), .ZN(n57) );
  ND2D1BWP30P140LVT U15 ( .A1(n60), .A2(n59), .ZN(N95) );
  ND2OPTIBD1BWP30P140LVT U16 ( .A1(n67), .A2(i_data_bus[35]), .ZN(n60) );
  ND2D1BWP30P140LVT U17 ( .A1(n68), .A2(i_data_bus[3]), .ZN(n59) );
  ND2D1BWP30P140LVT U18 ( .A1(n62), .A2(n61), .ZN(N96) );
  ND2OPTIBD1BWP30P140LVT U19 ( .A1(n67), .A2(i_data_bus[36]), .ZN(n62) );
  ND2D1BWP30P140LVT U20 ( .A1(n68), .A2(i_data_bus[4]), .ZN(n61) );
  ND2D1BWP30P140LVT U21 ( .A1(n64), .A2(n63), .ZN(N97) );
  ND2OPTIBD1BWP30P140LVT U22 ( .A1(n67), .A2(i_data_bus[37]), .ZN(n64) );
  ND2D1BWP30P140LVT U23 ( .A1(n68), .A2(i_data_bus[5]), .ZN(n63) );
  ND2D1BWP30P140LVT U24 ( .A1(n66), .A2(n65), .ZN(N98) );
  ND2OPTIBD1BWP30P140LVT U25 ( .A1(n67), .A2(i_data_bus[38]), .ZN(n66) );
  ND2D1BWP30P140LVT U26 ( .A1(n68), .A2(i_data_bus[6]), .ZN(n65) );
  ND2D1BWP30P140LVT U27 ( .A1(n70), .A2(n69), .ZN(N99) );
  ND2OPTIBD1BWP30P140LVT U28 ( .A1(n67), .A2(i_data_bus[39]), .ZN(n70) );
  ND2D1BWP30P140LVT U29 ( .A1(n68), .A2(i_data_bus[7]), .ZN(n69) );
  ND2D1BWP30P140LVT U30 ( .A1(n5), .A2(n4), .ZN(N100) );
  ND2OPTIBD1BWP30P140LVT U31 ( .A1(n67), .A2(i_data_bus[40]), .ZN(n5) );
  ND2D1BWP30P140LVT U32 ( .A1(n68), .A2(i_data_bus[8]), .ZN(n4) );
  ND2D1BWP30P140LVT U33 ( .A1(n7), .A2(n6), .ZN(N101) );
  ND2OPTIBD1BWP30P140LVT U34 ( .A1(n67), .A2(i_data_bus[41]), .ZN(n7) );
  ND2D1BWP30P140LVT U35 ( .A1(n68), .A2(i_data_bus[9]), .ZN(n6) );
  ND2D1BWP30P140LVT U36 ( .A1(n9), .A2(n8), .ZN(N102) );
  ND2OPTIBD1BWP30P140LVT U37 ( .A1(n67), .A2(i_data_bus[42]), .ZN(n9) );
  ND2D1BWP30P140LVT U38 ( .A1(n68), .A2(i_data_bus[10]), .ZN(n8) );
  ND2D1BWP30P140LVT U39 ( .A1(n11), .A2(n10), .ZN(N103) );
  ND2OPTIBD1BWP30P140LVT U40 ( .A1(n67), .A2(i_data_bus[43]), .ZN(n11) );
  ND2D1BWP30P140LVT U41 ( .A1(n68), .A2(i_data_bus[11]), .ZN(n10) );
  ND2D1BWP30P140LVT U42 ( .A1(n13), .A2(n12), .ZN(N104) );
  ND2OPTIBD1BWP30P140LVT U43 ( .A1(n67), .A2(i_data_bus[44]), .ZN(n13) );
  ND2D1BWP30P140LVT U44 ( .A1(n68), .A2(i_data_bus[12]), .ZN(n12) );
  ND2D1BWP30P140LVT U45 ( .A1(n15), .A2(n14), .ZN(N105) );
  ND2OPTIBD1BWP30P140LVT U46 ( .A1(n67), .A2(i_data_bus[45]), .ZN(n15) );
  ND2D1BWP30P140LVT U47 ( .A1(n68), .A2(i_data_bus[13]), .ZN(n14) );
  ND2D1BWP30P140LVT U48 ( .A1(n17), .A2(n16), .ZN(N106) );
  ND2OPTIBD1BWP30P140LVT U49 ( .A1(n67), .A2(i_data_bus[46]), .ZN(n17) );
  ND2D1BWP30P140LVT U50 ( .A1(n68), .A2(i_data_bus[14]), .ZN(n16) );
  ND2D1BWP30P140LVT U51 ( .A1(n19), .A2(n18), .ZN(N107) );
  ND2OPTIBD1BWP30P140LVT U52 ( .A1(n67), .A2(i_data_bus[47]), .ZN(n19) );
  ND2D1BWP30P140LVT U53 ( .A1(n68), .A2(i_data_bus[15]), .ZN(n18) );
  ND2D1BWP30P140LVT U54 ( .A1(n21), .A2(n20), .ZN(N108) );
  ND2OPTIBD1BWP30P140LVT U55 ( .A1(n67), .A2(i_data_bus[48]), .ZN(n21) );
  ND2D1BWP30P140LVT U56 ( .A1(n68), .A2(i_data_bus[16]), .ZN(n20) );
  ND2D1BWP30P140LVT U57 ( .A1(n23), .A2(n22), .ZN(N109) );
  ND2OPTIBD1BWP30P140LVT U58 ( .A1(n67), .A2(i_data_bus[49]), .ZN(n23) );
  ND2D1BWP30P140LVT U59 ( .A1(n68), .A2(i_data_bus[17]), .ZN(n22) );
  ND2D1BWP30P140LVT U60 ( .A1(n25), .A2(n24), .ZN(N110) );
  ND2OPTIBD1BWP30P140LVT U61 ( .A1(n67), .A2(i_data_bus[50]), .ZN(n25) );
  ND2D1BWP30P140LVT U62 ( .A1(n68), .A2(i_data_bus[18]), .ZN(n24) );
  ND2D1BWP30P140LVT U63 ( .A1(n27), .A2(n26), .ZN(N111) );
  ND2OPTIBD1BWP30P140LVT U64 ( .A1(n67), .A2(i_data_bus[51]), .ZN(n27) );
  ND2D1BWP30P140LVT U65 ( .A1(n68), .A2(i_data_bus[19]), .ZN(n26) );
  ND2D1BWP30P140LVT U66 ( .A1(n29), .A2(n28), .ZN(N112) );
  ND2OPTIBD1BWP30P140LVT U67 ( .A1(n67), .A2(i_data_bus[52]), .ZN(n29) );
  ND2D1BWP30P140LVT U68 ( .A1(n68), .A2(i_data_bus[20]), .ZN(n28) );
  ND2D1BWP30P140LVT U69 ( .A1(n31), .A2(n30), .ZN(N113) );
  ND2OPTIBD1BWP30P140LVT U70 ( .A1(n67), .A2(i_data_bus[53]), .ZN(n31) );
  ND2D1BWP30P140LVT U71 ( .A1(n68), .A2(i_data_bus[21]), .ZN(n30) );
  ND2D1BWP30P140LVT U72 ( .A1(n33), .A2(n32), .ZN(N114) );
  ND2OPTIBD1BWP30P140LVT U73 ( .A1(n67), .A2(i_data_bus[54]), .ZN(n33) );
  ND2D1BWP30P140LVT U74 ( .A1(n68), .A2(i_data_bus[22]), .ZN(n32) );
  ND2D1BWP30P140LVT U75 ( .A1(n35), .A2(n34), .ZN(N115) );
  ND2OPTIBD1BWP30P140LVT U76 ( .A1(n67), .A2(i_data_bus[55]), .ZN(n35) );
  ND2D1BWP30P140LVT U77 ( .A1(n68), .A2(i_data_bus[23]), .ZN(n34) );
  ND2D1BWP30P140LVT U78 ( .A1(n37), .A2(n36), .ZN(N116) );
  ND2OPTIBD1BWP30P140LVT U79 ( .A1(n67), .A2(i_data_bus[56]), .ZN(n37) );
  ND2D1BWP30P140LVT U80 ( .A1(n68), .A2(i_data_bus[24]), .ZN(n36) );
  ND2D1BWP30P140LVT U81 ( .A1(n39), .A2(n38), .ZN(N117) );
  ND2OPTIBD1BWP30P140LVT U82 ( .A1(n67), .A2(i_data_bus[57]), .ZN(n39) );
  ND2D1BWP30P140LVT U83 ( .A1(n68), .A2(i_data_bus[25]), .ZN(n38) );
  ND2D1BWP30P140LVT U84 ( .A1(n41), .A2(n40), .ZN(N118) );
  ND2OPTIBD1BWP30P140LVT U85 ( .A1(n67), .A2(i_data_bus[58]), .ZN(n41) );
  ND2D1BWP30P140LVT U86 ( .A1(n68), .A2(i_data_bus[26]), .ZN(n40) );
  ND2D1BWP30P140LVT U87 ( .A1(n43), .A2(n42), .ZN(N119) );
  ND2OPTIBD1BWP30P140LVT U88 ( .A1(n67), .A2(i_data_bus[59]), .ZN(n43) );
  ND2D1BWP30P140LVT U89 ( .A1(n68), .A2(i_data_bus[27]), .ZN(n42) );
  ND2D1BWP30P140LVT U90 ( .A1(n45), .A2(n44), .ZN(N120) );
  ND2OPTIBD1BWP30P140LVT U91 ( .A1(n67), .A2(i_data_bus[60]), .ZN(n45) );
  ND2D1BWP30P140LVT U92 ( .A1(n68), .A2(i_data_bus[28]), .ZN(n44) );
  ND2D1BWP30P140LVT U93 ( .A1(n47), .A2(n46), .ZN(N121) );
  ND2OPTIBD1BWP30P140LVT U94 ( .A1(n67), .A2(i_data_bus[61]), .ZN(n47) );
  ND2D1BWP30P140LVT U95 ( .A1(n68), .A2(i_data_bus[29]), .ZN(n46) );
  ND2D1BWP30P140LVT U96 ( .A1(n49), .A2(n48), .ZN(N122) );
  ND2OPTIBD1BWP30P140LVT U97 ( .A1(n67), .A2(i_data_bus[62]), .ZN(n49) );
  ND2D1BWP30P140LVT U98 ( .A1(n68), .A2(i_data_bus[30]), .ZN(n48) );
  ND2D1BWP30P140LVT U99 ( .A1(n51), .A2(n50), .ZN(N123) );
  ND2OPTIBD1BWP30P140LVT U100 ( .A1(n67), .A2(i_data_bus[63]), .ZN(n51) );
  ND2D1BWP30P140LVT U101 ( .A1(n68), .A2(i_data_bus[31]), .ZN(n50) );
  IND2D1BWP30P140LVT U102 ( .A1(n67), .B1(n52), .ZN(N91) );
  INVD1BWP30P140LVT U103 ( .I(n68), .ZN(n52) );
  ND3D1BWP30P140LVT U104 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n1)
         );
  NR2D1BWP30P140LVT U105 ( .A1(n1), .A2(rst), .ZN(n2) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_12 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_12 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_2 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_12 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_11 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_10 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_9 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_8 o_data_high ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_7 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_13 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n4), .A2(n3), .ZN(n2) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n4) );
  INVD1BWP30P140LVT U5 ( .I(n7), .ZN(n8) );
  NR2D1BWP30P140LVT U6 ( .A1(n4), .A2(n3), .ZN(n1) );
  INVD1BWP30P140LVT U7 ( .I(n8), .ZN(n36) );
  INVD1BWP30P140LVT U8 ( .I(n8), .ZN(n41) );
  OR2D1BWP30P140LVT U9 ( .A1(rst), .A2(i_cmd[0]), .Z(n3) );
  ND3D1BWP30P140LVT U10 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n6)
         );
  INVD1BWP30P140LVT U11 ( .I(rst), .ZN(n5) );
  IND2D1BWP30P140LVT U12 ( .A1(n6), .B1(n5), .ZN(n7) );
  IND2D1BWP30P140LVT U13 ( .A1(n2), .B1(n41), .ZN(N91) );
  INVD1BWP30P140LVT U14 ( .I(i_data_bus[54]), .ZN(n9) );
  MOAI22D1BWP30P140LVT U15 ( .A1(n9), .A2(n36), .B1(i_data_bus[22]), .B2(n2), 
        .ZN(N114) );
  INVD1BWP30P140LVT U16 ( .I(i_data_bus[50]), .ZN(n10) );
  MOAI22D1BWP30P140LVT U17 ( .A1(n10), .A2(n36), .B1(i_data_bus[18]), .B2(n1), 
        .ZN(N110) );
  INVD1BWP30P140LVT U18 ( .I(i_data_bus[48]), .ZN(n11) );
  MOAI22D1BWP30P140LVT U19 ( .A1(n11), .A2(n36), .B1(i_data_bus[16]), .B2(n2), 
        .ZN(N108) );
  INVD1BWP30P140LVT U20 ( .I(i_data_bus[52]), .ZN(n12) );
  MOAI22D1BWP30P140LVT U21 ( .A1(n12), .A2(n36), .B1(i_data_bus[20]), .B2(n1), 
        .ZN(N112) );
  INVD1BWP30P140LVT U22 ( .I(i_data_bus[41]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U23 ( .A1(n13), .A2(n41), .B1(i_data_bus[9]), .B2(n2), 
        .ZN(N101) );
  INVD1BWP30P140LVT U24 ( .I(i_data_bus[42]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U25 ( .A1(n14), .A2(n41), .B1(i_data_bus[10]), .B2(n1), 
        .ZN(N102) );
  INVD1BWP30P140LVT U26 ( .I(i_data_bus[43]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U27 ( .A1(n15), .A2(n41), .B1(i_data_bus[11]), .B2(n2), 
        .ZN(N103) );
  INVD1BWP30P140LVT U28 ( .I(i_data_bus[40]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U29 ( .A1(n16), .A2(n41), .B1(i_data_bus[8]), .B2(n1), 
        .ZN(N100) );
  INVD1BWP30P140LVT U30 ( .I(i_data_bus[34]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U31 ( .A1(n17), .A2(n41), .B1(i_data_bus[2]), .B2(n2), 
        .ZN(N94) );
  INVD1BWP30P140LVT U32 ( .I(i_data_bus[35]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U33 ( .A1(n18), .A2(n41), .B1(i_data_bus[3]), .B2(n1), 
        .ZN(N95) );
  INVD1BWP30P140LVT U34 ( .I(i_data_bus[36]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U35 ( .A1(n19), .A2(n41), .B1(i_data_bus[4]), .B2(n2), 
        .ZN(N96) );
  INVD1BWP30P140LVT U36 ( .I(i_data_bus[32]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U37 ( .A1(n20), .A2(n41), .B1(i_data_bus[0]), .B2(n1), 
        .ZN(N92) );
  INVD1BWP30P140LVT U38 ( .I(i_data_bus[33]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U39 ( .A1(n21), .A2(n41), .B1(i_data_bus[1]), .B2(n2), 
        .ZN(N93) );
  INVD1BWP30P140LVT U40 ( .I(i_data_bus[39]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U41 ( .A1(n22), .A2(n41), .B1(i_data_bus[7]), .B2(n1), 
        .ZN(N99) );
  INVD1BWP30P140LVT U42 ( .I(i_data_bus[37]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U43 ( .A1(n23), .A2(n41), .B1(i_data_bus[5]), .B2(n2), 
        .ZN(N97) );
  INVD1BWP30P140LVT U44 ( .I(i_data_bus[38]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U45 ( .A1(n24), .A2(n41), .B1(i_data_bus[6]), .B2(n1), 
        .ZN(N98) );
  INVD1BWP30P140LVT U46 ( .I(i_data_bus[57]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U47 ( .A1(n25), .A2(n36), .B1(i_data_bus[25]), .B2(n1), 
        .ZN(N117) );
  INVD1BWP30P140LVT U48 ( .I(i_data_bus[61]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U49 ( .A1(n26), .A2(n36), .B1(i_data_bus[29]), .B2(n2), 
        .ZN(N121) );
  INVD1BWP30P140LVT U50 ( .I(i_data_bus[59]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U51 ( .A1(n27), .A2(n36), .B1(i_data_bus[27]), .B2(n1), 
        .ZN(N119) );
  INVD1BWP30P140LVT U52 ( .I(i_data_bus[55]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U53 ( .A1(n28), .A2(n36), .B1(i_data_bus[23]), .B2(n2), 
        .ZN(N115) );
  INVD1BWP30P140LVT U54 ( .I(i_data_bus[44]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U55 ( .A1(n29), .A2(n36), .B1(i_data_bus[12]), .B2(n1), 
        .ZN(N104) );
  INVD1BWP30P140LVT U56 ( .I(i_data_bus[63]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U57 ( .A1(n30), .A2(n36), .B1(i_data_bus[31]), .B2(n2), 
        .ZN(N123) );
  INVD1BWP30P140LVT U58 ( .I(i_data_bus[45]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U59 ( .A1(n31), .A2(n36), .B1(i_data_bus[13]), .B2(n1), 
        .ZN(N105) );
  INVD1BWP30P140LVT U60 ( .I(i_data_bus[53]), .ZN(n32) );
  MOAI22D1BWP30P140LVT U61 ( .A1(n32), .A2(n36), .B1(i_data_bus[21]), .B2(n2), 
        .ZN(N113) );
  INVD1BWP30P140LVT U62 ( .I(i_data_bus[47]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U63 ( .A1(n33), .A2(n36), .B1(i_data_bus[15]), .B2(n1), 
        .ZN(N107) );
  INVD1BWP30P140LVT U64 ( .I(i_data_bus[46]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U65 ( .A1(n34), .A2(n36), .B1(i_data_bus[14]), .B2(n2), 
        .ZN(N106) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[51]), .ZN(n35) );
  MOAI22D1BWP30P140LVT U67 ( .A1(n35), .A2(n36), .B1(i_data_bus[19]), .B2(n1), 
        .ZN(N111) );
  INVD1BWP30P140LVT U68 ( .I(i_data_bus[49]), .ZN(n37) );
  MOAI22D1BWP30P140LVT U69 ( .A1(n37), .A2(n36), .B1(i_data_bus[17]), .B2(n2), 
        .ZN(N109) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[56]), .ZN(n38) );
  MOAI22D1BWP30P140LVT U71 ( .A1(n38), .A2(n41), .B1(i_data_bus[24]), .B2(n1), 
        .ZN(N116) );
  INVD1BWP30P140LVT U72 ( .I(i_data_bus[62]), .ZN(n39) );
  MOAI22D1BWP30P140LVT U73 ( .A1(n39), .A2(n41), .B1(i_data_bus[30]), .B2(n2), 
        .ZN(N122) );
  INVD1BWP30P140LVT U74 ( .I(i_data_bus[58]), .ZN(n40) );
  MOAI22D1BWP30P140LVT U75 ( .A1(n40), .A2(n41), .B1(i_data_bus[26]), .B2(n1), 
        .ZN(N118) );
  INVD1BWP30P140LVT U76 ( .I(i_data_bus[60]), .ZN(n42) );
  MOAI22D1BWP30P140LVT U77 ( .A1(n42), .A2(n41), .B1(i_data_bus[28]), .B2(n2), 
        .ZN(N120) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_13 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_13 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_14 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n4), .A2(n3), .ZN(n2) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n4) );
  INVD1BWP30P140LVT U5 ( .I(n7), .ZN(n8) );
  NR2D1BWP30P140LVT U6 ( .A1(n4), .A2(n3), .ZN(n1) );
  INVD1BWP30P140LVT U7 ( .I(n8), .ZN(n36) );
  INVD1BWP30P140LVT U8 ( .I(n8), .ZN(n41) );
  OR2D1BWP30P140LVT U9 ( .A1(rst), .A2(i_cmd[0]), .Z(n3) );
  ND3D1BWP30P140LVT U10 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n6)
         );
  INVD1BWP30P140LVT U11 ( .I(rst), .ZN(n5) );
  IND2D1BWP30P140LVT U12 ( .A1(n6), .B1(n5), .ZN(n7) );
  IND2D1BWP30P140LVT U13 ( .A1(n2), .B1(n41), .ZN(N91) );
  INVD1BWP30P140LVT U14 ( .I(i_data_bus[50]), .ZN(n9) );
  MOAI22D1BWP30P140LVT U15 ( .A1(n9), .A2(n36), .B1(i_data_bus[18]), .B2(n2), 
        .ZN(N110) );
  INVD1BWP30P140LVT U16 ( .I(i_data_bus[48]), .ZN(n10) );
  MOAI22D1BWP30P140LVT U17 ( .A1(n10), .A2(n36), .B1(i_data_bus[16]), .B2(n1), 
        .ZN(N108) );
  INVD1BWP30P140LVT U18 ( .I(i_data_bus[54]), .ZN(n11) );
  MOAI22D1BWP30P140LVT U19 ( .A1(n11), .A2(n36), .B1(i_data_bus[22]), .B2(n2), 
        .ZN(N114) );
  INVD1BWP30P140LVT U20 ( .I(i_data_bus[52]), .ZN(n12) );
  MOAI22D1BWP30P140LVT U21 ( .A1(n12), .A2(n36), .B1(i_data_bus[20]), .B2(n1), 
        .ZN(N112) );
  INVD1BWP30P140LVT U22 ( .I(i_data_bus[36]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U23 ( .A1(n13), .A2(n41), .B1(i_data_bus[4]), .B2(n2), 
        .ZN(N96) );
  INVD1BWP30P140LVT U24 ( .I(i_data_bus[35]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U25 ( .A1(n14), .A2(n41), .B1(i_data_bus[3]), .B2(n1), 
        .ZN(N95) );
  INVD1BWP30P140LVT U26 ( .I(i_data_bus[34]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U27 ( .A1(n15), .A2(n41), .B1(i_data_bus[2]), .B2(n2), 
        .ZN(N94) );
  INVD1BWP30P140LVT U28 ( .I(i_data_bus[42]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U29 ( .A1(n16), .A2(n41), .B1(i_data_bus[10]), .B2(n1), 
        .ZN(N102) );
  INVD1BWP30P140LVT U30 ( .I(i_data_bus[41]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U31 ( .A1(n17), .A2(n41), .B1(i_data_bus[9]), .B2(n2), 
        .ZN(N101) );
  INVD1BWP30P140LVT U32 ( .I(i_data_bus[40]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U33 ( .A1(n18), .A2(n41), .B1(i_data_bus[8]), .B2(n1), 
        .ZN(N100) );
  INVD1BWP30P140LVT U34 ( .I(i_data_bus[39]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U35 ( .A1(n19), .A2(n41), .B1(i_data_bus[7]), .B2(n2), 
        .ZN(N99) );
  INVD1BWP30P140LVT U36 ( .I(i_data_bus[38]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U37 ( .A1(n20), .A2(n41), .B1(i_data_bus[6]), .B2(n1), 
        .ZN(N98) );
  INVD1BWP30P140LVT U38 ( .I(i_data_bus[43]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U39 ( .A1(n21), .A2(n41), .B1(i_data_bus[11]), .B2(n2), 
        .ZN(N103) );
  INVD1BWP30P140LVT U40 ( .I(i_data_bus[33]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U41 ( .A1(n22), .A2(n41), .B1(i_data_bus[1]), .B2(n1), 
        .ZN(N93) );
  INVD1BWP30P140LVT U42 ( .I(i_data_bus[37]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U43 ( .A1(n23), .A2(n41), .B1(i_data_bus[5]), .B2(n2), 
        .ZN(N97) );
  INVD1BWP30P140LVT U44 ( .I(i_data_bus[32]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U45 ( .A1(n24), .A2(n41), .B1(i_data_bus[0]), .B2(n1), 
        .ZN(N92) );
  INVD1BWP30P140LVT U46 ( .I(i_data_bus[44]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U47 ( .A1(n25), .A2(n36), .B1(i_data_bus[12]), .B2(n1), 
        .ZN(N104) );
  INVD1BWP30P140LVT U48 ( .I(i_data_bus[45]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U49 ( .A1(n26), .A2(n36), .B1(i_data_bus[13]), .B2(n2), 
        .ZN(N105) );
  INVD1BWP30P140LVT U50 ( .I(i_data_bus[46]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U51 ( .A1(n27), .A2(n36), .B1(i_data_bus[14]), .B2(n1), 
        .ZN(N106) );
  INVD1BWP30P140LVT U52 ( .I(i_data_bus[47]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U53 ( .A1(n28), .A2(n36), .B1(i_data_bus[15]), .B2(n2), 
        .ZN(N107) );
  INVD1BWP30P140LVT U54 ( .I(i_data_bus[49]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U55 ( .A1(n29), .A2(n36), .B1(i_data_bus[17]), .B2(n1), 
        .ZN(N109) );
  INVD1BWP30P140LVT U56 ( .I(i_data_bus[51]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U57 ( .A1(n30), .A2(n36), .B1(i_data_bus[19]), .B2(n2), 
        .ZN(N111) );
  INVD1BWP30P140LVT U58 ( .I(i_data_bus[53]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U59 ( .A1(n31), .A2(n36), .B1(i_data_bus[21]), .B2(n1), 
        .ZN(N113) );
  INVD1BWP30P140LVT U60 ( .I(i_data_bus[55]), .ZN(n32) );
  MOAI22D1BWP30P140LVT U61 ( .A1(n32), .A2(n36), .B1(i_data_bus[23]), .B2(n2), 
        .ZN(N115) );
  INVD1BWP30P140LVT U62 ( .I(i_data_bus[57]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U63 ( .A1(n33), .A2(n36), .B1(i_data_bus[25]), .B2(n1), 
        .ZN(N117) );
  INVD1BWP30P140LVT U64 ( .I(i_data_bus[59]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U65 ( .A1(n34), .A2(n36), .B1(i_data_bus[27]), .B2(n2), 
        .ZN(N119) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[63]), .ZN(n35) );
  MOAI22D1BWP30P140LVT U67 ( .A1(n35), .A2(n36), .B1(i_data_bus[31]), .B2(n1), 
        .ZN(N123) );
  INVD1BWP30P140LVT U68 ( .I(i_data_bus[61]), .ZN(n37) );
  MOAI22D1BWP30P140LVT U69 ( .A1(n37), .A2(n36), .B1(i_data_bus[29]), .B2(n2), 
        .ZN(N121) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[56]), .ZN(n38) );
  MOAI22D1BWP30P140LVT U71 ( .A1(n38), .A2(n41), .B1(i_data_bus[24]), .B2(n1), 
        .ZN(N116) );
  INVD1BWP30P140LVT U72 ( .I(i_data_bus[60]), .ZN(n39) );
  MOAI22D1BWP30P140LVT U73 ( .A1(n39), .A2(n41), .B1(i_data_bus[28]), .B2(n2), 
        .ZN(N120) );
  INVD1BWP30P140LVT U74 ( .I(i_data_bus[58]), .ZN(n40) );
  MOAI22D1BWP30P140LVT U75 ( .A1(n40), .A2(n41), .B1(i_data_bus[26]), .B2(n1), 
        .ZN(N118) );
  INVD1BWP30P140LVT U76 ( .I(i_data_bus[62]), .ZN(n42) );
  MOAI22D1BWP30P140LVT U77 ( .A1(n42), .A2(n41), .B1(i_data_bus[30]), .B2(n2), 
        .ZN(N122) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_14 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_14 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_15 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U36 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_15 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_15 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_16 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  IND2D1BWP30P140LVT U3 ( .A1(n1), .B1(i_valid[0]), .ZN(n2) );
  INVD1BWP30P140LVT U4 ( .I(i_en), .ZN(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  NR3D1P5BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n6) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  BUFFD2BWP30P140LVT U8 ( .I(n4), .Z(n5) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n5), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n5), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n5), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n5), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n5), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n5), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n5), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n5), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n5), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n5), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n5), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n5), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n5), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n5), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n5), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n5), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n5), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n5), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n5), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n5), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n5), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n5), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n5), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n5), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n5), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n5), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n5), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n5), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n5), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n5), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n5), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n5), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n5), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_16 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_16 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_17 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n33, n34, n35,
         n36, n37;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  NR2D1BWP30P140LVT U3 ( .A1(n35), .A2(rst), .ZN(n36) );
  NR3D1P5BWP30P140LVT U4 ( .A1(n34), .A2(i_cmd[0]), .A3(rst), .ZN(n33) );
  ND2OPTIBD2BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n34) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n35)
         );
  BUFFD2BWP30P140LVT U7 ( .I(n36), .Z(n37) );
  AO22D1BWP30P140LVT U8 ( .A1(n33), .A2(i_data_bus[0]), .B1(n37), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n33), .A2(i_data_bus[1]), .B1(n37), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n33), .A2(i_data_bus[2]), .B1(n37), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n33), .A2(i_data_bus[3]), .B1(n37), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n33), .A2(i_data_bus[4]), .B1(n37), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n33), .A2(i_data_bus[5]), .B1(n37), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n33), .A2(i_data_bus[6]), .B1(n37), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n33), .A2(i_data_bus[7]), .B1(n37), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n33), .A2(i_data_bus[8]), .B1(n37), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n33), .A2(i_data_bus[9]), .B1(n37), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n33), .A2(i_data_bus[10]), .B1(n37), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n33), .A2(i_data_bus[11]), .B1(n37), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n33), .A2(i_data_bus[12]), .B1(n37), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n33), .A2(i_data_bus[13]), .B1(n37), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n33), .A2(i_data_bus[14]), .B1(n37), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n33), .A2(i_data_bus[15]), .B1(n37), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n33), .A2(i_data_bus[16]), .B1(n37), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n33), .A2(i_data_bus[17]), .B1(n37), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n33), .A2(i_data_bus[18]), .B1(n37), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n33), .A2(i_data_bus[19]), .B1(n37), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n33), .A2(i_data_bus[20]), .B1(n37), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n33), .A2(i_data_bus[21]), .B1(n37), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n33), .A2(i_data_bus[22]), .B1(n37), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n33), .A2(i_data_bus[23]), .B1(n37), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n33), .A2(i_data_bus[24]), .B1(n37), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n33), .A2(i_data_bus[25]), .B1(n37), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n33), .A2(i_data_bus[26]), .B1(n37), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n33), .A2(i_data_bus[27]), .B1(n37), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n33), .A2(i_data_bus[28]), .B1(n37), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n33), .A2(i_data_bus[29]), .B1(n37), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n33), .A2(i_data_bus[30]), .B1(n37), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n33), .A2(i_data_bus[31]), .B1(n37), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n33), .A2(n37), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_17 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_17 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_18 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n33, n34, n35,
         n36, n37;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  ND2OPTIBD1BWP30P140LVT U3 ( .A1(i_valid[0]), .A2(i_en), .ZN(n34) );
  NR2D1BWP30P140LVT U4 ( .A1(n35), .A2(rst), .ZN(n36) );
  NR3D1P5BWP30P140LVT U5 ( .A1(n34), .A2(i_cmd[0]), .A3(rst), .ZN(n33) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n35)
         );
  BUFFD2BWP30P140LVT U7 ( .I(n36), .Z(n37) );
  AO22D1BWP30P140LVT U8 ( .A1(n33), .A2(i_data_bus[0]), .B1(n37), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n33), .A2(i_data_bus[1]), .B1(n37), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n33), .A2(i_data_bus[2]), .B1(n37), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n33), .A2(i_data_bus[3]), .B1(n37), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n33), .A2(i_data_bus[4]), .B1(n37), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n33), .A2(i_data_bus[5]), .B1(n37), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n33), .A2(i_data_bus[6]), .B1(n37), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n33), .A2(i_data_bus[7]), .B1(n37), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n33), .A2(i_data_bus[8]), .B1(n37), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n33), .A2(i_data_bus[9]), .B1(n37), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n33), .A2(i_data_bus[10]), .B1(n37), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n33), .A2(i_data_bus[11]), .B1(n37), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n33), .A2(i_data_bus[12]), .B1(n37), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n33), .A2(i_data_bus[13]), .B1(n37), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n33), .A2(i_data_bus[14]), .B1(n37), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n33), .A2(i_data_bus[15]), .B1(n37), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n33), .A2(i_data_bus[16]), .B1(n37), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n33), .A2(i_data_bus[17]), .B1(n37), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n33), .A2(i_data_bus[18]), .B1(n37), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n33), .A2(i_data_bus[19]), .B1(n37), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n33), .A2(i_data_bus[20]), .B1(n37), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n33), .A2(i_data_bus[21]), .B1(n37), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n33), .A2(i_data_bus[22]), .B1(n37), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n33), .A2(i_data_bus[23]), .B1(n37), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n33), .A2(i_data_bus[24]), .B1(n37), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n33), .A2(i_data_bus[25]), .B1(n37), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n33), .A2(i_data_bus[26]), .B1(n37), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n33), .A2(i_data_bus[27]), .B1(n37), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n33), .A2(i_data_bus[28]), .B1(n37), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n33), .A2(i_data_bus[29]), .B1(n37), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n33), .A2(i_data_bus[30]), .B1(n37), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n33), .A2(i_data_bus[31]), .B1(n37), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n33), .A2(n37), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_18 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_18 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_3 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_18 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_17 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_16 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_15 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_14 o_data_high ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_13 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_19 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n4), .A2(n3), .ZN(n2) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n4) );
  INVD1BWP30P140LVT U5 ( .I(n7), .ZN(n8) );
  IND2D1BWP30P140LVT U6 ( .A1(n6), .B1(n5), .ZN(n7) );
  NR2D1BWP30P140LVT U7 ( .A1(n4), .A2(n3), .ZN(n1) );
  INVD1BWP30P140LVT U8 ( .I(n8), .ZN(n36) );
  INVD1BWP30P140LVT U9 ( .I(n8), .ZN(n41) );
  OR2D1BWP30P140LVT U10 ( .A1(rst), .A2(i_cmd[0]), .Z(n3) );
  ND3D1BWP30P140LVT U11 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n6)
         );
  INVD1BWP30P140LVT U12 ( .I(rst), .ZN(n5) );
  IND2D1BWP30P140LVT U13 ( .A1(n2), .B1(n41), .ZN(N91) );
  INVD1BWP30P140LVT U14 ( .I(i_data_bus[50]), .ZN(n9) );
  MOAI22D1BWP30P140LVT U15 ( .A1(n9), .A2(n36), .B1(i_data_bus[18]), .B2(n2), 
        .ZN(N110) );
  INVD1BWP30P140LVT U16 ( .I(i_data_bus[52]), .ZN(n10) );
  MOAI22D1BWP30P140LVT U17 ( .A1(n10), .A2(n36), .B1(i_data_bus[20]), .B2(n1), 
        .ZN(N112) );
  INVD1BWP30P140LVT U18 ( .I(i_data_bus[48]), .ZN(n11) );
  MOAI22D1BWP30P140LVT U19 ( .A1(n11), .A2(n36), .B1(i_data_bus[16]), .B2(n2), 
        .ZN(N108) );
  INVD1BWP30P140LVT U20 ( .I(i_data_bus[54]), .ZN(n12) );
  MOAI22D1BWP30P140LVT U21 ( .A1(n12), .A2(n36), .B1(i_data_bus[22]), .B2(n1), 
        .ZN(N114) );
  INVD1BWP30P140LVT U22 ( .I(i_data_bus[42]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U23 ( .A1(n13), .A2(n41), .B1(i_data_bus[10]), .B2(n2), 
        .ZN(N102) );
  INVD1BWP30P140LVT U24 ( .I(i_data_bus[32]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U25 ( .A1(n14), .A2(n41), .B1(i_data_bus[0]), .B2(n1), 
        .ZN(N92) );
  INVD1BWP30P140LVT U26 ( .I(i_data_bus[39]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U27 ( .A1(n15), .A2(n41), .B1(i_data_bus[7]), .B2(n2), 
        .ZN(N99) );
  INVD1BWP30P140LVT U28 ( .I(i_data_bus[41]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U29 ( .A1(n16), .A2(n41), .B1(i_data_bus[9]), .B2(n1), 
        .ZN(N101) );
  INVD1BWP30P140LVT U30 ( .I(i_data_bus[34]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U31 ( .A1(n17), .A2(n41), .B1(i_data_bus[2]), .B2(n2), 
        .ZN(N94) );
  INVD1BWP30P140LVT U32 ( .I(i_data_bus[38]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U33 ( .A1(n18), .A2(n41), .B1(i_data_bus[6]), .B2(n1), 
        .ZN(N98) );
  INVD1BWP30P140LVT U34 ( .I(i_data_bus[37]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U35 ( .A1(n19), .A2(n41), .B1(i_data_bus[5]), .B2(n2), 
        .ZN(N97) );
  INVD1BWP30P140LVT U36 ( .I(i_data_bus[36]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U37 ( .A1(n20), .A2(n41), .B1(i_data_bus[4]), .B2(n1), 
        .ZN(N96) );
  INVD1BWP30P140LVT U38 ( .I(i_data_bus[40]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U39 ( .A1(n21), .A2(n41), .B1(i_data_bus[8]), .B2(n2), 
        .ZN(N100) );
  INVD1BWP30P140LVT U40 ( .I(i_data_bus[43]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U41 ( .A1(n22), .A2(n41), .B1(i_data_bus[11]), .B2(n1), 
        .ZN(N103) );
  INVD1BWP30P140LVT U42 ( .I(i_data_bus[33]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U43 ( .A1(n23), .A2(n41), .B1(i_data_bus[1]), .B2(n2), 
        .ZN(N93) );
  INVD1BWP30P140LVT U44 ( .I(i_data_bus[35]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U45 ( .A1(n24), .A2(n41), .B1(i_data_bus[3]), .B2(n1), 
        .ZN(N95) );
  INVD1BWP30P140LVT U46 ( .I(i_data_bus[44]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U47 ( .A1(n25), .A2(n36), .B1(i_data_bus[12]), .B2(n1), 
        .ZN(N104) );
  INVD1BWP30P140LVT U48 ( .I(i_data_bus[47]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U49 ( .A1(n26), .A2(n36), .B1(i_data_bus[15]), .B2(n2), 
        .ZN(N107) );
  INVD1BWP30P140LVT U50 ( .I(i_data_bus[51]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U51 ( .A1(n27), .A2(n36), .B1(i_data_bus[19]), .B2(n1), 
        .ZN(N111) );
  INVD1BWP30P140LVT U52 ( .I(i_data_bus[63]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U53 ( .A1(n28), .A2(n36), .B1(i_data_bus[31]), .B2(n2), 
        .ZN(N123) );
  INVD1BWP30P140LVT U54 ( .I(i_data_bus[61]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U55 ( .A1(n29), .A2(n36), .B1(i_data_bus[29]), .B2(n1), 
        .ZN(N121) );
  INVD1BWP30P140LVT U56 ( .I(i_data_bus[57]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U57 ( .A1(n30), .A2(n36), .B1(i_data_bus[25]), .B2(n2), 
        .ZN(N117) );
  INVD1BWP30P140LVT U58 ( .I(i_data_bus[59]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U59 ( .A1(n31), .A2(n36), .B1(i_data_bus[27]), .B2(n1), 
        .ZN(N119) );
  INVD1BWP30P140LVT U60 ( .I(i_data_bus[55]), .ZN(n32) );
  MOAI22D1BWP30P140LVT U61 ( .A1(n32), .A2(n36), .B1(i_data_bus[23]), .B2(n2), 
        .ZN(N115) );
  INVD1BWP30P140LVT U62 ( .I(i_data_bus[45]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U63 ( .A1(n33), .A2(n36), .B1(i_data_bus[13]), .B2(n1), 
        .ZN(N105) );
  INVD1BWP30P140LVT U64 ( .I(i_data_bus[53]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U65 ( .A1(n34), .A2(n36), .B1(i_data_bus[21]), .B2(n2), 
        .ZN(N113) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[49]), .ZN(n35) );
  MOAI22D1BWP30P140LVT U67 ( .A1(n35), .A2(n36), .B1(i_data_bus[17]), .B2(n1), 
        .ZN(N109) );
  INVD1BWP30P140LVT U68 ( .I(i_data_bus[46]), .ZN(n37) );
  MOAI22D1BWP30P140LVT U69 ( .A1(n37), .A2(n36), .B1(i_data_bus[14]), .B2(n2), 
        .ZN(N106) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[58]), .ZN(n38) );
  MOAI22D1BWP30P140LVT U71 ( .A1(n38), .A2(n41), .B1(i_data_bus[26]), .B2(n1), 
        .ZN(N118) );
  INVD1BWP30P140LVT U72 ( .I(i_data_bus[62]), .ZN(n39) );
  MOAI22D1BWP30P140LVT U73 ( .A1(n39), .A2(n41), .B1(i_data_bus[30]), .B2(n2), 
        .ZN(N122) );
  INVD1BWP30P140LVT U74 ( .I(i_data_bus[56]), .ZN(n40) );
  MOAI22D1BWP30P140LVT U75 ( .A1(n40), .A2(n41), .B1(i_data_bus[24]), .B2(n1), 
        .ZN(N116) );
  INVD1BWP30P140LVT U76 ( .I(i_data_bus[60]), .ZN(n42) );
  MOAI22D1BWP30P140LVT U77 ( .A1(n42), .A2(n41), .B1(i_data_bus[28]), .B2(n2), 
        .ZN(N120) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_19 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_19 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_20 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n4), .A2(n3), .ZN(n2) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n4) );
  INVD1BWP30P140LVT U5 ( .I(n7), .ZN(n8) );
  IND2D1BWP30P140LVT U6 ( .A1(n6), .B1(n5), .ZN(n7) );
  NR2D1BWP30P140LVT U7 ( .A1(n4), .A2(n3), .ZN(n1) );
  INVD1BWP30P140LVT U8 ( .I(n8), .ZN(n36) );
  INVD1BWP30P140LVT U9 ( .I(n8), .ZN(n41) );
  OR2D1BWP30P140LVT U10 ( .A1(rst), .A2(i_cmd[0]), .Z(n3) );
  ND3D1BWP30P140LVT U11 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n6)
         );
  INVD1BWP30P140LVT U12 ( .I(rst), .ZN(n5) );
  IND2D1BWP30P140LVT U13 ( .A1(n2), .B1(n41), .ZN(N91) );
  INVD1BWP30P140LVT U14 ( .I(i_data_bus[54]), .ZN(n9) );
  MOAI22D1BWP30P140LVT U15 ( .A1(n9), .A2(n36), .B1(i_data_bus[22]), .B2(n2), 
        .ZN(N114) );
  INVD1BWP30P140LVT U16 ( .I(i_data_bus[52]), .ZN(n10) );
  MOAI22D1BWP30P140LVT U17 ( .A1(n10), .A2(n36), .B1(i_data_bus[20]), .B2(n1), 
        .ZN(N112) );
  INVD1BWP30P140LVT U18 ( .I(i_data_bus[50]), .ZN(n11) );
  MOAI22D1BWP30P140LVT U19 ( .A1(n11), .A2(n36), .B1(i_data_bus[18]), .B2(n2), 
        .ZN(N110) );
  INVD1BWP30P140LVT U20 ( .I(i_data_bus[48]), .ZN(n12) );
  MOAI22D1BWP30P140LVT U21 ( .A1(n12), .A2(n36), .B1(i_data_bus[16]), .B2(n1), 
        .ZN(N108) );
  INVD1BWP30P140LVT U22 ( .I(i_data_bus[38]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U23 ( .A1(n13), .A2(n41), .B1(i_data_bus[6]), .B2(n2), 
        .ZN(N98) );
  INVD1BWP30P140LVT U24 ( .I(i_data_bus[39]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U25 ( .A1(n14), .A2(n41), .B1(i_data_bus[7]), .B2(n1), 
        .ZN(N99) );
  INVD1BWP30P140LVT U26 ( .I(i_data_bus[35]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U27 ( .A1(n15), .A2(n41), .B1(i_data_bus[3]), .B2(n2), 
        .ZN(N95) );
  INVD1BWP30P140LVT U28 ( .I(i_data_bus[34]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U29 ( .A1(n16), .A2(n41), .B1(i_data_bus[2]), .B2(n1), 
        .ZN(N94) );
  INVD1BWP30P140LVT U30 ( .I(i_data_bus[36]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U31 ( .A1(n17), .A2(n41), .B1(i_data_bus[4]), .B2(n2), 
        .ZN(N96) );
  INVD1BWP30P140LVT U32 ( .I(i_data_bus[33]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U33 ( .A1(n18), .A2(n41), .B1(i_data_bus[1]), .B2(n1), 
        .ZN(N93) );
  INVD1BWP30P140LVT U34 ( .I(i_data_bus[32]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U35 ( .A1(n19), .A2(n41), .B1(i_data_bus[0]), .B2(n2), 
        .ZN(N92) );
  INVD1BWP30P140LVT U36 ( .I(i_data_bus[37]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U37 ( .A1(n20), .A2(n41), .B1(i_data_bus[5]), .B2(n1), 
        .ZN(N97) );
  INVD1BWP30P140LVT U38 ( .I(i_data_bus[43]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U39 ( .A1(n21), .A2(n41), .B1(i_data_bus[11]), .B2(n2), 
        .ZN(N103) );
  INVD1BWP30P140LVT U40 ( .I(i_data_bus[42]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U41 ( .A1(n22), .A2(n41), .B1(i_data_bus[10]), .B2(n1), 
        .ZN(N102) );
  INVD1BWP30P140LVT U42 ( .I(i_data_bus[41]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U43 ( .A1(n23), .A2(n41), .B1(i_data_bus[9]), .B2(n2), 
        .ZN(N101) );
  INVD1BWP30P140LVT U44 ( .I(i_data_bus[40]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U45 ( .A1(n24), .A2(n41), .B1(i_data_bus[8]), .B2(n1), 
        .ZN(N100) );
  INVD1BWP30P140LVT U46 ( .I(i_data_bus[57]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U47 ( .A1(n25), .A2(n36), .B1(i_data_bus[25]), .B2(n1), 
        .ZN(N117) );
  INVD1BWP30P140LVT U48 ( .I(i_data_bus[59]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U49 ( .A1(n26), .A2(n36), .B1(i_data_bus[27]), .B2(n2), 
        .ZN(N119) );
  INVD1BWP30P140LVT U50 ( .I(i_data_bus[46]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U51 ( .A1(n27), .A2(n36), .B1(i_data_bus[14]), .B2(n1), 
        .ZN(N106) );
  INVD1BWP30P140LVT U52 ( .I(i_data_bus[44]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U53 ( .A1(n28), .A2(n36), .B1(i_data_bus[12]), .B2(n2), 
        .ZN(N104) );
  INVD1BWP30P140LVT U54 ( .I(i_data_bus[47]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U55 ( .A1(n29), .A2(n36), .B1(i_data_bus[15]), .B2(n1), 
        .ZN(N107) );
  INVD1BWP30P140LVT U56 ( .I(i_data_bus[53]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U57 ( .A1(n30), .A2(n36), .B1(i_data_bus[21]), .B2(n2), 
        .ZN(N113) );
  INVD1BWP30P140LVT U58 ( .I(i_data_bus[45]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U59 ( .A1(n31), .A2(n36), .B1(i_data_bus[13]), .B2(n1), 
        .ZN(N105) );
  INVD1BWP30P140LVT U60 ( .I(i_data_bus[63]), .ZN(n32) );
  MOAI22D1BWP30P140LVT U61 ( .A1(n32), .A2(n36), .B1(i_data_bus[31]), .B2(n2), 
        .ZN(N123) );
  INVD1BWP30P140LVT U62 ( .I(i_data_bus[49]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U63 ( .A1(n33), .A2(n36), .B1(i_data_bus[17]), .B2(n1), 
        .ZN(N109) );
  INVD1BWP30P140LVT U64 ( .I(i_data_bus[51]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U65 ( .A1(n34), .A2(n36), .B1(i_data_bus[19]), .B2(n2), 
        .ZN(N111) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[61]), .ZN(n35) );
  MOAI22D1BWP30P140LVT U67 ( .A1(n35), .A2(n36), .B1(i_data_bus[29]), .B2(n1), 
        .ZN(N121) );
  INVD1BWP30P140LVT U68 ( .I(i_data_bus[55]), .ZN(n37) );
  MOAI22D1BWP30P140LVT U69 ( .A1(n37), .A2(n36), .B1(i_data_bus[23]), .B2(n2), 
        .ZN(N115) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[62]), .ZN(n38) );
  MOAI22D1BWP30P140LVT U71 ( .A1(n38), .A2(n41), .B1(i_data_bus[30]), .B2(n1), 
        .ZN(N122) );
  INVD1BWP30P140LVT U72 ( .I(i_data_bus[58]), .ZN(n39) );
  MOAI22D1BWP30P140LVT U73 ( .A1(n39), .A2(n41), .B1(i_data_bus[26]), .B2(n2), 
        .ZN(N118) );
  INVD1BWP30P140LVT U74 ( .I(i_data_bus[56]), .ZN(n40) );
  MOAI22D1BWP30P140LVT U75 ( .A1(n40), .A2(n41), .B1(i_data_bus[24]), .B2(n1), 
        .ZN(N116) );
  INVD1BWP30P140LVT U76 ( .I(i_data_bus[60]), .ZN(n42) );
  MOAI22D1BWP30P140LVT U77 ( .A1(n42), .A2(n41), .B1(i_data_bus[28]), .B2(n2), 
        .ZN(N120) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_20 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_20 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_21 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U36 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_21 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_21 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_22 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_22 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_22 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_23 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_23 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_23 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_24 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_24 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_24 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_4 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_24 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_23 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_22 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_21 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_20 o_data_high ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_19 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_25 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  INVD1BWP30P140LVT U3 ( .I(n5), .ZN(n6) );
  IND2D1BWP30P140LVT U4 ( .A1(n4), .B1(n3), .ZN(n5) );
  INVD1BWP30P140LVT U5 ( .I(n6), .ZN(n35) );
  ND2D1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  INVD1BWP30P140LVT U7 ( .I(n6), .ZN(n41) );
  OR2D1BWP30P140LVT U8 ( .A1(rst), .A2(i_cmd[0]), .Z(n1) );
  OR2D1BWP30P140LVT U9 ( .A1(n2), .A2(n1), .Z(n7) );
  INVD2BWP30P140LVT U10 ( .I(n7), .ZN(n40) );
  ND3D1BWP30P140LVT U11 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n4)
         );
  INVD1BWP30P140LVT U12 ( .I(rst), .ZN(n3) );
  IND2D1BWP30P140LVT U13 ( .A1(n40), .B1(n41), .ZN(N91) );
  INVD1BWP30P140LVT U14 ( .I(i_data_bus[52]), .ZN(n8) );
  MOAI22D1BWP30P140LVT U15 ( .A1(n8), .A2(n35), .B1(i_data_bus[20]), .B2(n40), 
        .ZN(N112) );
  INVD1BWP30P140LVT U16 ( .I(i_data_bus[54]), .ZN(n9) );
  MOAI22D1BWP30P140LVT U17 ( .A1(n9), .A2(n35), .B1(i_data_bus[22]), .B2(n40), 
        .ZN(N114) );
  INVD1BWP30P140LVT U18 ( .I(i_data_bus[48]), .ZN(n10) );
  MOAI22D1BWP30P140LVT U19 ( .A1(n10), .A2(n35), .B1(i_data_bus[16]), .B2(n40), 
        .ZN(N108) );
  INVD1BWP30P140LVT U20 ( .I(i_data_bus[50]), .ZN(n11) );
  MOAI22D1BWP30P140LVT U21 ( .A1(n11), .A2(n35), .B1(i_data_bus[18]), .B2(n40), 
        .ZN(N110) );
  INVD1BWP30P140LVT U22 ( .I(i_data_bus[41]), .ZN(n12) );
  MOAI22D1BWP30P140LVT U23 ( .A1(n12), .A2(n41), .B1(i_data_bus[9]), .B2(n40), 
        .ZN(N101) );
  INVD1BWP30P140LVT U24 ( .I(i_data_bus[43]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U25 ( .A1(n13), .A2(n41), .B1(i_data_bus[11]), .B2(n40), 
        .ZN(N103) );
  INVD1BWP30P140LVT U26 ( .I(i_data_bus[35]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U27 ( .A1(n14), .A2(n41), .B1(i_data_bus[3]), .B2(n40), 
        .ZN(N95) );
  INVD1BWP30P140LVT U28 ( .I(i_data_bus[34]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U29 ( .A1(n15), .A2(n41), .B1(i_data_bus[2]), .B2(n40), 
        .ZN(N94) );
  INVD1BWP30P140LVT U30 ( .I(i_data_bus[42]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U31 ( .A1(n16), .A2(n41), .B1(i_data_bus[10]), .B2(n40), 
        .ZN(N102) );
  INVD1BWP30P140LVT U32 ( .I(i_data_bus[36]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U33 ( .A1(n17), .A2(n41), .B1(i_data_bus[4]), .B2(n40), 
        .ZN(N96) );
  INVD1BWP30P140LVT U34 ( .I(i_data_bus[39]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U35 ( .A1(n18), .A2(n41), .B1(i_data_bus[7]), .B2(n40), 
        .ZN(N99) );
  INVD1BWP30P140LVT U36 ( .I(i_data_bus[38]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U37 ( .A1(n19), .A2(n41), .B1(i_data_bus[6]), .B2(n40), 
        .ZN(N98) );
  INVD1BWP30P140LVT U38 ( .I(i_data_bus[37]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U39 ( .A1(n20), .A2(n41), .B1(i_data_bus[5]), .B2(n40), 
        .ZN(N97) );
  INVD1BWP30P140LVT U40 ( .I(i_data_bus[40]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U41 ( .A1(n21), .A2(n41), .B1(i_data_bus[8]), .B2(n40), 
        .ZN(N100) );
  INVD1BWP30P140LVT U42 ( .I(i_data_bus[33]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U43 ( .A1(n22), .A2(n41), .B1(i_data_bus[1]), .B2(n40), 
        .ZN(N93) );
  INVD1BWP30P140LVT U44 ( .I(i_data_bus[32]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U45 ( .A1(n23), .A2(n41), .B1(i_data_bus[0]), .B2(n40), 
        .ZN(N92) );
  INVD1BWP30P140LVT U46 ( .I(i_data_bus[44]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U47 ( .A1(n24), .A2(n35), .B1(i_data_bus[12]), .B2(n40), 
        .ZN(N104) );
  INVD1BWP30P140LVT U48 ( .I(i_data_bus[55]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U49 ( .A1(n25), .A2(n35), .B1(i_data_bus[23]), .B2(n40), 
        .ZN(N115) );
  INVD1BWP30P140LVT U50 ( .I(i_data_bus[53]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U51 ( .A1(n26), .A2(n35), .B1(i_data_bus[21]), .B2(n40), 
        .ZN(N113) );
  INVD1BWP30P140LVT U52 ( .I(i_data_bus[51]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U53 ( .A1(n27), .A2(n35), .B1(i_data_bus[19]), .B2(n40), 
        .ZN(N111) );
  INVD1BWP30P140LVT U54 ( .I(i_data_bus[47]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U55 ( .A1(n28), .A2(n35), .B1(i_data_bus[15]), .B2(n40), 
        .ZN(N107) );
  INVD1BWP30P140LVT U56 ( .I(i_data_bus[61]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U57 ( .A1(n29), .A2(n35), .B1(i_data_bus[29]), .B2(n40), 
        .ZN(N121) );
  INVD1BWP30P140LVT U58 ( .I(i_data_bus[59]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U59 ( .A1(n30), .A2(n35), .B1(i_data_bus[27]), .B2(n40), 
        .ZN(N119) );
  INVD1BWP30P140LVT U60 ( .I(i_data_bus[63]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U61 ( .A1(n31), .A2(n35), .B1(i_data_bus[31]), .B2(n40), 
        .ZN(N123) );
  INVD1BWP30P140LVT U62 ( .I(i_data_bus[49]), .ZN(n32) );
  MOAI22D1BWP30P140LVT U63 ( .A1(n32), .A2(n35), .B1(i_data_bus[17]), .B2(n40), 
        .ZN(N109) );
  INVD1BWP30P140LVT U64 ( .I(i_data_bus[46]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U65 ( .A1(n33), .A2(n35), .B1(i_data_bus[14]), .B2(n40), 
        .ZN(N106) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[57]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U67 ( .A1(n34), .A2(n35), .B1(i_data_bus[25]), .B2(n40), 
        .ZN(N117) );
  INVD1BWP30P140LVT U68 ( .I(i_data_bus[45]), .ZN(n36) );
  MOAI22D1BWP30P140LVT U69 ( .A1(n36), .A2(n35), .B1(i_data_bus[13]), .B2(n40), 
        .ZN(N105) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[62]), .ZN(n37) );
  MOAI22D1BWP30P140LVT U71 ( .A1(n37), .A2(n41), .B1(i_data_bus[30]), .B2(n40), 
        .ZN(N122) );
  INVD1BWP30P140LVT U72 ( .I(i_data_bus[58]), .ZN(n38) );
  MOAI22D1BWP30P140LVT U73 ( .A1(n38), .A2(n41), .B1(i_data_bus[26]), .B2(n40), 
        .ZN(N118) );
  INVD1BWP30P140LVT U74 ( .I(i_data_bus[60]), .ZN(n39) );
  MOAI22D1BWP30P140LVT U75 ( .A1(n39), .A2(n41), .B1(i_data_bus[28]), .B2(n40), 
        .ZN(N120) );
  INVD1BWP30P140LVT U76 ( .I(i_data_bus[56]), .ZN(n42) );
  MOAI22D1BWP30P140LVT U77 ( .A1(n42), .A2(n41), .B1(i_data_bus[24]), .B2(n40), 
        .ZN(N116) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_25 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_25 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_26 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D3BWP30P140LVT U3 ( .A1(n3), .A2(n2), .ZN(n1) );
  INVD1BWP30P140LVT U4 ( .I(n6), .ZN(n7) );
  IND2D1BWP30P140LVT U5 ( .A1(n5), .B1(n4), .ZN(n6) );
  INVD1BWP30P140LVT U6 ( .I(n7), .ZN(n35) );
  ND2D1BWP30P140LVT U7 ( .A1(i_en), .A2(i_valid[0]), .ZN(n3) );
  INVD1BWP30P140LVT U8 ( .I(n7), .ZN(n40) );
  OR2D1BWP30P140LVT U9 ( .A1(rst), .A2(i_cmd[0]), .Z(n2) );
  ND3D1BWP30P140LVT U10 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n5)
         );
  INVD1BWP30P140LVT U11 ( .I(rst), .ZN(n4) );
  IND2D1BWP30P140LVT U12 ( .A1(n1), .B1(n40), .ZN(N91) );
  INVD1BWP30P140LVT U13 ( .I(i_data_bus[48]), .ZN(n8) );
  MOAI22D1BWP30P140LVT U14 ( .A1(n8), .A2(n35), .B1(i_data_bus[16]), .B2(n1), 
        .ZN(N108) );
  INVD1BWP30P140LVT U15 ( .I(i_data_bus[54]), .ZN(n9) );
  MOAI22D1BWP30P140LVT U16 ( .A1(n9), .A2(n35), .B1(i_data_bus[22]), .B2(n1), 
        .ZN(N114) );
  INVD1BWP30P140LVT U17 ( .I(i_data_bus[52]), .ZN(n10) );
  MOAI22D1BWP30P140LVT U18 ( .A1(n10), .A2(n35), .B1(i_data_bus[20]), .B2(n1), 
        .ZN(N112) );
  INVD1BWP30P140LVT U19 ( .I(i_data_bus[50]), .ZN(n11) );
  MOAI22D1BWP30P140LVT U20 ( .A1(n11), .A2(n35), .B1(i_data_bus[18]), .B2(n1), 
        .ZN(N110) );
  INVD1BWP30P140LVT U21 ( .I(i_data_bus[36]), .ZN(n12) );
  MOAI22D1BWP30P140LVT U22 ( .A1(n12), .A2(n40), .B1(i_data_bus[4]), .B2(n1), 
        .ZN(N96) );
  INVD1BWP30P140LVT U23 ( .I(i_data_bus[37]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U24 ( .A1(n13), .A2(n40), .B1(i_data_bus[5]), .B2(n1), 
        .ZN(N97) );
  INVD1BWP30P140LVT U25 ( .I(i_data_bus[38]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U26 ( .A1(n14), .A2(n40), .B1(i_data_bus[6]), .B2(n1), 
        .ZN(N98) );
  INVD1BWP30P140LVT U27 ( .I(i_data_bus[34]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U28 ( .A1(n15), .A2(n40), .B1(i_data_bus[2]), .B2(n1), 
        .ZN(N94) );
  INVD1BWP30P140LVT U29 ( .I(i_data_bus[35]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U30 ( .A1(n16), .A2(n40), .B1(i_data_bus[3]), .B2(n1), 
        .ZN(N95) );
  INVD1BWP30P140LVT U31 ( .I(i_data_bus[41]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U32 ( .A1(n17), .A2(n40), .B1(i_data_bus[9]), .B2(n1), 
        .ZN(N101) );
  INVD1BWP30P140LVT U33 ( .I(i_data_bus[32]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U34 ( .A1(n18), .A2(n40), .B1(i_data_bus[0]), .B2(n1), 
        .ZN(N92) );
  INVD1BWP30P140LVT U35 ( .I(i_data_bus[40]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U36 ( .A1(n19), .A2(n40), .B1(i_data_bus[8]), .B2(n1), 
        .ZN(N100) );
  INVD1BWP30P140LVT U37 ( .I(i_data_bus[39]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U38 ( .A1(n20), .A2(n40), .B1(i_data_bus[7]), .B2(n1), 
        .ZN(N99) );
  INVD1BWP30P140LVT U39 ( .I(i_data_bus[42]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U40 ( .A1(n21), .A2(n40), .B1(i_data_bus[10]), .B2(n1), 
        .ZN(N102) );
  INVD1BWP30P140LVT U41 ( .I(i_data_bus[33]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U42 ( .A1(n22), .A2(n40), .B1(i_data_bus[1]), .B2(n1), 
        .ZN(N93) );
  INVD1BWP30P140LVT U43 ( .I(i_data_bus[43]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U44 ( .A1(n23), .A2(n40), .B1(i_data_bus[11]), .B2(n1), 
        .ZN(N103) );
  INVD1BWP30P140LVT U45 ( .I(i_data_bus[44]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U46 ( .A1(n24), .A2(n35), .B1(i_data_bus[12]), .B2(n1), 
        .ZN(N104) );
  INVD1BWP30P140LVT U47 ( .I(i_data_bus[55]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U48 ( .A1(n25), .A2(n35), .B1(i_data_bus[23]), .B2(n1), 
        .ZN(N115) );
  INVD1BWP30P140LVT U49 ( .I(i_data_bus[63]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U50 ( .A1(n26), .A2(n35), .B1(i_data_bus[31]), .B2(n1), 
        .ZN(N123) );
  INVD1BWP30P140LVT U51 ( .I(i_data_bus[57]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U52 ( .A1(n27), .A2(n35), .B1(i_data_bus[25]), .B2(n1), 
        .ZN(N117) );
  INVD1BWP30P140LVT U53 ( .I(i_data_bus[45]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U54 ( .A1(n28), .A2(n35), .B1(i_data_bus[13]), .B2(n1), 
        .ZN(N105) );
  INVD1BWP30P140LVT U55 ( .I(i_data_bus[59]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U56 ( .A1(n29), .A2(n35), .B1(i_data_bus[27]), .B2(n1), 
        .ZN(N119) );
  INVD1BWP30P140LVT U57 ( .I(i_data_bus[49]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U58 ( .A1(n30), .A2(n35), .B1(i_data_bus[17]), .B2(n1), 
        .ZN(N109) );
  INVD1BWP30P140LVT U59 ( .I(i_data_bus[61]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U60 ( .A1(n31), .A2(n35), .B1(i_data_bus[29]), .B2(n1), 
        .ZN(N121) );
  INVD1BWP30P140LVT U61 ( .I(i_data_bus[53]), .ZN(n32) );
  MOAI22D1BWP30P140LVT U62 ( .A1(n32), .A2(n35), .B1(i_data_bus[21]), .B2(n1), 
        .ZN(N113) );
  INVD1BWP30P140LVT U63 ( .I(i_data_bus[51]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U64 ( .A1(n33), .A2(n35), .B1(i_data_bus[19]), .B2(n1), 
        .ZN(N111) );
  INVD1BWP30P140LVT U65 ( .I(i_data_bus[47]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U66 ( .A1(n34), .A2(n35), .B1(i_data_bus[15]), .B2(n1), 
        .ZN(N107) );
  INVD1BWP30P140LVT U67 ( .I(i_data_bus[46]), .ZN(n36) );
  MOAI22D1BWP30P140LVT U68 ( .A1(n36), .A2(n35), .B1(i_data_bus[14]), .B2(n1), 
        .ZN(N106) );
  INVD1BWP30P140LVT U69 ( .I(i_data_bus[58]), .ZN(n37) );
  MOAI22D1BWP30P140LVT U70 ( .A1(n37), .A2(n40), .B1(i_data_bus[26]), .B2(n1), 
        .ZN(N118) );
  INVD1BWP30P140LVT U71 ( .I(i_data_bus[60]), .ZN(n38) );
  MOAI22D1BWP30P140LVT U72 ( .A1(n38), .A2(n40), .B1(i_data_bus[28]), .B2(n1), 
        .ZN(N120) );
  INVD1BWP30P140LVT U73 ( .I(i_data_bus[56]), .ZN(n39) );
  MOAI22D1BWP30P140LVT U74 ( .A1(n39), .A2(n40), .B1(i_data_bus[24]), .B2(n1), 
        .ZN(N116) );
  INVD1BWP30P140LVT U75 ( .I(i_data_bus[62]), .ZN(n41) );
  MOAI22D1BWP30P140LVT U76 ( .A1(n41), .A2(n40), .B1(i_data_bus[30]), .B2(n1), 
        .ZN(N122) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_26 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_26 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_27 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(i_cmd[0]), .A2(n2), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2OPTIBD1BWP30P140LVT U24 ( .A1(i_valid[0]), .A2(n1), .ZN(n2) );
  INR2D1BWP30P140LVT U25 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U36 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U37 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_27 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_27 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_28 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2OPTPAD1BWP30P140LVT U3 ( .A1(i_cmd[0]), .A2(n2), .ZN(n6) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_valid[0]), .A2(n1), .ZN(n2) );
  INR2D1BWP30P140LVT U5 ( .A1(i_en), .B1(rst), .ZN(n1) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  NR2D1BWP30P140LVT U7 ( .A1(n3), .A2(rst), .ZN(n4) );
  BUFFD2BWP30P140LVT U8 ( .I(n4), .Z(n5) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n5), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n5), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n5), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n5), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n5), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n5), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n5), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n5), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n5), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n5), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n5), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n5), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n5), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n5), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n5), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n5), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n5), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n5), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n5), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n5), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n5), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n5), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n5), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n5), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n5), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n5), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n5), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n5), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n5), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n5), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n5), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n5), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n5), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_28 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_28 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_29 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  INVD1BWP30P140LVT U3 ( .I(n4), .ZN(n69) );
  OR3D1BWP30P140LVT U4 ( .A1(n3), .A2(rst), .A3(i_cmd[0]), .Z(n4) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n3) );
  CKBD1BWP30P140LVT U6 ( .I(n68), .Z(n1) );
  NR2D1BWP30P140LVT U7 ( .A1(n2), .A2(rst), .ZN(n68) );
  IND2D1BWP30P140LVT U8 ( .A1(n1), .B1(n57), .ZN(N91) );
  INVD1BWP30P140LVT U9 ( .I(n69), .ZN(n57) );
  ND2OPTIBD1BWP30P140LVT U10 ( .A1(n59), .A2(n58), .ZN(N92) );
  ND2OPTIBD1BWP30P140LVT U11 ( .A1(n69), .A2(i_data_bus[0]), .ZN(n58) );
  ND2OPTIBD1BWP30P140LVT U12 ( .A1(n1), .A2(i_data_bus[32]), .ZN(n59) );
  ND2OPTIBD1BWP30P140LVT U13 ( .A1(n61), .A2(n60), .ZN(N93) );
  ND2OPTIBD1BWP30P140LVT U14 ( .A1(n69), .A2(i_data_bus[1]), .ZN(n60) );
  ND2OPTIBD1BWP30P140LVT U15 ( .A1(n1), .A2(i_data_bus[33]), .ZN(n61) );
  ND2OPTIBD1BWP30P140LVT U16 ( .A1(n63), .A2(n62), .ZN(N94) );
  ND2OPTIBD1BWP30P140LVT U17 ( .A1(n69), .A2(i_data_bus[2]), .ZN(n62) );
  ND2OPTIBD1BWP30P140LVT U18 ( .A1(n1), .A2(i_data_bus[34]), .ZN(n63) );
  ND2OPTIBD1BWP30P140LVT U19 ( .A1(n65), .A2(n64), .ZN(N95) );
  ND2OPTIBD1BWP30P140LVT U20 ( .A1(n69), .A2(i_data_bus[3]), .ZN(n64) );
  ND2OPTIBD1BWP30P140LVT U21 ( .A1(n1), .A2(i_data_bus[35]), .ZN(n65) );
  ND2OPTIBD1BWP30P140LVT U22 ( .A1(n67), .A2(n66), .ZN(N96) );
  ND2OPTIBD1BWP30P140LVT U23 ( .A1(n69), .A2(i_data_bus[4]), .ZN(n66) );
  ND2OPTIBD1BWP30P140LVT U24 ( .A1(n1), .A2(i_data_bus[36]), .ZN(n67) );
  ND2OPTIBD1BWP30P140LVT U25 ( .A1(n71), .A2(n70), .ZN(N97) );
  ND2OPTIBD1BWP30P140LVT U26 ( .A1(n69), .A2(i_data_bus[5]), .ZN(n70) );
  ND2OPTIBD1BWP30P140LVT U27 ( .A1(n1), .A2(i_data_bus[37]), .ZN(n71) );
  ND2OPTIBD1BWP30P140LVT U28 ( .A1(n6), .A2(n5), .ZN(N98) );
  ND2OPTIBD1BWP30P140LVT U29 ( .A1(n69), .A2(i_data_bus[6]), .ZN(n5) );
  ND2OPTIBD1BWP30P140LVT U30 ( .A1(n1), .A2(i_data_bus[38]), .ZN(n6) );
  ND2OPTIBD1BWP30P140LVT U31 ( .A1(n8), .A2(n7), .ZN(N99) );
  ND2OPTIBD1BWP30P140LVT U32 ( .A1(n69), .A2(i_data_bus[7]), .ZN(n7) );
  ND2OPTIBD1BWP30P140LVT U33 ( .A1(n1), .A2(i_data_bus[39]), .ZN(n8) );
  ND2OPTIBD1BWP30P140LVT U34 ( .A1(n10), .A2(n9), .ZN(N100) );
  ND2OPTIBD1BWP30P140LVT U35 ( .A1(n69), .A2(i_data_bus[8]), .ZN(n9) );
  ND2OPTIBD1BWP30P140LVT U36 ( .A1(n1), .A2(i_data_bus[40]), .ZN(n10) );
  ND2OPTIBD1BWP30P140LVT U37 ( .A1(n12), .A2(n11), .ZN(N101) );
  ND2OPTIBD1BWP30P140LVT U38 ( .A1(n69), .A2(i_data_bus[9]), .ZN(n11) );
  ND2OPTIBD1BWP30P140LVT U39 ( .A1(n1), .A2(i_data_bus[41]), .ZN(n12) );
  ND2OPTIBD1BWP30P140LVT U40 ( .A1(n14), .A2(n13), .ZN(N102) );
  ND2OPTIBD1BWP30P140LVT U41 ( .A1(n69), .A2(i_data_bus[10]), .ZN(n13) );
  ND2OPTIBD1BWP30P140LVT U42 ( .A1(n1), .A2(i_data_bus[42]), .ZN(n14) );
  ND2OPTIBD1BWP30P140LVT U43 ( .A1(n16), .A2(n15), .ZN(N103) );
  ND2OPTIBD1BWP30P140LVT U44 ( .A1(n69), .A2(i_data_bus[11]), .ZN(n15) );
  ND2OPTIBD1BWP30P140LVT U45 ( .A1(n1), .A2(i_data_bus[43]), .ZN(n16) );
  ND2OPTIBD1BWP30P140LVT U46 ( .A1(n18), .A2(n17), .ZN(N104) );
  ND2OPTIBD1BWP30P140LVT U47 ( .A1(n69), .A2(i_data_bus[12]), .ZN(n17) );
  ND2OPTIBD1BWP30P140LVT U48 ( .A1(n1), .A2(i_data_bus[44]), .ZN(n18) );
  ND2OPTIBD1BWP30P140LVT U49 ( .A1(n20), .A2(n19), .ZN(N105) );
  ND2OPTIBD1BWP30P140LVT U50 ( .A1(n69), .A2(i_data_bus[13]), .ZN(n19) );
  ND2OPTIBD1BWP30P140LVT U51 ( .A1(n1), .A2(i_data_bus[45]), .ZN(n20) );
  ND2OPTIBD1BWP30P140LVT U52 ( .A1(n22), .A2(n21), .ZN(N106) );
  ND2OPTIBD1BWP30P140LVT U53 ( .A1(n69), .A2(i_data_bus[14]), .ZN(n21) );
  ND2OPTIBD1BWP30P140LVT U54 ( .A1(n1), .A2(i_data_bus[46]), .ZN(n22) );
  ND2OPTIBD1BWP30P140LVT U55 ( .A1(n24), .A2(n23), .ZN(N107) );
  ND2OPTIBD1BWP30P140LVT U56 ( .A1(n69), .A2(i_data_bus[15]), .ZN(n23) );
  ND2OPTIBD1BWP30P140LVT U57 ( .A1(n1), .A2(i_data_bus[47]), .ZN(n24) );
  ND2OPTIBD1BWP30P140LVT U58 ( .A1(n26), .A2(n25), .ZN(N108) );
  ND2OPTIBD1BWP30P140LVT U59 ( .A1(n69), .A2(i_data_bus[16]), .ZN(n25) );
  ND2OPTIBD1BWP30P140LVT U60 ( .A1(n1), .A2(i_data_bus[48]), .ZN(n26) );
  ND2OPTIBD1BWP30P140LVT U61 ( .A1(n28), .A2(n27), .ZN(N109) );
  ND2OPTIBD1BWP30P140LVT U62 ( .A1(n69), .A2(i_data_bus[17]), .ZN(n27) );
  ND2OPTIBD1BWP30P140LVT U63 ( .A1(n1), .A2(i_data_bus[49]), .ZN(n28) );
  ND2OPTIBD1BWP30P140LVT U64 ( .A1(n30), .A2(n29), .ZN(N110) );
  ND2OPTIBD1BWP30P140LVT U65 ( .A1(n69), .A2(i_data_bus[18]), .ZN(n29) );
  ND2OPTIBD1BWP30P140LVT U66 ( .A1(n1), .A2(i_data_bus[50]), .ZN(n30) );
  ND2OPTIBD1BWP30P140LVT U67 ( .A1(n32), .A2(n31), .ZN(N111) );
  ND2OPTIBD1BWP30P140LVT U68 ( .A1(n69), .A2(i_data_bus[19]), .ZN(n31) );
  ND2OPTIBD1BWP30P140LVT U69 ( .A1(n1), .A2(i_data_bus[51]), .ZN(n32) );
  ND2OPTIBD1BWP30P140LVT U70 ( .A1(n34), .A2(n33), .ZN(N112) );
  ND2OPTIBD1BWP30P140LVT U71 ( .A1(n69), .A2(i_data_bus[20]), .ZN(n33) );
  ND2OPTIBD1BWP30P140LVT U72 ( .A1(n1), .A2(i_data_bus[52]), .ZN(n34) );
  ND2OPTIBD1BWP30P140LVT U73 ( .A1(n36), .A2(n35), .ZN(N113) );
  ND2OPTIBD1BWP30P140LVT U74 ( .A1(n69), .A2(i_data_bus[21]), .ZN(n35) );
  ND2OPTIBD1BWP30P140LVT U75 ( .A1(n1), .A2(i_data_bus[53]), .ZN(n36) );
  ND2OPTIBD1BWP30P140LVT U76 ( .A1(n38), .A2(n37), .ZN(N114) );
  ND2OPTIBD1BWP30P140LVT U77 ( .A1(n69), .A2(i_data_bus[22]), .ZN(n37) );
  ND2OPTIBD1BWP30P140LVT U78 ( .A1(n1), .A2(i_data_bus[54]), .ZN(n38) );
  ND2OPTIBD1BWP30P140LVT U79 ( .A1(n40), .A2(n39), .ZN(N115) );
  ND2OPTIBD1BWP30P140LVT U80 ( .A1(n69), .A2(i_data_bus[23]), .ZN(n39) );
  ND2OPTIBD1BWP30P140LVT U81 ( .A1(n1), .A2(i_data_bus[55]), .ZN(n40) );
  ND2OPTIBD1BWP30P140LVT U82 ( .A1(n42), .A2(n41), .ZN(N116) );
  ND2OPTIBD1BWP30P140LVT U83 ( .A1(n69), .A2(i_data_bus[24]), .ZN(n41) );
  ND2OPTIBD1BWP30P140LVT U84 ( .A1(n1), .A2(i_data_bus[56]), .ZN(n42) );
  ND2OPTIBD1BWP30P140LVT U85 ( .A1(n44), .A2(n43), .ZN(N117) );
  ND2OPTIBD1BWP30P140LVT U86 ( .A1(n69), .A2(i_data_bus[25]), .ZN(n43) );
  ND2OPTIBD1BWP30P140LVT U87 ( .A1(n1), .A2(i_data_bus[57]), .ZN(n44) );
  ND2OPTIBD1BWP30P140LVT U88 ( .A1(n46), .A2(n45), .ZN(N118) );
  ND2OPTIBD1BWP30P140LVT U89 ( .A1(n69), .A2(i_data_bus[26]), .ZN(n45) );
  ND2OPTIBD1BWP30P140LVT U90 ( .A1(n1), .A2(i_data_bus[58]), .ZN(n46) );
  ND2OPTIBD1BWP30P140LVT U91 ( .A1(n48), .A2(n47), .ZN(N119) );
  ND2OPTIBD1BWP30P140LVT U92 ( .A1(n69), .A2(i_data_bus[27]), .ZN(n47) );
  ND2OPTIBD1BWP30P140LVT U93 ( .A1(n1), .A2(i_data_bus[59]), .ZN(n48) );
  ND2OPTIBD1BWP30P140LVT U94 ( .A1(n50), .A2(n49), .ZN(N120) );
  ND2OPTIBD1BWP30P140LVT U95 ( .A1(n69), .A2(i_data_bus[28]), .ZN(n49) );
  ND2OPTIBD1BWP30P140LVT U96 ( .A1(n1), .A2(i_data_bus[60]), .ZN(n50) );
  ND2OPTIBD1BWP30P140LVT U97 ( .A1(n52), .A2(n51), .ZN(N121) );
  ND2OPTIBD1BWP30P140LVT U98 ( .A1(n69), .A2(i_data_bus[29]), .ZN(n51) );
  ND2OPTIBD1BWP30P140LVT U99 ( .A1(n1), .A2(i_data_bus[61]), .ZN(n52) );
  ND2OPTIBD1BWP30P140LVT U100 ( .A1(n54), .A2(n53), .ZN(N122) );
  ND2OPTIBD1BWP30P140LVT U101 ( .A1(n69), .A2(i_data_bus[30]), .ZN(n53) );
  ND2OPTIBD1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[62]), .ZN(n54) );
  ND2OPTIBD1BWP30P140LVT U103 ( .A1(n56), .A2(n55), .ZN(N123) );
  ND2OPTIBD1BWP30P140LVT U104 ( .A1(n69), .A2(i_data_bus[31]), .ZN(n55) );
  ND2OPTIBD1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[63]), .ZN(n56) );
  ND3D1BWP30P140LVT U106 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2)
         );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_29 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_29 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_30 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n2), .A2(rst), .ZN(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n2), .A2(rst), .ZN(n71) );
  INVD1BWP30P140LVT U5 ( .I(n4), .ZN(n69) );
  OR3D1BWP30P140LVT U6 ( .A1(n3), .A2(rst), .A3(i_cmd[0]), .Z(n4) );
  ND2D1BWP30P140LVT U7 ( .A1(i_en), .A2(i_valid[0]), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U8 ( .A1(n6), .A2(n5), .ZN(N92) );
  ND2OPTIBD1BWP30P140LVT U9 ( .A1(n69), .A2(i_data_bus[0]), .ZN(n5) );
  ND2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_data_bus[32]), .ZN(n6) );
  ND2OPTIBD1BWP30P140LVT U11 ( .A1(n8), .A2(n7), .ZN(N93) );
  ND2OPTIBD1BWP30P140LVT U12 ( .A1(n69), .A2(i_data_bus[1]), .ZN(n7) );
  ND2D1BWP30P140LVT U13 ( .A1(n71), .A2(i_data_bus[33]), .ZN(n8) );
  ND2OPTIBD1BWP30P140LVT U14 ( .A1(n10), .A2(n9), .ZN(N94) );
  ND2OPTIBD1BWP30P140LVT U15 ( .A1(n69), .A2(i_data_bus[2]), .ZN(n9) );
  ND2D1BWP30P140LVT U16 ( .A1(n1), .A2(i_data_bus[34]), .ZN(n10) );
  ND2OPTIBD1BWP30P140LVT U17 ( .A1(n12), .A2(n11), .ZN(N95) );
  ND2OPTIBD1BWP30P140LVT U18 ( .A1(n69), .A2(i_data_bus[3]), .ZN(n11) );
  ND2D1BWP30P140LVT U19 ( .A1(n71), .A2(i_data_bus[35]), .ZN(n12) );
  ND2OPTIBD1BWP30P140LVT U20 ( .A1(n14), .A2(n13), .ZN(N96) );
  ND2OPTIBD1BWP30P140LVT U21 ( .A1(n69), .A2(i_data_bus[4]), .ZN(n13) );
  ND2D1BWP30P140LVT U22 ( .A1(n1), .A2(i_data_bus[36]), .ZN(n14) );
  ND2OPTIBD1BWP30P140LVT U23 ( .A1(n16), .A2(n15), .ZN(N97) );
  ND2OPTIBD1BWP30P140LVT U24 ( .A1(n69), .A2(i_data_bus[5]), .ZN(n15) );
  ND2D1BWP30P140LVT U25 ( .A1(n71), .A2(i_data_bus[37]), .ZN(n16) );
  ND2OPTIBD1BWP30P140LVT U26 ( .A1(n18), .A2(n17), .ZN(N98) );
  ND2OPTIBD1BWP30P140LVT U27 ( .A1(n69), .A2(i_data_bus[6]), .ZN(n17) );
  ND2D1BWP30P140LVT U28 ( .A1(n1), .A2(i_data_bus[38]), .ZN(n18) );
  ND2OPTIBD1BWP30P140LVT U29 ( .A1(n20), .A2(n19), .ZN(N99) );
  ND2OPTIBD1BWP30P140LVT U30 ( .A1(n69), .A2(i_data_bus[7]), .ZN(n19) );
  ND2D1BWP30P140LVT U31 ( .A1(n71), .A2(i_data_bus[39]), .ZN(n20) );
  ND2OPTIBD1BWP30P140LVT U32 ( .A1(n22), .A2(n21), .ZN(N100) );
  ND2OPTIBD1BWP30P140LVT U33 ( .A1(n69), .A2(i_data_bus[8]), .ZN(n21) );
  ND2D1BWP30P140LVT U34 ( .A1(n1), .A2(i_data_bus[40]), .ZN(n22) );
  ND2OPTIBD1BWP30P140LVT U35 ( .A1(n24), .A2(n23), .ZN(N101) );
  ND2OPTIBD1BWP30P140LVT U36 ( .A1(n69), .A2(i_data_bus[9]), .ZN(n23) );
  ND2D1BWP30P140LVT U37 ( .A1(n71), .A2(i_data_bus[41]), .ZN(n24) );
  ND2OPTIBD1BWP30P140LVT U38 ( .A1(n26), .A2(n25), .ZN(N102) );
  ND2OPTIBD1BWP30P140LVT U39 ( .A1(n69), .A2(i_data_bus[10]), .ZN(n25) );
  ND2D1BWP30P140LVT U40 ( .A1(n1), .A2(i_data_bus[42]), .ZN(n26) );
  ND2OPTIBD1BWP30P140LVT U41 ( .A1(n28), .A2(n27), .ZN(N103) );
  ND2OPTIBD1BWP30P140LVT U42 ( .A1(n69), .A2(i_data_bus[11]), .ZN(n27) );
  ND2D1BWP30P140LVT U43 ( .A1(n71), .A2(i_data_bus[43]), .ZN(n28) );
  ND2OPTIBD1BWP30P140LVT U44 ( .A1(n30), .A2(n29), .ZN(N104) );
  ND2OPTIBD1BWP30P140LVT U45 ( .A1(n69), .A2(i_data_bus[12]), .ZN(n29) );
  ND2D1BWP30P140LVT U46 ( .A1(n1), .A2(i_data_bus[44]), .ZN(n30) );
  ND2OPTIBD1BWP30P140LVT U47 ( .A1(n32), .A2(n31), .ZN(N105) );
  ND2OPTIBD1BWP30P140LVT U48 ( .A1(n69), .A2(i_data_bus[13]), .ZN(n31) );
  ND2D1BWP30P140LVT U49 ( .A1(n71), .A2(i_data_bus[45]), .ZN(n32) );
  ND2OPTIBD1BWP30P140LVT U50 ( .A1(n34), .A2(n33), .ZN(N106) );
  ND2OPTIBD1BWP30P140LVT U51 ( .A1(n69), .A2(i_data_bus[14]), .ZN(n33) );
  ND2D1BWP30P140LVT U52 ( .A1(n1), .A2(i_data_bus[46]), .ZN(n34) );
  ND2OPTIBD1BWP30P140LVT U53 ( .A1(n36), .A2(n35), .ZN(N107) );
  ND2OPTIBD1BWP30P140LVT U54 ( .A1(n69), .A2(i_data_bus[15]), .ZN(n35) );
  ND2D1BWP30P140LVT U55 ( .A1(n71), .A2(i_data_bus[47]), .ZN(n36) );
  ND2OPTIBD1BWP30P140LVT U56 ( .A1(n38), .A2(n37), .ZN(N108) );
  ND2OPTIBD1BWP30P140LVT U57 ( .A1(n69), .A2(i_data_bus[16]), .ZN(n37) );
  ND2D1BWP30P140LVT U58 ( .A1(n1), .A2(i_data_bus[48]), .ZN(n38) );
  ND2OPTIBD1BWP30P140LVT U59 ( .A1(n40), .A2(n39), .ZN(N109) );
  ND2OPTIBD1BWP30P140LVT U60 ( .A1(n69), .A2(i_data_bus[17]), .ZN(n39) );
  ND2D1BWP30P140LVT U61 ( .A1(n71), .A2(i_data_bus[49]), .ZN(n40) );
  ND2OPTIBD1BWP30P140LVT U62 ( .A1(n42), .A2(n41), .ZN(N110) );
  ND2OPTIBD1BWP30P140LVT U63 ( .A1(n69), .A2(i_data_bus[18]), .ZN(n41) );
  ND2D1BWP30P140LVT U64 ( .A1(n1), .A2(i_data_bus[50]), .ZN(n42) );
  ND2OPTIBD1BWP30P140LVT U65 ( .A1(n44), .A2(n43), .ZN(N111) );
  ND2OPTIBD1BWP30P140LVT U66 ( .A1(n69), .A2(i_data_bus[19]), .ZN(n43) );
  ND2D1BWP30P140LVT U67 ( .A1(n71), .A2(i_data_bus[51]), .ZN(n44) );
  ND2OPTIBD1BWP30P140LVT U68 ( .A1(n46), .A2(n45), .ZN(N112) );
  ND2OPTIBD1BWP30P140LVT U69 ( .A1(n69), .A2(i_data_bus[20]), .ZN(n45) );
  ND2D1BWP30P140LVT U70 ( .A1(n1), .A2(i_data_bus[52]), .ZN(n46) );
  ND2OPTIBD1BWP30P140LVT U71 ( .A1(n48), .A2(n47), .ZN(N113) );
  ND2OPTIBD1BWP30P140LVT U72 ( .A1(n69), .A2(i_data_bus[21]), .ZN(n47) );
  ND2D1BWP30P140LVT U73 ( .A1(n71), .A2(i_data_bus[53]), .ZN(n48) );
  ND2OPTIBD1BWP30P140LVT U74 ( .A1(n50), .A2(n49), .ZN(N114) );
  ND2OPTIBD1BWP30P140LVT U75 ( .A1(n69), .A2(i_data_bus[22]), .ZN(n49) );
  ND2D1BWP30P140LVT U76 ( .A1(n1), .A2(i_data_bus[54]), .ZN(n50) );
  ND2OPTIBD1BWP30P140LVT U77 ( .A1(n52), .A2(n51), .ZN(N115) );
  ND2OPTIBD1BWP30P140LVT U78 ( .A1(n69), .A2(i_data_bus[23]), .ZN(n51) );
  ND2D1BWP30P140LVT U79 ( .A1(n71), .A2(i_data_bus[55]), .ZN(n52) );
  ND2OPTIBD1BWP30P140LVT U80 ( .A1(n54), .A2(n53), .ZN(N116) );
  ND2OPTIBD1BWP30P140LVT U81 ( .A1(n69), .A2(i_data_bus[24]), .ZN(n53) );
  ND2D1BWP30P140LVT U82 ( .A1(n1), .A2(i_data_bus[56]), .ZN(n54) );
  ND2OPTIBD1BWP30P140LVT U83 ( .A1(n56), .A2(n55), .ZN(N117) );
  ND2OPTIBD1BWP30P140LVT U84 ( .A1(n69), .A2(i_data_bus[25]), .ZN(n55) );
  ND2D1BWP30P140LVT U85 ( .A1(n71), .A2(i_data_bus[57]), .ZN(n56) );
  ND2OPTIBD1BWP30P140LVT U86 ( .A1(n58), .A2(n57), .ZN(N118) );
  ND2OPTIBD1BWP30P140LVT U87 ( .A1(n69), .A2(i_data_bus[26]), .ZN(n57) );
  ND2D1BWP30P140LVT U88 ( .A1(n1), .A2(i_data_bus[58]), .ZN(n58) );
  ND2OPTIBD1BWP30P140LVT U89 ( .A1(n60), .A2(n59), .ZN(N119) );
  ND2OPTIBD1BWP30P140LVT U90 ( .A1(n69), .A2(i_data_bus[27]), .ZN(n59) );
  ND2D1BWP30P140LVT U91 ( .A1(n71), .A2(i_data_bus[59]), .ZN(n60) );
  ND2OPTIBD1BWP30P140LVT U92 ( .A1(n62), .A2(n61), .ZN(N120) );
  ND2OPTIBD1BWP30P140LVT U93 ( .A1(n69), .A2(i_data_bus[28]), .ZN(n61) );
  ND2D1BWP30P140LVT U94 ( .A1(n1), .A2(i_data_bus[60]), .ZN(n62) );
  ND2OPTIBD1BWP30P140LVT U95 ( .A1(n64), .A2(n63), .ZN(N121) );
  ND2OPTIBD1BWP30P140LVT U96 ( .A1(n69), .A2(i_data_bus[29]), .ZN(n63) );
  ND2D1BWP30P140LVT U97 ( .A1(n71), .A2(i_data_bus[61]), .ZN(n64) );
  ND2OPTIBD1BWP30P140LVT U98 ( .A1(n66), .A2(n65), .ZN(N122) );
  ND2OPTIBD1BWP30P140LVT U99 ( .A1(n69), .A2(i_data_bus[30]), .ZN(n65) );
  ND2D1BWP30P140LVT U100 ( .A1(n1), .A2(i_data_bus[62]), .ZN(n66) );
  ND2OPTIBD1BWP30P140LVT U101 ( .A1(n68), .A2(n67), .ZN(N123) );
  ND2OPTIBD1BWP30P140LVT U102 ( .A1(n69), .A2(i_data_bus[31]), .ZN(n67) );
  ND2D1BWP30P140LVT U103 ( .A1(n71), .A2(i_data_bus[63]), .ZN(n68) );
  IND2D1BWP30P140LVT U104 ( .A1(n71), .B1(n70), .ZN(N91) );
  INVD1BWP30P140LVT U105 ( .I(n69), .ZN(n70) );
  ND3D1BWP30P140LVT U106 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2)
         );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_30 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_30 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_5 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_30 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_29 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_28 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_27 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_26 o_data_high ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_25 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_31 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n4), .A2(n3), .ZN(n2) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n4) );
  INVD1BWP30P140LVT U5 ( .I(n7), .ZN(n8) );
  NR2D1BWP30P140LVT U6 ( .A1(n4), .A2(n3), .ZN(n1) );
  INVD1BWP30P140LVT U7 ( .I(n8), .ZN(n36) );
  INVD1BWP30P140LVT U8 ( .I(n8), .ZN(n41) );
  OR2D1BWP30P140LVT U9 ( .A1(rst), .A2(i_cmd[0]), .Z(n3) );
  ND3D1BWP30P140LVT U10 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n6)
         );
  INVD1BWP30P140LVT U11 ( .I(rst), .ZN(n5) );
  IND2D1BWP30P140LVT U12 ( .A1(n6), .B1(n5), .ZN(n7) );
  IND2D1BWP30P140LVT U13 ( .A1(n2), .B1(n41), .ZN(N91) );
  INVD1BWP30P140LVT U14 ( .I(i_data_bus[52]), .ZN(n9) );
  MOAI22D1BWP30P140LVT U15 ( .A1(n9), .A2(n36), .B1(i_data_bus[20]), .B2(n2), 
        .ZN(N112) );
  INVD1BWP30P140LVT U16 ( .I(i_data_bus[54]), .ZN(n10) );
  MOAI22D1BWP30P140LVT U17 ( .A1(n10), .A2(n36), .B1(i_data_bus[22]), .B2(n1), 
        .ZN(N114) );
  INVD1BWP30P140LVT U18 ( .I(i_data_bus[48]), .ZN(n11) );
  MOAI22D1BWP30P140LVT U19 ( .A1(n11), .A2(n36), .B1(i_data_bus[16]), .B2(n2), 
        .ZN(N108) );
  INVD1BWP30P140LVT U20 ( .I(i_data_bus[50]), .ZN(n12) );
  MOAI22D1BWP30P140LVT U21 ( .A1(n12), .A2(n36), .B1(i_data_bus[18]), .B2(n1), 
        .ZN(N110) );
  INVD1BWP30P140LVT U22 ( .I(i_data_bus[32]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U23 ( .A1(n13), .A2(n41), .B1(i_data_bus[0]), .B2(n2), 
        .ZN(N92) );
  INVD1BWP30P140LVT U24 ( .I(i_data_bus[33]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U25 ( .A1(n14), .A2(n41), .B1(i_data_bus[1]), .B2(n1), 
        .ZN(N93) );
  INVD1BWP30P140LVT U26 ( .I(i_data_bus[34]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U27 ( .A1(n15), .A2(n41), .B1(i_data_bus[2]), .B2(n2), 
        .ZN(N94) );
  INVD1BWP30P140LVT U28 ( .I(i_data_bus[35]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U29 ( .A1(n16), .A2(n41), .B1(i_data_bus[3]), .B2(n1), 
        .ZN(N95) );
  INVD1BWP30P140LVT U30 ( .I(i_data_bus[36]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U31 ( .A1(n17), .A2(n41), .B1(i_data_bus[4]), .B2(n2), 
        .ZN(N96) );
  INVD1BWP30P140LVT U32 ( .I(i_data_bus[37]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U33 ( .A1(n18), .A2(n41), .B1(i_data_bus[5]), .B2(n1), 
        .ZN(N97) );
  INVD1BWP30P140LVT U34 ( .I(i_data_bus[38]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U35 ( .A1(n19), .A2(n41), .B1(i_data_bus[6]), .B2(n2), 
        .ZN(N98) );
  INVD1BWP30P140LVT U36 ( .I(i_data_bus[39]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U37 ( .A1(n20), .A2(n41), .B1(i_data_bus[7]), .B2(n1), 
        .ZN(N99) );
  INVD1BWP30P140LVT U38 ( .I(i_data_bus[40]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U39 ( .A1(n21), .A2(n41), .B1(i_data_bus[8]), .B2(n2), 
        .ZN(N100) );
  INVD1BWP30P140LVT U40 ( .I(i_data_bus[41]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U41 ( .A1(n22), .A2(n41), .B1(i_data_bus[9]), .B2(n1), 
        .ZN(N101) );
  INVD1BWP30P140LVT U42 ( .I(i_data_bus[42]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U43 ( .A1(n23), .A2(n41), .B1(i_data_bus[10]), .B2(n2), 
        .ZN(N102) );
  INVD1BWP30P140LVT U44 ( .I(i_data_bus[43]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U45 ( .A1(n24), .A2(n41), .B1(i_data_bus[11]), .B2(n1), 
        .ZN(N103) );
  INVD1BWP30P140LVT U46 ( .I(i_data_bus[47]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U47 ( .A1(n25), .A2(n36), .B1(i_data_bus[15]), .B2(n1), 
        .ZN(N107) );
  INVD1BWP30P140LVT U48 ( .I(i_data_bus[44]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U49 ( .A1(n26), .A2(n36), .B1(i_data_bus[12]), .B2(n2), 
        .ZN(N104) );
  INVD1BWP30P140LVT U50 ( .I(i_data_bus[55]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U51 ( .A1(n27), .A2(n36), .B1(i_data_bus[23]), .B2(n1), 
        .ZN(N115) );
  INVD1BWP30P140LVT U52 ( .I(i_data_bus[61]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U53 ( .A1(n28), .A2(n36), .B1(i_data_bus[29]), .B2(n2), 
        .ZN(N121) );
  INVD1BWP30P140LVT U54 ( .I(i_data_bus[46]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U55 ( .A1(n29), .A2(n36), .B1(i_data_bus[14]), .B2(n1), 
        .ZN(N106) );
  INVD1BWP30P140LVT U56 ( .I(i_data_bus[59]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U57 ( .A1(n30), .A2(n36), .B1(i_data_bus[27]), .B2(n2), 
        .ZN(N119) );
  INVD1BWP30P140LVT U58 ( .I(i_data_bus[45]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U59 ( .A1(n31), .A2(n36), .B1(i_data_bus[13]), .B2(n1), 
        .ZN(N105) );
  INVD1BWP30P140LVT U60 ( .I(i_data_bus[51]), .ZN(n32) );
  MOAI22D1BWP30P140LVT U61 ( .A1(n32), .A2(n36), .B1(i_data_bus[19]), .B2(n2), 
        .ZN(N111) );
  INVD1BWP30P140LVT U62 ( .I(i_data_bus[57]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U63 ( .A1(n33), .A2(n36), .B1(i_data_bus[25]), .B2(n1), 
        .ZN(N117) );
  INVD1BWP30P140LVT U64 ( .I(i_data_bus[49]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U65 ( .A1(n34), .A2(n36), .B1(i_data_bus[17]), .B2(n2), 
        .ZN(N109) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[63]), .ZN(n35) );
  MOAI22D1BWP30P140LVT U67 ( .A1(n35), .A2(n36), .B1(i_data_bus[31]), .B2(n1), 
        .ZN(N123) );
  INVD1BWP30P140LVT U68 ( .I(i_data_bus[53]), .ZN(n37) );
  MOAI22D1BWP30P140LVT U69 ( .A1(n37), .A2(n36), .B1(i_data_bus[21]), .B2(n2), 
        .ZN(N113) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[56]), .ZN(n38) );
  MOAI22D1BWP30P140LVT U71 ( .A1(n38), .A2(n41), .B1(i_data_bus[24]), .B2(n1), 
        .ZN(N116) );
  INVD1BWP30P140LVT U72 ( .I(i_data_bus[60]), .ZN(n39) );
  MOAI22D1BWP30P140LVT U73 ( .A1(n39), .A2(n41), .B1(i_data_bus[28]), .B2(n2), 
        .ZN(N120) );
  INVD1BWP30P140LVT U74 ( .I(i_data_bus[62]), .ZN(n40) );
  MOAI22D1BWP30P140LVT U75 ( .A1(n40), .A2(n41), .B1(i_data_bus[30]), .B2(n1), 
        .ZN(N122) );
  INVD1BWP30P140LVT U76 ( .I(i_data_bus[58]), .ZN(n42) );
  MOAI22D1BWP30P140LVT U77 ( .A1(n42), .A2(n41), .B1(i_data_bus[26]), .B2(n2), 
        .ZN(N118) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_31 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_31 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_32 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n4), .A2(n3), .ZN(n2) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n4) );
  INVD1BWP30P140LVT U5 ( .I(n7), .ZN(n8) );
  NR2D1BWP30P140LVT U6 ( .A1(n4), .A2(n3), .ZN(n1) );
  INVD1BWP30P140LVT U7 ( .I(n8), .ZN(n36) );
  INVD1BWP30P140LVT U8 ( .I(n8), .ZN(n41) );
  OR2D1BWP30P140LVT U9 ( .A1(rst), .A2(i_cmd[0]), .Z(n3) );
  ND3D1BWP30P140LVT U10 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n6)
         );
  INVD1BWP30P140LVT U11 ( .I(rst), .ZN(n5) );
  IND2D1BWP30P140LVT U12 ( .A1(n6), .B1(n5), .ZN(n7) );
  IND2D1BWP30P140LVT U13 ( .A1(n2), .B1(n41), .ZN(N91) );
  INVD1BWP30P140LVT U14 ( .I(i_data_bus[48]), .ZN(n9) );
  MOAI22D1BWP30P140LVT U15 ( .A1(n9), .A2(n36), .B1(i_data_bus[16]), .B2(n2), 
        .ZN(N108) );
  INVD1BWP30P140LVT U16 ( .I(i_data_bus[52]), .ZN(n10) );
  MOAI22D1BWP30P140LVT U17 ( .A1(n10), .A2(n36), .B1(i_data_bus[20]), .B2(n1), 
        .ZN(N112) );
  INVD1BWP30P140LVT U18 ( .I(i_data_bus[50]), .ZN(n11) );
  MOAI22D1BWP30P140LVT U19 ( .A1(n11), .A2(n36), .B1(i_data_bus[18]), .B2(n2), 
        .ZN(N110) );
  INVD1BWP30P140LVT U20 ( .I(i_data_bus[54]), .ZN(n12) );
  MOAI22D1BWP30P140LVT U21 ( .A1(n12), .A2(n36), .B1(i_data_bus[22]), .B2(n1), 
        .ZN(N114) );
  INVD1BWP30P140LVT U22 ( .I(i_data_bus[37]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U23 ( .A1(n13), .A2(n41), .B1(i_data_bus[5]), .B2(n2), 
        .ZN(N97) );
  INVD1BWP30P140LVT U24 ( .I(i_data_bus[36]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U25 ( .A1(n14), .A2(n41), .B1(i_data_bus[4]), .B2(n1), 
        .ZN(N96) );
  INVD1BWP30P140LVT U26 ( .I(i_data_bus[34]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U27 ( .A1(n15), .A2(n41), .B1(i_data_bus[2]), .B2(n2), 
        .ZN(N94) );
  INVD1BWP30P140LVT U28 ( .I(i_data_bus[40]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U29 ( .A1(n16), .A2(n41), .B1(i_data_bus[8]), .B2(n1), 
        .ZN(N100) );
  INVD1BWP30P140LVT U30 ( .I(i_data_bus[43]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U31 ( .A1(n17), .A2(n41), .B1(i_data_bus[11]), .B2(n2), 
        .ZN(N103) );
  INVD1BWP30P140LVT U32 ( .I(i_data_bus[38]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U33 ( .A1(n18), .A2(n41), .B1(i_data_bus[6]), .B2(n1), 
        .ZN(N98) );
  INVD1BWP30P140LVT U34 ( .I(i_data_bus[33]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U35 ( .A1(n19), .A2(n41), .B1(i_data_bus[1]), .B2(n2), 
        .ZN(N93) );
  INVD1BWP30P140LVT U36 ( .I(i_data_bus[39]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U37 ( .A1(n20), .A2(n41), .B1(i_data_bus[7]), .B2(n1), 
        .ZN(N99) );
  INVD1BWP30P140LVT U38 ( .I(i_data_bus[41]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U39 ( .A1(n21), .A2(n41), .B1(i_data_bus[9]), .B2(n2), 
        .ZN(N101) );
  INVD1BWP30P140LVT U40 ( .I(i_data_bus[32]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U41 ( .A1(n22), .A2(n41), .B1(i_data_bus[0]), .B2(n1), 
        .ZN(N92) );
  INVD1BWP30P140LVT U42 ( .I(i_data_bus[35]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U43 ( .A1(n23), .A2(n41), .B1(i_data_bus[3]), .B2(n2), 
        .ZN(N95) );
  INVD1BWP30P140LVT U44 ( .I(i_data_bus[42]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U45 ( .A1(n24), .A2(n41), .B1(i_data_bus[10]), .B2(n1), 
        .ZN(N102) );
  INVD1BWP30P140LVT U46 ( .I(i_data_bus[55]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U47 ( .A1(n25), .A2(n36), .B1(i_data_bus[23]), .B2(n1), 
        .ZN(N115) );
  INVD1BWP30P140LVT U48 ( .I(i_data_bus[53]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U49 ( .A1(n26), .A2(n36), .B1(i_data_bus[21]), .B2(n2), 
        .ZN(N113) );
  INVD1BWP30P140LVT U50 ( .I(i_data_bus[51]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U51 ( .A1(n27), .A2(n36), .B1(i_data_bus[19]), .B2(n1), 
        .ZN(N111) );
  INVD1BWP30P140LVT U52 ( .I(i_data_bus[49]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U53 ( .A1(n28), .A2(n36), .B1(i_data_bus[17]), .B2(n2), 
        .ZN(N109) );
  INVD1BWP30P140LVT U54 ( .I(i_data_bus[46]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U55 ( .A1(n29), .A2(n36), .B1(i_data_bus[14]), .B2(n1), 
        .ZN(N106) );
  INVD1BWP30P140LVT U56 ( .I(i_data_bus[45]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U57 ( .A1(n30), .A2(n36), .B1(i_data_bus[13]), .B2(n2), 
        .ZN(N105) );
  INVD1BWP30P140LVT U58 ( .I(i_data_bus[44]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U59 ( .A1(n31), .A2(n36), .B1(i_data_bus[12]), .B2(n1), 
        .ZN(N104) );
  INVD1BWP30P140LVT U60 ( .I(i_data_bus[63]), .ZN(n32) );
  MOAI22D1BWP30P140LVT U61 ( .A1(n32), .A2(n36), .B1(i_data_bus[31]), .B2(n2), 
        .ZN(N123) );
  INVD1BWP30P140LVT U62 ( .I(i_data_bus[61]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U63 ( .A1(n33), .A2(n36), .B1(i_data_bus[29]), .B2(n1), 
        .ZN(N121) );
  INVD1BWP30P140LVT U64 ( .I(i_data_bus[59]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U65 ( .A1(n34), .A2(n36), .B1(i_data_bus[27]), .B2(n2), 
        .ZN(N119) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[57]), .ZN(n35) );
  MOAI22D1BWP30P140LVT U67 ( .A1(n35), .A2(n36), .B1(i_data_bus[25]), .B2(n1), 
        .ZN(N117) );
  INVD1BWP30P140LVT U68 ( .I(i_data_bus[47]), .ZN(n37) );
  MOAI22D1BWP30P140LVT U69 ( .A1(n37), .A2(n36), .B1(i_data_bus[15]), .B2(n2), 
        .ZN(N107) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[60]), .ZN(n38) );
  MOAI22D1BWP30P140LVT U71 ( .A1(n38), .A2(n41), .B1(i_data_bus[28]), .B2(n1), 
        .ZN(N120) );
  INVD1BWP30P140LVT U72 ( .I(i_data_bus[62]), .ZN(n39) );
  MOAI22D1BWP30P140LVT U73 ( .A1(n39), .A2(n41), .B1(i_data_bus[30]), .B2(n2), 
        .ZN(N122) );
  INVD1BWP30P140LVT U74 ( .I(i_data_bus[56]), .ZN(n40) );
  MOAI22D1BWP30P140LVT U75 ( .A1(n40), .A2(n41), .B1(i_data_bus[24]), .B2(n1), 
        .ZN(N116) );
  INVD1BWP30P140LVT U76 ( .I(i_data_bus[58]), .ZN(n42) );
  MOAI22D1BWP30P140LVT U77 ( .A1(n42), .A2(n41), .B1(i_data_bus[26]), .B2(n2), 
        .ZN(N118) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_32 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_32 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_33 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U36 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_33 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_33 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_34 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  IND2D1BWP30P140LVT U3 ( .A1(n1), .B1(i_valid[0]), .ZN(n2) );
  INVD1BWP30P140LVT U4 ( .I(i_en), .ZN(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  NR3D1P5BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n6) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  BUFFD2BWP30P140LVT U8 ( .I(n4), .Z(n5) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n5), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n5), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n5), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n5), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n5), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n5), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n5), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n5), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n5), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n5), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n5), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n5), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n5), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n5), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n5), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n5), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n5), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n5), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n5), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n5), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n5), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n5), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n5), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n5), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n5), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n5), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n5), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n5), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n5), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n5), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n5), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n5), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n5), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_34 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_34 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_35 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3OPTPAD2BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  NR2D1BWP30P140LVT U4 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U5 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U8 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_35 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_35 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_36 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3OPTPAD2BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  NR2D1BWP30P140LVT U4 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U5 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U8 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_36 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_36 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_6 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_36 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_35 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_34 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_33 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_32 o_data_high ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_31 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_37 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n4), .A2(n3), .ZN(n2) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n4) );
  INVD1BWP30P140LVT U5 ( .I(n7), .ZN(n8) );
  IND2D1BWP30P140LVT U6 ( .A1(n6), .B1(n5), .ZN(n7) );
  NR2D1BWP30P140LVT U7 ( .A1(n4), .A2(n3), .ZN(n1) );
  INVD1BWP30P140LVT U8 ( .I(n8), .ZN(n36) );
  INVD1BWP30P140LVT U9 ( .I(n8), .ZN(n41) );
  OR2D1BWP30P140LVT U10 ( .A1(rst), .A2(i_cmd[0]), .Z(n3) );
  ND3D1BWP30P140LVT U11 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n6)
         );
  INVD1BWP30P140LVT U12 ( .I(rst), .ZN(n5) );
  IND2D1BWP30P140LVT U13 ( .A1(n2), .B1(n41), .ZN(N91) );
  INVD1BWP30P140LVT U14 ( .I(i_data_bus[54]), .ZN(n9) );
  MOAI22D1BWP30P140LVT U15 ( .A1(n9), .A2(n36), .B1(i_data_bus[22]), .B2(n2), 
        .ZN(N114) );
  INVD1BWP30P140LVT U16 ( .I(i_data_bus[50]), .ZN(n10) );
  MOAI22D1BWP30P140LVT U17 ( .A1(n10), .A2(n36), .B1(i_data_bus[18]), .B2(n1), 
        .ZN(N110) );
  INVD1BWP30P140LVT U18 ( .I(i_data_bus[48]), .ZN(n11) );
  MOAI22D1BWP30P140LVT U19 ( .A1(n11), .A2(n36), .B1(i_data_bus[16]), .B2(n2), 
        .ZN(N108) );
  INVD1BWP30P140LVT U20 ( .I(i_data_bus[52]), .ZN(n12) );
  MOAI22D1BWP30P140LVT U21 ( .A1(n12), .A2(n36), .B1(i_data_bus[20]), .B2(n1), 
        .ZN(N112) );
  INVD1BWP30P140LVT U22 ( .I(i_data_bus[38]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U23 ( .A1(n13), .A2(n41), .B1(i_data_bus[6]), .B2(n2), 
        .ZN(N98) );
  INVD1BWP30P140LVT U24 ( .I(i_data_bus[39]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U25 ( .A1(n14), .A2(n41), .B1(i_data_bus[7]), .B2(n1), 
        .ZN(N99) );
  INVD1BWP30P140LVT U26 ( .I(i_data_bus[40]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U27 ( .A1(n15), .A2(n41), .B1(i_data_bus[8]), .B2(n2), 
        .ZN(N100) );
  INVD1BWP30P140LVT U28 ( .I(i_data_bus[41]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U29 ( .A1(n16), .A2(n41), .B1(i_data_bus[9]), .B2(n1), 
        .ZN(N101) );
  INVD1BWP30P140LVT U30 ( .I(i_data_bus[42]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U31 ( .A1(n17), .A2(n41), .B1(i_data_bus[10]), .B2(n2), 
        .ZN(N102) );
  INVD1BWP30P140LVT U32 ( .I(i_data_bus[43]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U33 ( .A1(n18), .A2(n41), .B1(i_data_bus[11]), .B2(n1), 
        .ZN(N103) );
  INVD1BWP30P140LVT U34 ( .I(i_data_bus[35]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U35 ( .A1(n19), .A2(n41), .B1(i_data_bus[3]), .B2(n2), 
        .ZN(N95) );
  INVD1BWP30P140LVT U36 ( .I(i_data_bus[32]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U37 ( .A1(n20), .A2(n41), .B1(i_data_bus[0]), .B2(n1), 
        .ZN(N92) );
  INVD1BWP30P140LVT U38 ( .I(i_data_bus[33]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U39 ( .A1(n21), .A2(n41), .B1(i_data_bus[1]), .B2(n2), 
        .ZN(N93) );
  INVD1BWP30P140LVT U40 ( .I(i_data_bus[34]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U41 ( .A1(n22), .A2(n41), .B1(i_data_bus[2]), .B2(n1), 
        .ZN(N94) );
  INVD1BWP30P140LVT U42 ( .I(i_data_bus[36]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U43 ( .A1(n23), .A2(n41), .B1(i_data_bus[4]), .B2(n2), 
        .ZN(N96) );
  INVD1BWP30P140LVT U44 ( .I(i_data_bus[37]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U45 ( .A1(n24), .A2(n41), .B1(i_data_bus[5]), .B2(n1), 
        .ZN(N97) );
  INVD1BWP30P140LVT U46 ( .I(i_data_bus[46]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U47 ( .A1(n25), .A2(n36), .B1(i_data_bus[14]), .B2(n1), 
        .ZN(N106) );
  INVD1BWP30P140LVT U48 ( .I(i_data_bus[61]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U49 ( .A1(n26), .A2(n36), .B1(i_data_bus[29]), .B2(n2), 
        .ZN(N121) );
  INVD1BWP30P140LVT U50 ( .I(i_data_bus[45]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U51 ( .A1(n27), .A2(n36), .B1(i_data_bus[13]), .B2(n1), 
        .ZN(N105) );
  INVD1BWP30P140LVT U52 ( .I(i_data_bus[44]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U53 ( .A1(n28), .A2(n36), .B1(i_data_bus[12]), .B2(n2), 
        .ZN(N104) );
  INVD1BWP30P140LVT U54 ( .I(i_data_bus[51]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U55 ( .A1(n29), .A2(n36), .B1(i_data_bus[19]), .B2(n1), 
        .ZN(N111) );
  INVD1BWP30P140LVT U56 ( .I(i_data_bus[63]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U57 ( .A1(n30), .A2(n36), .B1(i_data_bus[31]), .B2(n2), 
        .ZN(N123) );
  INVD1BWP30P140LVT U58 ( .I(i_data_bus[49]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U59 ( .A1(n31), .A2(n36), .B1(i_data_bus[17]), .B2(n1), 
        .ZN(N109) );
  INVD1BWP30P140LVT U60 ( .I(i_data_bus[59]), .ZN(n32) );
  MOAI22D1BWP30P140LVT U61 ( .A1(n32), .A2(n36), .B1(i_data_bus[27]), .B2(n2), 
        .ZN(N119) );
  INVD1BWP30P140LVT U62 ( .I(i_data_bus[53]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U63 ( .A1(n33), .A2(n36), .B1(i_data_bus[21]), .B2(n1), 
        .ZN(N113) );
  INVD1BWP30P140LVT U64 ( .I(i_data_bus[57]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U65 ( .A1(n34), .A2(n36), .B1(i_data_bus[25]), .B2(n2), 
        .ZN(N117) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[47]), .ZN(n35) );
  MOAI22D1BWP30P140LVT U67 ( .A1(n35), .A2(n36), .B1(i_data_bus[15]), .B2(n1), 
        .ZN(N107) );
  INVD1BWP30P140LVT U68 ( .I(i_data_bus[55]), .ZN(n37) );
  MOAI22D1BWP30P140LVT U69 ( .A1(n37), .A2(n36), .B1(i_data_bus[23]), .B2(n2), 
        .ZN(N115) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[58]), .ZN(n38) );
  MOAI22D1BWP30P140LVT U71 ( .A1(n38), .A2(n41), .B1(i_data_bus[26]), .B2(n1), 
        .ZN(N118) );
  INVD1BWP30P140LVT U72 ( .I(i_data_bus[60]), .ZN(n39) );
  MOAI22D1BWP30P140LVT U73 ( .A1(n39), .A2(n41), .B1(i_data_bus[28]), .B2(n2), 
        .ZN(N120) );
  INVD1BWP30P140LVT U74 ( .I(i_data_bus[62]), .ZN(n40) );
  MOAI22D1BWP30P140LVT U75 ( .A1(n40), .A2(n41), .B1(i_data_bus[30]), .B2(n1), 
        .ZN(N122) );
  INVD1BWP30P140LVT U76 ( .I(i_data_bus[56]), .ZN(n42) );
  MOAI22D1BWP30P140LVT U77 ( .A1(n42), .A2(n41), .B1(i_data_bus[24]), .B2(n2), 
        .ZN(N116) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_37 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_37 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_38 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n4), .A2(n3), .ZN(n2) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n4) );
  INVD1BWP30P140LVT U5 ( .I(n7), .ZN(n8) );
  IND2D1BWP30P140LVT U6 ( .A1(n6), .B1(n5), .ZN(n7) );
  NR2D1BWP30P140LVT U7 ( .A1(n4), .A2(n3), .ZN(n1) );
  INVD1BWP30P140LVT U8 ( .I(n8), .ZN(n36) );
  INVD1BWP30P140LVT U9 ( .I(n8), .ZN(n41) );
  OR2D1BWP30P140LVT U10 ( .A1(rst), .A2(i_cmd[0]), .Z(n3) );
  ND3D1BWP30P140LVT U11 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n6)
         );
  INVD1BWP30P140LVT U12 ( .I(rst), .ZN(n5) );
  IND2D1BWP30P140LVT U13 ( .A1(n2), .B1(n41), .ZN(N91) );
  INVD1BWP30P140LVT U14 ( .I(i_data_bus[54]), .ZN(n9) );
  MOAI22D1BWP30P140LVT U15 ( .A1(n9), .A2(n36), .B1(i_data_bus[22]), .B2(n2), 
        .ZN(N114) );
  INVD1BWP30P140LVT U16 ( .I(i_data_bus[50]), .ZN(n10) );
  MOAI22D1BWP30P140LVT U17 ( .A1(n10), .A2(n36), .B1(i_data_bus[18]), .B2(n1), 
        .ZN(N110) );
  INVD1BWP30P140LVT U18 ( .I(i_data_bus[52]), .ZN(n11) );
  MOAI22D1BWP30P140LVT U19 ( .A1(n11), .A2(n36), .B1(i_data_bus[20]), .B2(n2), 
        .ZN(N112) );
  INVD1BWP30P140LVT U20 ( .I(i_data_bus[48]), .ZN(n12) );
  MOAI22D1BWP30P140LVT U21 ( .A1(n12), .A2(n36), .B1(i_data_bus[16]), .B2(n1), 
        .ZN(N108) );
  INVD1BWP30P140LVT U22 ( .I(i_data_bus[42]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U23 ( .A1(n13), .A2(n41), .B1(i_data_bus[10]), .B2(n2), 
        .ZN(N102) );
  INVD1BWP30P140LVT U24 ( .I(i_data_bus[41]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U25 ( .A1(n14), .A2(n41), .B1(i_data_bus[9]), .B2(n1), 
        .ZN(N101) );
  INVD1BWP30P140LVT U26 ( .I(i_data_bus[32]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U27 ( .A1(n15), .A2(n41), .B1(i_data_bus[0]), .B2(n2), 
        .ZN(N92) );
  INVD1BWP30P140LVT U28 ( .I(i_data_bus[33]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U29 ( .A1(n16), .A2(n41), .B1(i_data_bus[1]), .B2(n1), 
        .ZN(N93) );
  INVD1BWP30P140LVT U30 ( .I(i_data_bus[34]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U31 ( .A1(n17), .A2(n41), .B1(i_data_bus[2]), .B2(n2), 
        .ZN(N94) );
  INVD1BWP30P140LVT U32 ( .I(i_data_bus[43]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U33 ( .A1(n18), .A2(n41), .B1(i_data_bus[11]), .B2(n1), 
        .ZN(N103) );
  INVD1BWP30P140LVT U34 ( .I(i_data_bus[35]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U35 ( .A1(n19), .A2(n41), .B1(i_data_bus[3]), .B2(n2), 
        .ZN(N95) );
  INVD1BWP30P140LVT U36 ( .I(i_data_bus[36]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U37 ( .A1(n20), .A2(n41), .B1(i_data_bus[4]), .B2(n1), 
        .ZN(N96) );
  INVD1BWP30P140LVT U38 ( .I(i_data_bus[37]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U39 ( .A1(n21), .A2(n41), .B1(i_data_bus[5]), .B2(n2), 
        .ZN(N97) );
  INVD1BWP30P140LVT U40 ( .I(i_data_bus[38]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U41 ( .A1(n22), .A2(n41), .B1(i_data_bus[6]), .B2(n1), 
        .ZN(N98) );
  INVD1BWP30P140LVT U42 ( .I(i_data_bus[39]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U43 ( .A1(n23), .A2(n41), .B1(i_data_bus[7]), .B2(n2), 
        .ZN(N99) );
  INVD1BWP30P140LVT U44 ( .I(i_data_bus[40]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U45 ( .A1(n24), .A2(n41), .B1(i_data_bus[8]), .B2(n1), 
        .ZN(N100) );
  INVD1BWP30P140LVT U46 ( .I(i_data_bus[63]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U47 ( .A1(n25), .A2(n36), .B1(i_data_bus[31]), .B2(n1), 
        .ZN(N123) );
  INVD1BWP30P140LVT U48 ( .I(i_data_bus[44]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U49 ( .A1(n26), .A2(n36), .B1(i_data_bus[12]), .B2(n2), 
        .ZN(N104) );
  INVD1BWP30P140LVT U50 ( .I(i_data_bus[61]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U51 ( .A1(n27), .A2(n36), .B1(i_data_bus[29]), .B2(n1), 
        .ZN(N121) );
  INVD1BWP30P140LVT U52 ( .I(i_data_bus[59]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U53 ( .A1(n28), .A2(n36), .B1(i_data_bus[27]), .B2(n2), 
        .ZN(N119) );
  INVD1BWP30P140LVT U54 ( .I(i_data_bus[57]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U55 ( .A1(n29), .A2(n36), .B1(i_data_bus[25]), .B2(n1), 
        .ZN(N117) );
  INVD1BWP30P140LVT U56 ( .I(i_data_bus[55]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U57 ( .A1(n30), .A2(n36), .B1(i_data_bus[23]), .B2(n2), 
        .ZN(N115) );
  INVD1BWP30P140LVT U58 ( .I(i_data_bus[47]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U59 ( .A1(n31), .A2(n36), .B1(i_data_bus[15]), .B2(n1), 
        .ZN(N107) );
  INVD1BWP30P140LVT U60 ( .I(i_data_bus[45]), .ZN(n32) );
  MOAI22D1BWP30P140LVT U61 ( .A1(n32), .A2(n36), .B1(i_data_bus[13]), .B2(n2), 
        .ZN(N105) );
  INVD1BWP30P140LVT U62 ( .I(i_data_bus[51]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U63 ( .A1(n33), .A2(n36), .B1(i_data_bus[19]), .B2(n1), 
        .ZN(N111) );
  INVD1BWP30P140LVT U64 ( .I(i_data_bus[53]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U65 ( .A1(n34), .A2(n36), .B1(i_data_bus[21]), .B2(n2), 
        .ZN(N113) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[46]), .ZN(n35) );
  MOAI22D1BWP30P140LVT U67 ( .A1(n35), .A2(n36), .B1(i_data_bus[14]), .B2(n1), 
        .ZN(N106) );
  INVD1BWP30P140LVT U68 ( .I(i_data_bus[49]), .ZN(n37) );
  MOAI22D1BWP30P140LVT U69 ( .A1(n37), .A2(n36), .B1(i_data_bus[17]), .B2(n2), 
        .ZN(N109) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[56]), .ZN(n38) );
  MOAI22D1BWP30P140LVT U71 ( .A1(n38), .A2(n41), .B1(i_data_bus[24]), .B2(n1), 
        .ZN(N116) );
  INVD1BWP30P140LVT U72 ( .I(i_data_bus[60]), .ZN(n39) );
  MOAI22D1BWP30P140LVT U73 ( .A1(n39), .A2(n41), .B1(i_data_bus[28]), .B2(n2), 
        .ZN(N120) );
  INVD1BWP30P140LVT U74 ( .I(i_data_bus[58]), .ZN(n40) );
  MOAI22D1BWP30P140LVT U75 ( .A1(n40), .A2(n41), .B1(i_data_bus[26]), .B2(n1), 
        .ZN(N118) );
  INVD1BWP30P140LVT U76 ( .I(i_data_bus[62]), .ZN(n42) );
  MOAI22D1BWP30P140LVT U77 ( .A1(n42), .A2(n41), .B1(i_data_bus[30]), .B2(n2), 
        .ZN(N122) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_38 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_38 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_39 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U36 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_39 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_39 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_40 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_40 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_40 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_41 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_41 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_41 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_42 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_42 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_42 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_7 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_42 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_41 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_40 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_39 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_38 o_data_high ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_37 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_43 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n4), .A2(n3), .ZN(n2) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n4) );
  INVD1BWP30P140LVT U5 ( .I(n7), .ZN(n8) );
  NR2D1BWP30P140LVT U6 ( .A1(n4), .A2(n3), .ZN(n1) );
  INVD1BWP30P140LVT U7 ( .I(n8), .ZN(n36) );
  INVD1BWP30P140LVT U8 ( .I(n8), .ZN(n41) );
  OR2D1BWP30P140LVT U9 ( .A1(rst), .A2(i_cmd[0]), .Z(n3) );
  ND3D1BWP30P140LVT U10 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n6)
         );
  INVD1BWP30P140LVT U11 ( .I(rst), .ZN(n5) );
  IND2D1BWP30P140LVT U12 ( .A1(n6), .B1(n5), .ZN(n7) );
  IND2D1BWP30P140LVT U13 ( .A1(n2), .B1(n41), .ZN(N91) );
  INVD1BWP30P140LVT U14 ( .I(i_data_bus[52]), .ZN(n9) );
  MOAI22D1BWP30P140LVT U15 ( .A1(n9), .A2(n36), .B1(i_data_bus[20]), .B2(n2), 
        .ZN(N112) );
  INVD1BWP30P140LVT U16 ( .I(i_data_bus[48]), .ZN(n10) );
  MOAI22D1BWP30P140LVT U17 ( .A1(n10), .A2(n36), .B1(i_data_bus[16]), .B2(n1), 
        .ZN(N108) );
  INVD1BWP30P140LVT U18 ( .I(i_data_bus[54]), .ZN(n11) );
  MOAI22D1BWP30P140LVT U19 ( .A1(n11), .A2(n36), .B1(i_data_bus[22]), .B2(n2), 
        .ZN(N114) );
  INVD1BWP30P140LVT U20 ( .I(i_data_bus[50]), .ZN(n12) );
  MOAI22D1BWP30P140LVT U21 ( .A1(n12), .A2(n36), .B1(i_data_bus[18]), .B2(n1), 
        .ZN(N110) );
  INVD1BWP30P140LVT U22 ( .I(i_data_bus[43]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U23 ( .A1(n13), .A2(n41), .B1(i_data_bus[11]), .B2(n2), 
        .ZN(N103) );
  INVD1BWP30P140LVT U24 ( .I(i_data_bus[32]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U25 ( .A1(n14), .A2(n41), .B1(i_data_bus[0]), .B2(n1), 
        .ZN(N92) );
  INVD1BWP30P140LVT U26 ( .I(i_data_bus[38]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U27 ( .A1(n15), .A2(n41), .B1(i_data_bus[6]), .B2(n2), 
        .ZN(N98) );
  INVD1BWP30P140LVT U28 ( .I(i_data_bus[37]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U29 ( .A1(n16), .A2(n41), .B1(i_data_bus[5]), .B2(n1), 
        .ZN(N97) );
  INVD1BWP30P140LVT U30 ( .I(i_data_bus[36]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U31 ( .A1(n17), .A2(n41), .B1(i_data_bus[4]), .B2(n2), 
        .ZN(N96) );
  INVD1BWP30P140LVT U32 ( .I(i_data_bus[35]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U33 ( .A1(n18), .A2(n41), .B1(i_data_bus[3]), .B2(n1), 
        .ZN(N95) );
  INVD1BWP30P140LVT U34 ( .I(i_data_bus[34]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U35 ( .A1(n19), .A2(n41), .B1(i_data_bus[2]), .B2(n2), 
        .ZN(N94) );
  INVD1BWP30P140LVT U36 ( .I(i_data_bus[33]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U37 ( .A1(n20), .A2(n41), .B1(i_data_bus[1]), .B2(n1), 
        .ZN(N93) );
  INVD1BWP30P140LVT U38 ( .I(i_data_bus[42]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U39 ( .A1(n21), .A2(n41), .B1(i_data_bus[10]), .B2(n2), 
        .ZN(N102) );
  INVD1BWP30P140LVT U40 ( .I(i_data_bus[41]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U41 ( .A1(n22), .A2(n41), .B1(i_data_bus[9]), .B2(n1), 
        .ZN(N101) );
  INVD1BWP30P140LVT U42 ( .I(i_data_bus[40]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U43 ( .A1(n23), .A2(n41), .B1(i_data_bus[8]), .B2(n2), 
        .ZN(N100) );
  INVD1BWP30P140LVT U44 ( .I(i_data_bus[39]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U45 ( .A1(n24), .A2(n41), .B1(i_data_bus[7]), .B2(n1), 
        .ZN(N99) );
  INVD1BWP30P140LVT U46 ( .I(i_data_bus[45]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U47 ( .A1(n25), .A2(n36), .B1(i_data_bus[13]), .B2(n1), 
        .ZN(N105) );
  INVD1BWP30P140LVT U48 ( .I(i_data_bus[61]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U49 ( .A1(n26), .A2(n36), .B1(i_data_bus[29]), .B2(n2), 
        .ZN(N121) );
  INVD1BWP30P140LVT U50 ( .I(i_data_bus[63]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U51 ( .A1(n27), .A2(n36), .B1(i_data_bus[31]), .B2(n1), 
        .ZN(N123) );
  INVD1BWP30P140LVT U52 ( .I(i_data_bus[57]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U53 ( .A1(n28), .A2(n36), .B1(i_data_bus[25]), .B2(n2), 
        .ZN(N117) );
  INVD1BWP30P140LVT U54 ( .I(i_data_bus[46]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U55 ( .A1(n29), .A2(n36), .B1(i_data_bus[14]), .B2(n1), 
        .ZN(N106) );
  INVD1BWP30P140LVT U56 ( .I(i_data_bus[59]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U57 ( .A1(n30), .A2(n36), .B1(i_data_bus[27]), .B2(n2), 
        .ZN(N119) );
  INVD1BWP30P140LVT U58 ( .I(i_data_bus[44]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U59 ( .A1(n31), .A2(n36), .B1(i_data_bus[12]), .B2(n1), 
        .ZN(N104) );
  INVD1BWP30P140LVT U60 ( .I(i_data_bus[49]), .ZN(n32) );
  MOAI22D1BWP30P140LVT U61 ( .A1(n32), .A2(n36), .B1(i_data_bus[17]), .B2(n2), 
        .ZN(N109) );
  INVD1BWP30P140LVT U62 ( .I(i_data_bus[53]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U63 ( .A1(n33), .A2(n36), .B1(i_data_bus[21]), .B2(n1), 
        .ZN(N113) );
  INVD1BWP30P140LVT U64 ( .I(i_data_bus[55]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U65 ( .A1(n34), .A2(n36), .B1(i_data_bus[23]), .B2(n2), 
        .ZN(N115) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[51]), .ZN(n35) );
  MOAI22D1BWP30P140LVT U67 ( .A1(n35), .A2(n36), .B1(i_data_bus[19]), .B2(n1), 
        .ZN(N111) );
  INVD1BWP30P140LVT U68 ( .I(i_data_bus[47]), .ZN(n37) );
  MOAI22D1BWP30P140LVT U69 ( .A1(n37), .A2(n36), .B1(i_data_bus[15]), .B2(n2), 
        .ZN(N107) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[60]), .ZN(n38) );
  MOAI22D1BWP30P140LVT U71 ( .A1(n38), .A2(n41), .B1(i_data_bus[28]), .B2(n1), 
        .ZN(N120) );
  INVD1BWP30P140LVT U72 ( .I(i_data_bus[58]), .ZN(n39) );
  MOAI22D1BWP30P140LVT U73 ( .A1(n39), .A2(n41), .B1(i_data_bus[26]), .B2(n2), 
        .ZN(N118) );
  INVD1BWP30P140LVT U74 ( .I(i_data_bus[56]), .ZN(n40) );
  MOAI22D1BWP30P140LVT U75 ( .A1(n40), .A2(n41), .B1(i_data_bus[24]), .B2(n1), 
        .ZN(N116) );
  INVD1BWP30P140LVT U76 ( .I(i_data_bus[62]), .ZN(n42) );
  MOAI22D1BWP30P140LVT U77 ( .A1(n42), .A2(n41), .B1(i_data_bus[30]), .B2(n2), 
        .ZN(N122) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_43 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_43 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_44 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n4), .A2(n3), .ZN(n2) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n4) );
  INVD1BWP30P140LVT U5 ( .I(n7), .ZN(n8) );
  NR2D1BWP30P140LVT U6 ( .A1(n4), .A2(n3), .ZN(n1) );
  INVD1BWP30P140LVT U7 ( .I(n8), .ZN(n36) );
  INVD1BWP30P140LVT U8 ( .I(n8), .ZN(n41) );
  OR2D1BWP30P140LVT U9 ( .A1(rst), .A2(i_cmd[0]), .Z(n3) );
  ND3D1BWP30P140LVT U10 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n6)
         );
  INVD1BWP30P140LVT U11 ( .I(rst), .ZN(n5) );
  IND2D1BWP30P140LVT U12 ( .A1(n6), .B1(n5), .ZN(n7) );
  IND2D1BWP30P140LVT U13 ( .A1(n2), .B1(n41), .ZN(N91) );
  INVD1BWP30P140LVT U14 ( .I(i_data_bus[54]), .ZN(n9) );
  MOAI22D1BWP30P140LVT U15 ( .A1(n9), .A2(n36), .B1(i_data_bus[22]), .B2(n2), 
        .ZN(N114) );
  INVD1BWP30P140LVT U16 ( .I(i_data_bus[48]), .ZN(n10) );
  MOAI22D1BWP30P140LVT U17 ( .A1(n10), .A2(n36), .B1(i_data_bus[16]), .B2(n1), 
        .ZN(N108) );
  INVD1BWP30P140LVT U18 ( .I(i_data_bus[50]), .ZN(n11) );
  MOAI22D1BWP30P140LVT U19 ( .A1(n11), .A2(n36), .B1(i_data_bus[18]), .B2(n2), 
        .ZN(N110) );
  INVD1BWP30P140LVT U20 ( .I(i_data_bus[52]), .ZN(n12) );
  MOAI22D1BWP30P140LVT U21 ( .A1(n12), .A2(n36), .B1(i_data_bus[20]), .B2(n1), 
        .ZN(N112) );
  INVD1BWP30P140LVT U22 ( .I(i_data_bus[35]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U23 ( .A1(n13), .A2(n41), .B1(i_data_bus[3]), .B2(n2), 
        .ZN(N95) );
  INVD1BWP30P140LVT U24 ( .I(i_data_bus[34]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U25 ( .A1(n14), .A2(n41), .B1(i_data_bus[2]), .B2(n1), 
        .ZN(N94) );
  INVD1BWP30P140LVT U26 ( .I(i_data_bus[33]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U27 ( .A1(n15), .A2(n41), .B1(i_data_bus[1]), .B2(n2), 
        .ZN(N93) );
  INVD1BWP30P140LVT U28 ( .I(i_data_bus[43]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U29 ( .A1(n16), .A2(n41), .B1(i_data_bus[11]), .B2(n1), 
        .ZN(N103) );
  INVD1BWP30P140LVT U30 ( .I(i_data_bus[42]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U31 ( .A1(n17), .A2(n41), .B1(i_data_bus[10]), .B2(n2), 
        .ZN(N102) );
  INVD1BWP30P140LVT U32 ( .I(i_data_bus[32]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U33 ( .A1(n18), .A2(n41), .B1(i_data_bus[0]), .B2(n1), 
        .ZN(N92) );
  INVD1BWP30P140LVT U34 ( .I(i_data_bus[37]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U35 ( .A1(n19), .A2(n41), .B1(i_data_bus[5]), .B2(n2), 
        .ZN(N97) );
  INVD1BWP30P140LVT U36 ( .I(i_data_bus[41]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U37 ( .A1(n20), .A2(n41), .B1(i_data_bus[9]), .B2(n1), 
        .ZN(N101) );
  INVD1BWP30P140LVT U38 ( .I(i_data_bus[40]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U39 ( .A1(n21), .A2(n41), .B1(i_data_bus[8]), .B2(n2), 
        .ZN(N100) );
  INVD1BWP30P140LVT U40 ( .I(i_data_bus[39]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U41 ( .A1(n22), .A2(n41), .B1(i_data_bus[7]), .B2(n1), 
        .ZN(N99) );
  INVD1BWP30P140LVT U42 ( .I(i_data_bus[38]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U43 ( .A1(n23), .A2(n41), .B1(i_data_bus[6]), .B2(n2), 
        .ZN(N98) );
  INVD1BWP30P140LVT U44 ( .I(i_data_bus[36]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U45 ( .A1(n24), .A2(n41), .B1(i_data_bus[4]), .B2(n1), 
        .ZN(N96) );
  INVD1BWP30P140LVT U46 ( .I(i_data_bus[63]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U47 ( .A1(n25), .A2(n36), .B1(i_data_bus[31]), .B2(n1), 
        .ZN(N123) );
  INVD1BWP30P140LVT U48 ( .I(i_data_bus[44]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U49 ( .A1(n26), .A2(n36), .B1(i_data_bus[12]), .B2(n2), 
        .ZN(N104) );
  INVD1BWP30P140LVT U50 ( .I(i_data_bus[45]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U51 ( .A1(n27), .A2(n36), .B1(i_data_bus[13]), .B2(n1), 
        .ZN(N105) );
  INVD1BWP30P140LVT U52 ( .I(i_data_bus[46]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U53 ( .A1(n28), .A2(n36), .B1(i_data_bus[14]), .B2(n2), 
        .ZN(N106) );
  INVD1BWP30P140LVT U54 ( .I(i_data_bus[47]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U55 ( .A1(n29), .A2(n36), .B1(i_data_bus[15]), .B2(n1), 
        .ZN(N107) );
  INVD1BWP30P140LVT U56 ( .I(i_data_bus[49]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U57 ( .A1(n30), .A2(n36), .B1(i_data_bus[17]), .B2(n2), 
        .ZN(N109) );
  INVD1BWP30P140LVT U58 ( .I(i_data_bus[59]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U59 ( .A1(n31), .A2(n36), .B1(i_data_bus[27]), .B2(n1), 
        .ZN(N119) );
  INVD1BWP30P140LVT U60 ( .I(i_data_bus[51]), .ZN(n32) );
  MOAI22D1BWP30P140LVT U61 ( .A1(n32), .A2(n36), .B1(i_data_bus[19]), .B2(n2), 
        .ZN(N111) );
  INVD1BWP30P140LVT U62 ( .I(i_data_bus[53]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U63 ( .A1(n33), .A2(n36), .B1(i_data_bus[21]), .B2(n1), 
        .ZN(N113) );
  INVD1BWP30P140LVT U64 ( .I(i_data_bus[55]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U65 ( .A1(n34), .A2(n36), .B1(i_data_bus[23]), .B2(n2), 
        .ZN(N115) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[57]), .ZN(n35) );
  MOAI22D1BWP30P140LVT U67 ( .A1(n35), .A2(n36), .B1(i_data_bus[25]), .B2(n1), 
        .ZN(N117) );
  INVD1BWP30P140LVT U68 ( .I(i_data_bus[61]), .ZN(n37) );
  MOAI22D1BWP30P140LVT U69 ( .A1(n37), .A2(n36), .B1(i_data_bus[29]), .B2(n2), 
        .ZN(N121) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[58]), .ZN(n38) );
  MOAI22D1BWP30P140LVT U71 ( .A1(n38), .A2(n41), .B1(i_data_bus[26]), .B2(n1), 
        .ZN(N118) );
  INVD1BWP30P140LVT U72 ( .I(i_data_bus[62]), .ZN(n39) );
  MOAI22D1BWP30P140LVT U73 ( .A1(n39), .A2(n41), .B1(i_data_bus[30]), .B2(n2), 
        .ZN(N122) );
  INVD1BWP30P140LVT U74 ( .I(i_data_bus[56]), .ZN(n40) );
  MOAI22D1BWP30P140LVT U75 ( .A1(n40), .A2(n41), .B1(i_data_bus[24]), .B2(n1), 
        .ZN(N116) );
  INVD1BWP30P140LVT U76 ( .I(i_data_bus[60]), .ZN(n42) );
  MOAI22D1BWP30P140LVT U77 ( .A1(n42), .A2(n41), .B1(i_data_bus[28]), .B2(n2), 
        .ZN(N120) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_44 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_44 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_45 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U36 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_45 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_45 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_46 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  IND2D1BWP30P140LVT U3 ( .A1(n1), .B1(i_valid[0]), .ZN(n2) );
  INVD1BWP30P140LVT U4 ( .I(i_en), .ZN(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  NR3D1P5BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n6) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  BUFFD2BWP30P140LVT U8 ( .I(n4), .Z(n5) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n5), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n5), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n5), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n5), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n5), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n5), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n5), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n5), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n5), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n5), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n5), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n5), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n5), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n5), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n5), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n5), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n5), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n5), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n5), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n5), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n5), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n5), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n5), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n5), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n5), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n5), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n5), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n5), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n5), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n5), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n5), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n5), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n5), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_46 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_46 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_47 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3OPTPAD2BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  NR2D1BWP30P140LVT U4 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U5 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U8 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_47 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_47 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_48 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3OPTPAD2BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  NR2D1BWP30P140LVT U4 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U5 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U8 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_48 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_48 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_8 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_48 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_47 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_46 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_45 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_44 o_data_high ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_43 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_49 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  CKBD1BWP30P140LVT U3 ( .I(n2), .Z(n70) );
  NR2D1BWP30P140LVT U4 ( .A1(n1), .A2(rst), .ZN(n2) );
  INVD1BWP30P140LVT U5 ( .I(n4), .ZN(n69) );
  OR3D1BWP30P140LVT U6 ( .A1(n3), .A2(rst), .A3(i_cmd[0]), .Z(n4) );
  ND2D1BWP30P140LVT U7 ( .A1(i_en), .A2(i_valid[0]), .ZN(n3) );
  ND2D1BWP30P140LVT U8 ( .A1(n68), .A2(n67), .ZN(N92) );
  ND2OPTIBD1BWP30P140LVT U9 ( .A1(n69), .A2(i_data_bus[0]), .ZN(n67) );
  ND2OPTIBD1BWP30P140LVT U10 ( .A1(n70), .A2(i_data_bus[32]), .ZN(n68) );
  ND2D1BWP30P140LVT U11 ( .A1(n6), .A2(n5), .ZN(N93) );
  ND2OPTIBD1BWP30P140LVT U12 ( .A1(n69), .A2(i_data_bus[1]), .ZN(n5) );
  ND2OPTIBD1BWP30P140LVT U13 ( .A1(n70), .A2(i_data_bus[33]), .ZN(n6) );
  ND2D1BWP30P140LVT U14 ( .A1(n8), .A2(n7), .ZN(N94) );
  ND2OPTIBD1BWP30P140LVT U15 ( .A1(n69), .A2(i_data_bus[2]), .ZN(n7) );
  ND2OPTIBD1BWP30P140LVT U16 ( .A1(n70), .A2(i_data_bus[34]), .ZN(n8) );
  ND2D1BWP30P140LVT U17 ( .A1(n10), .A2(n9), .ZN(N95) );
  ND2OPTIBD1BWP30P140LVT U18 ( .A1(n69), .A2(i_data_bus[3]), .ZN(n9) );
  ND2OPTIBD1BWP30P140LVT U19 ( .A1(n70), .A2(i_data_bus[35]), .ZN(n10) );
  ND2D1BWP30P140LVT U20 ( .A1(n12), .A2(n11), .ZN(N96) );
  ND2OPTIBD1BWP30P140LVT U21 ( .A1(n69), .A2(i_data_bus[4]), .ZN(n11) );
  ND2OPTIBD1BWP30P140LVT U22 ( .A1(n70), .A2(i_data_bus[36]), .ZN(n12) );
  ND2D1BWP30P140LVT U23 ( .A1(n14), .A2(n13), .ZN(N97) );
  ND2OPTIBD1BWP30P140LVT U24 ( .A1(n69), .A2(i_data_bus[5]), .ZN(n13) );
  ND2OPTIBD1BWP30P140LVT U25 ( .A1(n70), .A2(i_data_bus[37]), .ZN(n14) );
  ND2D1BWP30P140LVT U26 ( .A1(n16), .A2(n15), .ZN(N98) );
  ND2OPTIBD1BWP30P140LVT U27 ( .A1(n69), .A2(i_data_bus[6]), .ZN(n15) );
  ND2OPTIBD1BWP30P140LVT U28 ( .A1(n70), .A2(i_data_bus[38]), .ZN(n16) );
  ND2D1BWP30P140LVT U29 ( .A1(n18), .A2(n17), .ZN(N99) );
  ND2OPTIBD1BWP30P140LVT U30 ( .A1(n69), .A2(i_data_bus[7]), .ZN(n17) );
  ND2OPTIBD1BWP30P140LVT U31 ( .A1(n70), .A2(i_data_bus[39]), .ZN(n18) );
  ND2D1BWP30P140LVT U32 ( .A1(n20), .A2(n19), .ZN(N100) );
  ND2OPTIBD1BWP30P140LVT U33 ( .A1(n69), .A2(i_data_bus[8]), .ZN(n19) );
  ND2OPTIBD1BWP30P140LVT U34 ( .A1(n70), .A2(i_data_bus[40]), .ZN(n20) );
  ND2D1BWP30P140LVT U35 ( .A1(n22), .A2(n21), .ZN(N101) );
  ND2OPTIBD1BWP30P140LVT U36 ( .A1(n69), .A2(i_data_bus[9]), .ZN(n21) );
  ND2OPTIBD1BWP30P140LVT U37 ( .A1(n70), .A2(i_data_bus[41]), .ZN(n22) );
  ND2D1BWP30P140LVT U38 ( .A1(n24), .A2(n23), .ZN(N102) );
  ND2OPTIBD1BWP30P140LVT U39 ( .A1(n69), .A2(i_data_bus[10]), .ZN(n23) );
  ND2OPTIBD1BWP30P140LVT U40 ( .A1(n70), .A2(i_data_bus[42]), .ZN(n24) );
  ND2D1BWP30P140LVT U41 ( .A1(n26), .A2(n25), .ZN(N103) );
  ND2OPTIBD1BWP30P140LVT U42 ( .A1(n69), .A2(i_data_bus[11]), .ZN(n25) );
  ND2OPTIBD1BWP30P140LVT U43 ( .A1(n70), .A2(i_data_bus[43]), .ZN(n26) );
  ND2D1BWP30P140LVT U44 ( .A1(n28), .A2(n27), .ZN(N104) );
  ND2OPTIBD1BWP30P140LVT U45 ( .A1(n69), .A2(i_data_bus[12]), .ZN(n27) );
  ND2OPTIBD1BWP30P140LVT U46 ( .A1(n70), .A2(i_data_bus[44]), .ZN(n28) );
  ND2D1BWP30P140LVT U47 ( .A1(n30), .A2(n29), .ZN(N105) );
  ND2OPTIBD1BWP30P140LVT U48 ( .A1(n69), .A2(i_data_bus[13]), .ZN(n29) );
  ND2OPTIBD1BWP30P140LVT U49 ( .A1(n70), .A2(i_data_bus[45]), .ZN(n30) );
  ND2D1BWP30P140LVT U50 ( .A1(n32), .A2(n31), .ZN(N106) );
  ND2OPTIBD1BWP30P140LVT U51 ( .A1(n69), .A2(i_data_bus[14]), .ZN(n31) );
  ND2OPTIBD1BWP30P140LVT U52 ( .A1(n70), .A2(i_data_bus[46]), .ZN(n32) );
  ND2D1BWP30P140LVT U53 ( .A1(n34), .A2(n33), .ZN(N107) );
  ND2OPTIBD1BWP30P140LVT U54 ( .A1(n69), .A2(i_data_bus[15]), .ZN(n33) );
  ND2OPTIBD1BWP30P140LVT U55 ( .A1(n70), .A2(i_data_bus[47]), .ZN(n34) );
  ND2D1BWP30P140LVT U56 ( .A1(n36), .A2(n35), .ZN(N108) );
  ND2OPTIBD1BWP30P140LVT U57 ( .A1(n69), .A2(i_data_bus[16]), .ZN(n35) );
  ND2OPTIBD1BWP30P140LVT U58 ( .A1(n70), .A2(i_data_bus[48]), .ZN(n36) );
  ND2D1BWP30P140LVT U59 ( .A1(n38), .A2(n37), .ZN(N109) );
  ND2OPTIBD1BWP30P140LVT U60 ( .A1(n69), .A2(i_data_bus[17]), .ZN(n37) );
  ND2OPTIBD1BWP30P140LVT U61 ( .A1(n70), .A2(i_data_bus[49]), .ZN(n38) );
  ND2D1BWP30P140LVT U62 ( .A1(n40), .A2(n39), .ZN(N110) );
  ND2OPTIBD1BWP30P140LVT U63 ( .A1(n69), .A2(i_data_bus[18]), .ZN(n39) );
  ND2OPTIBD1BWP30P140LVT U64 ( .A1(n70), .A2(i_data_bus[50]), .ZN(n40) );
  ND2D1BWP30P140LVT U65 ( .A1(n42), .A2(n41), .ZN(N111) );
  ND2OPTIBD1BWP30P140LVT U66 ( .A1(n69), .A2(i_data_bus[19]), .ZN(n41) );
  ND2OPTIBD1BWP30P140LVT U67 ( .A1(n70), .A2(i_data_bus[51]), .ZN(n42) );
  ND2D1BWP30P140LVT U68 ( .A1(n44), .A2(n43), .ZN(N112) );
  ND2OPTIBD1BWP30P140LVT U69 ( .A1(n69), .A2(i_data_bus[20]), .ZN(n43) );
  ND2OPTIBD1BWP30P140LVT U70 ( .A1(n70), .A2(i_data_bus[52]), .ZN(n44) );
  ND2D1BWP30P140LVT U71 ( .A1(n46), .A2(n45), .ZN(N113) );
  ND2OPTIBD1BWP30P140LVT U72 ( .A1(n69), .A2(i_data_bus[21]), .ZN(n45) );
  ND2OPTIBD1BWP30P140LVT U73 ( .A1(n70), .A2(i_data_bus[53]), .ZN(n46) );
  ND2D1BWP30P140LVT U74 ( .A1(n48), .A2(n47), .ZN(N114) );
  ND2OPTIBD1BWP30P140LVT U75 ( .A1(n69), .A2(i_data_bus[22]), .ZN(n47) );
  ND2OPTIBD1BWP30P140LVT U76 ( .A1(n70), .A2(i_data_bus[54]), .ZN(n48) );
  ND2D1BWP30P140LVT U77 ( .A1(n50), .A2(n49), .ZN(N115) );
  ND2OPTIBD1BWP30P140LVT U78 ( .A1(n69), .A2(i_data_bus[23]), .ZN(n49) );
  ND2OPTIBD1BWP30P140LVT U79 ( .A1(n70), .A2(i_data_bus[55]), .ZN(n50) );
  ND2D1BWP30P140LVT U80 ( .A1(n52), .A2(n51), .ZN(N116) );
  ND2OPTIBD1BWP30P140LVT U81 ( .A1(n69), .A2(i_data_bus[24]), .ZN(n51) );
  ND2OPTIBD1BWP30P140LVT U82 ( .A1(n70), .A2(i_data_bus[56]), .ZN(n52) );
  ND2D1BWP30P140LVT U83 ( .A1(n54), .A2(n53), .ZN(N117) );
  ND2OPTIBD1BWP30P140LVT U84 ( .A1(n69), .A2(i_data_bus[25]), .ZN(n53) );
  ND2OPTIBD1BWP30P140LVT U85 ( .A1(n70), .A2(i_data_bus[57]), .ZN(n54) );
  ND2D1BWP30P140LVT U86 ( .A1(n56), .A2(n55), .ZN(N118) );
  ND2OPTIBD1BWP30P140LVT U87 ( .A1(n69), .A2(i_data_bus[26]), .ZN(n55) );
  ND2OPTIBD1BWP30P140LVT U88 ( .A1(n70), .A2(i_data_bus[58]), .ZN(n56) );
  ND2D1BWP30P140LVT U89 ( .A1(n58), .A2(n57), .ZN(N119) );
  ND2OPTIBD1BWP30P140LVT U90 ( .A1(n69), .A2(i_data_bus[27]), .ZN(n57) );
  ND2OPTIBD1BWP30P140LVT U91 ( .A1(n70), .A2(i_data_bus[59]), .ZN(n58) );
  ND2D1BWP30P140LVT U92 ( .A1(n60), .A2(n59), .ZN(N120) );
  ND2OPTIBD1BWP30P140LVT U93 ( .A1(n69), .A2(i_data_bus[28]), .ZN(n59) );
  ND2OPTIBD1BWP30P140LVT U94 ( .A1(n70), .A2(i_data_bus[60]), .ZN(n60) );
  ND2D1BWP30P140LVT U95 ( .A1(n62), .A2(n61), .ZN(N121) );
  ND2OPTIBD1BWP30P140LVT U96 ( .A1(n69), .A2(i_data_bus[29]), .ZN(n61) );
  ND2OPTIBD1BWP30P140LVT U97 ( .A1(n70), .A2(i_data_bus[61]), .ZN(n62) );
  ND2D1BWP30P140LVT U98 ( .A1(n64), .A2(n63), .ZN(N122) );
  ND2OPTIBD1BWP30P140LVT U99 ( .A1(n69), .A2(i_data_bus[30]), .ZN(n63) );
  ND2OPTIBD1BWP30P140LVT U100 ( .A1(n70), .A2(i_data_bus[62]), .ZN(n64) );
  ND2D1BWP30P140LVT U101 ( .A1(n66), .A2(n65), .ZN(N123) );
  ND2OPTIBD1BWP30P140LVT U102 ( .A1(n69), .A2(i_data_bus[31]), .ZN(n65) );
  ND2OPTIBD1BWP30P140LVT U103 ( .A1(n70), .A2(i_data_bus[63]), .ZN(n66) );
  IND2D1BWP30P140LVT U104 ( .A1(n70), .B1(n4), .ZN(N91) );
  ND3D1BWP30P140LVT U105 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n1)
         );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_49 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_49 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_50 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n34), .Z(n70) );
  INVD1BWP30P140LVT U4 ( .I(n36), .ZN(n69) );
  OR3D1BWP30P140LVT U5 ( .A1(n35), .A2(rst), .A3(i_cmd[0]), .Z(n36) );
  ND2D1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n35) );
  IND2D1BWP30P140LVT U7 ( .A1(n1), .B1(n37), .ZN(N92) );
  ND2OPTIBD1BWP30P140LVT U8 ( .A1(n69), .A2(i_data_bus[0]), .ZN(n37) );
  IND2D1BWP30P140LVT U9 ( .A1(n2), .B1(n38), .ZN(N93) );
  ND2OPTIBD1BWP30P140LVT U10 ( .A1(n69), .A2(i_data_bus[1]), .ZN(n38) );
  IND2D1BWP30P140LVT U11 ( .A1(n3), .B1(n39), .ZN(N94) );
  ND2OPTIBD1BWP30P140LVT U12 ( .A1(n69), .A2(i_data_bus[2]), .ZN(n39) );
  IND2D1BWP30P140LVT U13 ( .A1(n4), .B1(n40), .ZN(N95) );
  ND2OPTIBD1BWP30P140LVT U14 ( .A1(n69), .A2(i_data_bus[3]), .ZN(n40) );
  IND2D1BWP30P140LVT U15 ( .A1(n5), .B1(n41), .ZN(N96) );
  ND2OPTIBD1BWP30P140LVT U16 ( .A1(n69), .A2(i_data_bus[4]), .ZN(n41) );
  IND2D1BWP30P140LVT U17 ( .A1(n6), .B1(n42), .ZN(N97) );
  ND2OPTIBD1BWP30P140LVT U18 ( .A1(n69), .A2(i_data_bus[5]), .ZN(n42) );
  IND2D1BWP30P140LVT U19 ( .A1(n7), .B1(n43), .ZN(N98) );
  ND2OPTIBD1BWP30P140LVT U20 ( .A1(n69), .A2(i_data_bus[6]), .ZN(n43) );
  IND2D1BWP30P140LVT U21 ( .A1(n8), .B1(n44), .ZN(N99) );
  ND2OPTIBD1BWP30P140LVT U22 ( .A1(n69), .A2(i_data_bus[7]), .ZN(n44) );
  IND2D1BWP30P140LVT U23 ( .A1(n9), .B1(n45), .ZN(N100) );
  ND2OPTIBD1BWP30P140LVT U24 ( .A1(n69), .A2(i_data_bus[8]), .ZN(n45) );
  IND2D1BWP30P140LVT U25 ( .A1(n10), .B1(n46), .ZN(N101) );
  ND2OPTIBD1BWP30P140LVT U26 ( .A1(n69), .A2(i_data_bus[9]), .ZN(n46) );
  IND2D1BWP30P140LVT U27 ( .A1(n11), .B1(n47), .ZN(N102) );
  ND2OPTIBD1BWP30P140LVT U28 ( .A1(n69), .A2(i_data_bus[10]), .ZN(n47) );
  IND2D1BWP30P140LVT U29 ( .A1(n12), .B1(n48), .ZN(N103) );
  ND2OPTIBD1BWP30P140LVT U30 ( .A1(n69), .A2(i_data_bus[11]), .ZN(n48) );
  IND2D1BWP30P140LVT U31 ( .A1(n13), .B1(n49), .ZN(N104) );
  ND2OPTIBD1BWP30P140LVT U32 ( .A1(n69), .A2(i_data_bus[12]), .ZN(n49) );
  IND2D1BWP30P140LVT U33 ( .A1(n14), .B1(n50), .ZN(N105) );
  ND2OPTIBD1BWP30P140LVT U34 ( .A1(n69), .A2(i_data_bus[13]), .ZN(n50) );
  IND2D1BWP30P140LVT U35 ( .A1(n15), .B1(n51), .ZN(N106) );
  ND2OPTIBD1BWP30P140LVT U36 ( .A1(n69), .A2(i_data_bus[14]), .ZN(n51) );
  IND2D1BWP30P140LVT U37 ( .A1(n16), .B1(n52), .ZN(N107) );
  ND2OPTIBD1BWP30P140LVT U38 ( .A1(n69), .A2(i_data_bus[15]), .ZN(n52) );
  IND2D1BWP30P140LVT U39 ( .A1(n17), .B1(n53), .ZN(N108) );
  ND2OPTIBD1BWP30P140LVT U40 ( .A1(n69), .A2(i_data_bus[16]), .ZN(n53) );
  IND2D1BWP30P140LVT U41 ( .A1(n18), .B1(n54), .ZN(N109) );
  ND2OPTIBD1BWP30P140LVT U42 ( .A1(n69), .A2(i_data_bus[17]), .ZN(n54) );
  IND2D1BWP30P140LVT U43 ( .A1(n19), .B1(n55), .ZN(N110) );
  ND2OPTIBD1BWP30P140LVT U44 ( .A1(n69), .A2(i_data_bus[18]), .ZN(n55) );
  IND2D1BWP30P140LVT U45 ( .A1(n20), .B1(n56), .ZN(N111) );
  ND2OPTIBD1BWP30P140LVT U46 ( .A1(n69), .A2(i_data_bus[19]), .ZN(n56) );
  IND2D1BWP30P140LVT U47 ( .A1(n21), .B1(n57), .ZN(N112) );
  ND2OPTIBD1BWP30P140LVT U48 ( .A1(n69), .A2(i_data_bus[20]), .ZN(n57) );
  IND2D1BWP30P140LVT U49 ( .A1(n22), .B1(n58), .ZN(N113) );
  ND2OPTIBD1BWP30P140LVT U50 ( .A1(n69), .A2(i_data_bus[21]), .ZN(n58) );
  IND2D1BWP30P140LVT U51 ( .A1(n23), .B1(n59), .ZN(N114) );
  ND2OPTIBD1BWP30P140LVT U52 ( .A1(n69), .A2(i_data_bus[22]), .ZN(n59) );
  IND2D1BWP30P140LVT U53 ( .A1(n24), .B1(n60), .ZN(N115) );
  ND2OPTIBD1BWP30P140LVT U54 ( .A1(n69), .A2(i_data_bus[23]), .ZN(n60) );
  IND2D1BWP30P140LVT U55 ( .A1(n25), .B1(n61), .ZN(N116) );
  ND2OPTIBD1BWP30P140LVT U56 ( .A1(n69), .A2(i_data_bus[24]), .ZN(n61) );
  IND2D1BWP30P140LVT U57 ( .A1(n26), .B1(n62), .ZN(N117) );
  ND2OPTIBD1BWP30P140LVT U58 ( .A1(n69), .A2(i_data_bus[25]), .ZN(n62) );
  IND2D1BWP30P140LVT U59 ( .A1(n27), .B1(n63), .ZN(N118) );
  ND2OPTIBD1BWP30P140LVT U60 ( .A1(n69), .A2(i_data_bus[26]), .ZN(n63) );
  IND2D1BWP30P140LVT U61 ( .A1(n28), .B1(n64), .ZN(N119) );
  ND2OPTIBD1BWP30P140LVT U62 ( .A1(n69), .A2(i_data_bus[27]), .ZN(n64) );
  IND2D1BWP30P140LVT U63 ( .A1(n29), .B1(n65), .ZN(N120) );
  ND2OPTIBD1BWP30P140LVT U64 ( .A1(n69), .A2(i_data_bus[28]), .ZN(n65) );
  IND2D1BWP30P140LVT U65 ( .A1(n30), .B1(n66), .ZN(N121) );
  ND2OPTIBD1BWP30P140LVT U66 ( .A1(n69), .A2(i_data_bus[29]), .ZN(n66) );
  IND2D1BWP30P140LVT U67 ( .A1(n31), .B1(n67), .ZN(N122) );
  ND2OPTIBD1BWP30P140LVT U68 ( .A1(n69), .A2(i_data_bus[30]), .ZN(n67) );
  IND2D1BWP30P140LVT U69 ( .A1(n32), .B1(n68), .ZN(N123) );
  ND2OPTIBD1BWP30P140LVT U70 ( .A1(n69), .A2(i_data_bus[31]), .ZN(n68) );
  IND2D1BWP30P140LVT U71 ( .A1(n70), .B1(n36), .ZN(N91) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n70), .A2(i_data_bus[32]), .Z(n1) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n70), .A2(i_data_bus[33]), .Z(n2) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n70), .A2(i_data_bus[34]), .Z(n3) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n70), .A2(i_data_bus[35]), .Z(n4) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n70), .A2(i_data_bus[36]), .Z(n5) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n70), .A2(i_data_bus[37]), .Z(n6) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n70), .A2(i_data_bus[38]), .Z(n7) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n70), .A2(i_data_bus[39]), .Z(n8) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n70), .A2(i_data_bus[40]), .Z(n9) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n70), .A2(i_data_bus[41]), .Z(n10) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n70), .A2(i_data_bus[42]), .Z(n11) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n70), .A2(i_data_bus[43]), .Z(n12) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n70), .A2(i_data_bus[44]), .Z(n13) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n70), .A2(i_data_bus[45]), .Z(n14) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n70), .A2(i_data_bus[46]), .Z(n15) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n70), .A2(i_data_bus[47]), .Z(n16) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n70), .A2(i_data_bus[48]), .Z(n17) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n70), .A2(i_data_bus[49]), .Z(n18) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n70), .A2(i_data_bus[50]), .Z(n19) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n70), .A2(i_data_bus[51]), .Z(n20) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n70), .A2(i_data_bus[52]), .Z(n21) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n70), .A2(i_data_bus[53]), .Z(n22) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n70), .A2(i_data_bus[54]), .Z(n23) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n70), .A2(i_data_bus[55]), .Z(n24) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n70), .A2(i_data_bus[56]), .Z(n25) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n70), .A2(i_data_bus[57]), .Z(n26) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n70), .A2(i_data_bus[58]), .Z(n27) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n70), .A2(i_data_bus[59]), .Z(n28) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n70), .A2(i_data_bus[60]), .Z(n29) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n70), .A2(i_data_bus[61]), .Z(n30) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n70), .A2(i_data_bus[62]), .Z(n31) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n70), .A2(i_data_bus[63]), .Z(n32) );
  ND3D1BWP30P140LVT U104 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n33)
         );
  NR2D1BWP30P140LVT U105 ( .A1(n33), .A2(rst), .ZN(n34) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_50 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_50 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_51 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2D1BWP30P140LVT U3 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3D1P5BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U36 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_51 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_51 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_52 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2OPTPAD1BWP30P140LVT U3 ( .A1(i_cmd[0]), .A2(n2), .ZN(n6) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_valid[0]), .A2(n1), .ZN(n2) );
  INR2D1BWP30P140LVT U5 ( .A1(i_en), .B1(rst), .ZN(n1) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  NR2D1BWP30P140LVT U7 ( .A1(n3), .A2(rst), .ZN(n4) );
  BUFFD2BWP30P140LVT U8 ( .I(n4), .Z(n5) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n5), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n5), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n5), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n5), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n5), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n5), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n5), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n5), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n5), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n5), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n5), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n5), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n5), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n5), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n5), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n5), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n5), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n5), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n5), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n5), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n5), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n5), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n5), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n5), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n5), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n5), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n5), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n5), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n5), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n5), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n5), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n5), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n5), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_52 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_52 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_53 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  BUFFD2BWP30P140LVT U3 ( .I(n13), .Z(n70) );
  NR3D1P5BWP30P140LVT U4 ( .A1(n14), .A2(rst), .A3(i_cmd[0]), .ZN(n1) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n14) );
  IND2D1BWP30P140LVT U6 ( .A1(n70), .B1(n69), .ZN(N91) );
  INVD1BWP30P140LVT U7 ( .I(n1), .ZN(n69) );
  ND2OPTIBD1BWP30P140LVT U8 ( .A1(n26), .A2(n25), .ZN(N92) );
  ND2OPTIBD1BWP30P140LVT U9 ( .A1(n1), .A2(i_data_bus[0]), .ZN(n25) );
  ND2D1BWP30P140LVT U10 ( .A1(n70), .A2(i_data_bus[32]), .ZN(n26) );
  ND2OPTIBD1BWP30P140LVT U11 ( .A1(n28), .A2(n27), .ZN(N93) );
  ND2OPTIBD1BWP30P140LVT U12 ( .A1(n1), .A2(i_data_bus[1]), .ZN(n27) );
  ND2D1BWP30P140LVT U13 ( .A1(n70), .A2(i_data_bus[33]), .ZN(n28) );
  ND2OPTIBD1BWP30P140LVT U14 ( .A1(n30), .A2(n29), .ZN(N94) );
  ND2OPTIBD1BWP30P140LVT U15 ( .A1(n1), .A2(i_data_bus[2]), .ZN(n29) );
  ND2D1BWP30P140LVT U16 ( .A1(n70), .A2(i_data_bus[34]), .ZN(n30) );
  ND2OPTIBD1BWP30P140LVT U17 ( .A1(n32), .A2(n31), .ZN(N95) );
  ND2OPTIBD1BWP30P140LVT U18 ( .A1(n1), .A2(i_data_bus[3]), .ZN(n31) );
  ND2D1BWP30P140LVT U19 ( .A1(n70), .A2(i_data_bus[35]), .ZN(n32) );
  ND2OPTIBD1BWP30P140LVT U20 ( .A1(n34), .A2(n33), .ZN(N96) );
  ND2OPTIBD1BWP30P140LVT U21 ( .A1(n1), .A2(i_data_bus[4]), .ZN(n33) );
  ND2D1BWP30P140LVT U22 ( .A1(n70), .A2(i_data_bus[36]), .ZN(n34) );
  ND2OPTIBD1BWP30P140LVT U23 ( .A1(n36), .A2(n35), .ZN(N97) );
  ND2OPTIBD1BWP30P140LVT U24 ( .A1(n1), .A2(i_data_bus[5]), .ZN(n35) );
  ND2D1BWP30P140LVT U25 ( .A1(n70), .A2(i_data_bus[37]), .ZN(n36) );
  ND2OPTIBD1BWP30P140LVT U26 ( .A1(n38), .A2(n37), .ZN(N98) );
  ND2OPTIBD1BWP30P140LVT U27 ( .A1(n1), .A2(i_data_bus[6]), .ZN(n37) );
  ND2D1BWP30P140LVT U28 ( .A1(n70), .A2(i_data_bus[38]), .ZN(n38) );
  ND2OPTIBD1BWP30P140LVT U29 ( .A1(n40), .A2(n39), .ZN(N99) );
  ND2OPTIBD1BWP30P140LVT U30 ( .A1(n1), .A2(i_data_bus[7]), .ZN(n39) );
  ND2D1BWP30P140LVT U31 ( .A1(n70), .A2(i_data_bus[39]), .ZN(n40) );
  ND2OPTIBD1BWP30P140LVT U32 ( .A1(n42), .A2(n41), .ZN(N100) );
  ND2OPTIBD1BWP30P140LVT U33 ( .A1(n1), .A2(i_data_bus[8]), .ZN(n41) );
  ND2D1BWP30P140LVT U34 ( .A1(n70), .A2(i_data_bus[40]), .ZN(n42) );
  ND2OPTIBD1BWP30P140LVT U35 ( .A1(n44), .A2(n43), .ZN(N101) );
  ND2OPTIBD1BWP30P140LVT U36 ( .A1(n1), .A2(i_data_bus[9]), .ZN(n43) );
  ND2D1BWP30P140LVT U37 ( .A1(n70), .A2(i_data_bus[41]), .ZN(n44) );
  ND2OPTIBD1BWP30P140LVT U38 ( .A1(n46), .A2(n45), .ZN(N102) );
  ND2OPTIBD1BWP30P140LVT U39 ( .A1(n1), .A2(i_data_bus[10]), .ZN(n45) );
  ND2D1BWP30P140LVT U40 ( .A1(n70), .A2(i_data_bus[42]), .ZN(n46) );
  ND2OPTIBD1BWP30P140LVT U41 ( .A1(n48), .A2(n47), .ZN(N103) );
  ND2OPTIBD1BWP30P140LVT U42 ( .A1(n1), .A2(i_data_bus[11]), .ZN(n47) );
  ND2D1BWP30P140LVT U43 ( .A1(n70), .A2(i_data_bus[43]), .ZN(n48) );
  ND2OPTIBD1BWP30P140LVT U44 ( .A1(n50), .A2(n49), .ZN(N104) );
  ND2OPTIBD1BWP30P140LVT U45 ( .A1(n1), .A2(i_data_bus[12]), .ZN(n49) );
  ND2D1BWP30P140LVT U46 ( .A1(n70), .A2(i_data_bus[44]), .ZN(n50) );
  ND2OPTIBD1BWP30P140LVT U47 ( .A1(n52), .A2(n51), .ZN(N105) );
  ND2OPTIBD1BWP30P140LVT U48 ( .A1(n1), .A2(i_data_bus[13]), .ZN(n51) );
  ND2D1BWP30P140LVT U49 ( .A1(n70), .A2(i_data_bus[45]), .ZN(n52) );
  ND2OPTIBD1BWP30P140LVT U50 ( .A1(n54), .A2(n53), .ZN(N106) );
  ND2OPTIBD1BWP30P140LVT U51 ( .A1(n1), .A2(i_data_bus[14]), .ZN(n53) );
  ND2D1BWP30P140LVT U52 ( .A1(n70), .A2(i_data_bus[46]), .ZN(n54) );
  ND2OPTIBD1BWP30P140LVT U53 ( .A1(n56), .A2(n55), .ZN(N107) );
  ND2OPTIBD1BWP30P140LVT U54 ( .A1(n1), .A2(i_data_bus[15]), .ZN(n55) );
  ND2D1BWP30P140LVT U55 ( .A1(n70), .A2(i_data_bus[47]), .ZN(n56) );
  ND2OPTIBD1BWP30P140LVT U56 ( .A1(n58), .A2(n57), .ZN(N108) );
  ND2OPTIBD1BWP30P140LVT U57 ( .A1(n1), .A2(i_data_bus[16]), .ZN(n57) );
  ND2D1BWP30P140LVT U58 ( .A1(n70), .A2(i_data_bus[48]), .ZN(n58) );
  ND2OPTIBD1BWP30P140LVT U59 ( .A1(n60), .A2(n59), .ZN(N109) );
  ND2OPTIBD1BWP30P140LVT U60 ( .A1(n1), .A2(i_data_bus[17]), .ZN(n59) );
  ND2D1BWP30P140LVT U61 ( .A1(n70), .A2(i_data_bus[49]), .ZN(n60) );
  ND2OPTIBD1BWP30P140LVT U62 ( .A1(n62), .A2(n61), .ZN(N110) );
  ND2OPTIBD1BWP30P140LVT U63 ( .A1(n1), .A2(i_data_bus[18]), .ZN(n61) );
  ND2D1BWP30P140LVT U64 ( .A1(n70), .A2(i_data_bus[50]), .ZN(n62) );
  ND2OPTIBD1BWP30P140LVT U65 ( .A1(n64), .A2(n63), .ZN(N111) );
  ND2OPTIBD1BWP30P140LVT U66 ( .A1(n1), .A2(i_data_bus[19]), .ZN(n63) );
  ND2D1BWP30P140LVT U67 ( .A1(n70), .A2(i_data_bus[51]), .ZN(n64) );
  ND2OPTIBD1BWP30P140LVT U68 ( .A1(n66), .A2(n65), .ZN(N112) );
  ND2OPTIBD1BWP30P140LVT U69 ( .A1(n1), .A2(i_data_bus[20]), .ZN(n65) );
  ND2D1BWP30P140LVT U70 ( .A1(n70), .A2(i_data_bus[52]), .ZN(n66) );
  ND2OPTIBD1BWP30P140LVT U71 ( .A1(n68), .A2(n67), .ZN(N113) );
  ND2OPTIBD1BWP30P140LVT U72 ( .A1(n1), .A2(i_data_bus[21]), .ZN(n67) );
  ND2D1BWP30P140LVT U73 ( .A1(n70), .A2(i_data_bus[53]), .ZN(n68) );
  IND2D1BWP30P140LVT U74 ( .A1(n2), .B1(n15), .ZN(N114) );
  ND2OPTIBD1BWP30P140LVT U75 ( .A1(n1), .A2(i_data_bus[22]), .ZN(n15) );
  IND2D1BWP30P140LVT U76 ( .A1(n3), .B1(n16), .ZN(N115) );
  ND2OPTIBD1BWP30P140LVT U77 ( .A1(n1), .A2(i_data_bus[23]), .ZN(n16) );
  IND2D1BWP30P140LVT U78 ( .A1(n4), .B1(n17), .ZN(N116) );
  ND2OPTIBD1BWP30P140LVT U79 ( .A1(n1), .A2(i_data_bus[24]), .ZN(n17) );
  IND2D1BWP30P140LVT U80 ( .A1(n5), .B1(n18), .ZN(N117) );
  ND2OPTIBD1BWP30P140LVT U81 ( .A1(n1), .A2(i_data_bus[25]), .ZN(n18) );
  IND2D1BWP30P140LVT U82 ( .A1(n6), .B1(n19), .ZN(N118) );
  ND2OPTIBD1BWP30P140LVT U83 ( .A1(n1), .A2(i_data_bus[26]), .ZN(n19) );
  IND2D1BWP30P140LVT U84 ( .A1(n7), .B1(n20), .ZN(N119) );
  ND2OPTIBD1BWP30P140LVT U85 ( .A1(n1), .A2(i_data_bus[27]), .ZN(n20) );
  IND2D1BWP30P140LVT U86 ( .A1(n8), .B1(n21), .ZN(N120) );
  ND2OPTIBD1BWP30P140LVT U87 ( .A1(n1), .A2(i_data_bus[28]), .ZN(n21) );
  IND2D1BWP30P140LVT U88 ( .A1(n9), .B1(n22), .ZN(N121) );
  ND2OPTIBD1BWP30P140LVT U89 ( .A1(n1), .A2(i_data_bus[29]), .ZN(n22) );
  IND2D1BWP30P140LVT U90 ( .A1(n10), .B1(n23), .ZN(N122) );
  ND2OPTIBD1BWP30P140LVT U91 ( .A1(n1), .A2(i_data_bus[30]), .ZN(n23) );
  IND2D1BWP30P140LVT U92 ( .A1(n11), .B1(n24), .ZN(N123) );
  ND2OPTIBD1BWP30P140LVT U93 ( .A1(n1), .A2(i_data_bus[31]), .ZN(n24) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n70), .A2(i_data_bus[54]), .Z(n2) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n70), .A2(i_data_bus[55]), .Z(n3) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n70), .A2(i_data_bus[56]), .Z(n4) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n70), .A2(i_data_bus[57]), .Z(n5) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n70), .A2(i_data_bus[58]), .Z(n6) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n70), .A2(i_data_bus[59]), .Z(n7) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n70), .A2(i_data_bus[60]), .Z(n8) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n70), .A2(i_data_bus[61]), .Z(n9) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n70), .A2(i_data_bus[62]), .Z(n10) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n70), .A2(i_data_bus[63]), .Z(n11) );
  ND3D1BWP30P140LVT U104 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n12)
         );
  NR2D1BWP30P140LVT U105 ( .A1(n12), .A2(rst), .ZN(n13) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_53 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_53 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_54 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n5), .Z(n1) );
  NR2OPTPAD1BWP30P140LVT U4 ( .A1(i_cmd[0]), .A2(n3), .ZN(n6) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(i_valid[0]), .A2(n2), .ZN(n3) );
  INR2D1BWP30P140LVT U6 ( .A1(i_en), .B1(rst), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n4) );
  NR2D1BWP30P140LVT U8 ( .A1(n4), .A2(rst), .ZN(n5) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_54 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_54 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_9 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_54 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_53 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_52 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_51 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_50 o_data_high ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_49 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_55 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  NR2D1BWP30P140LVT U3 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_55 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_55 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_56 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_56 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_56 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_57 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  NR3D0P7BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n1) );
  NR3D0P7BWP30P140LVT U4 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U36 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(i_data_bus[31]), .Z(N123) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_57 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_57 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_58 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  IND2D1BWP30P140LVT U3 ( .A1(n1), .B1(i_valid[0]), .ZN(n2) );
  INVD1BWP30P140LVT U4 ( .I(i_en), .ZN(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  NR3D1P5BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n6) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  BUFFD2BWP30P140LVT U8 ( .I(n4), .Z(n5) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n5), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n5), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n5), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n5), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n5), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n5), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n5), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n5), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n5), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n5), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n5), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n5), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n5), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n5), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n5), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n5), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n5), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n5), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n5), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n5), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n5), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n5), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n5), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n5), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n5), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n5), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n5), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n5), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n5), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n5), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n5), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n5), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n5), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_58 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_58 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_59 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3OPTPAD2BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  NR2D1BWP30P140LVT U4 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U5 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U8 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_59 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_59 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_60 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3OPTPAD2BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  NR2D1BWP30P140LVT U4 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U5 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U8 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_60 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_60 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_10 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_60 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_59 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_58 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_57 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_56 o_data_high ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_55 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_61 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  NR2D1BWP30P140LVT U3 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_61 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_61 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_62 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_62 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_62 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_63 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2D1BWP30P140LVT U36 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_63 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_63 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_64 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_64 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_64 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_65 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_65 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_65 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_66 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_66 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_66 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_11 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_66 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_65 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_64 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_63 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_62 o_data_high ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_61 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_67 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2OPTPAD1BWP30P140LVT U3 ( .A1(i_cmd[0]), .A2(n3), .ZN(n6) );
  BUFFD2BWP30P140LVT U4 ( .I(n5), .Z(n1) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(i_valid[0]), .A2(n2), .ZN(n3) );
  INR2D1BWP30P140LVT U6 ( .A1(i_en), .B1(rst), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n4) );
  NR2D1BWP30P140LVT U8 ( .A1(n4), .A2(rst), .ZN(n5) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_67 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_67 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_68 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n5), .Z(n1) );
  INVD2BWP30P140LVT U4 ( .I(n3), .ZN(n6) );
  OR3D1BWP30P140LVT U5 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .Z(n3) );
  ND2D1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n4) );
  NR2D1BWP30P140LVT U8 ( .A1(n4), .A2(rst), .ZN(n5) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_68 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_68 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_69 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2D1BWP30P140LVT U24 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U36 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_69 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_69 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_70 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n5), .Z(n1) );
  NR2OPTPAD1BWP30P140LVT U4 ( .A1(i_cmd[0]), .A2(n3), .ZN(n6) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(i_valid[0]), .A2(n2), .ZN(n3) );
  INR2D1BWP30P140LVT U6 ( .A1(i_en), .B1(rst), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n4) );
  NR2D1BWP30P140LVT U8 ( .A1(n4), .A2(rst), .ZN(n5) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_70 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_70 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_71 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  CKBD1BWP30P140LVT U3 ( .I(n35), .Z(n77) );
  NR3D1P5BWP30P140LVT U4 ( .A1(n19), .A2(rst), .A3(i_cmd[0]), .ZN(n1) );
  IND2D1BWP30P140LVT U5 ( .A1(n40), .B1(n41), .ZN(N96) );
  IND2D1BWP30P140LVT U6 ( .A1(n38), .B1(n39), .ZN(N93) );
  IND2D1BWP30P140LVT U7 ( .A1(n36), .B1(n37), .ZN(N92) );
  IND2D1BWP30P140LVT U8 ( .A1(n42), .B1(n43), .ZN(N97) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n77), .A2(i_data_bus[37]), .Z(n42) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n77), .A2(i_data_bus[36]), .Z(n40) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n77), .A2(i_data_bus[33]), .Z(n38) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n77), .A2(i_data_bus[32]), .Z(n36) );
  NR2D1BWP30P140LVT U13 ( .A1(n18), .A2(rst), .ZN(n35) );
  CKBD1BWP30P140LVT U14 ( .I(n35), .Z(n83) );
  IND2D1BWP30P140LVT U15 ( .A1(n83), .B1(n82), .ZN(N91) );
  INVD1BWP30P140LVT U16 ( .I(n1), .ZN(n82) );
  ND2D1BWP30P140LVT U17 ( .A1(n1), .A2(i_data_bus[2]), .ZN(n20) );
  ND2D1BWP30P140LVT U18 ( .A1(n1), .A2(i_data_bus[3]), .ZN(n21) );
  ND2D1BWP30P140LVT U19 ( .A1(n1), .A2(i_data_bus[6]), .ZN(n22) );
  ND2D1BWP30P140LVT U20 ( .A1(n1), .A2(i_data_bus[7]), .ZN(n23) );
  ND2D1BWP30P140LVT U21 ( .A1(n1), .A2(i_data_bus[10]), .ZN(n24) );
  ND2D1BWP30P140LVT U22 ( .A1(n1), .A2(i_data_bus[11]), .ZN(n25) );
  ND2D1BWP30P140LVT U23 ( .A1(n1), .A2(i_data_bus[14]), .ZN(n26) );
  ND2D1BWP30P140LVT U24 ( .A1(n1), .A2(i_data_bus[15]), .ZN(n27) );
  ND2D1BWP30P140LVT U25 ( .A1(n1), .A2(i_data_bus[18]), .ZN(n28) );
  ND2D1BWP30P140LVT U26 ( .A1(n1), .A2(i_data_bus[19]), .ZN(n29) );
  ND2D1BWP30P140LVT U27 ( .A1(n1), .A2(i_data_bus[22]), .ZN(n30) );
  ND2D1BWP30P140LVT U28 ( .A1(n1), .A2(i_data_bus[23]), .ZN(n31) );
  ND2D1BWP30P140LVT U29 ( .A1(n1), .A2(i_data_bus[26]), .ZN(n32) );
  ND2D1BWP30P140LVT U30 ( .A1(n1), .A2(i_data_bus[27]), .ZN(n33) );
  ND2D1BWP30P140LVT U31 ( .A1(n1), .A2(i_data_bus[30]), .ZN(n34) );
  IND2D1BWP30P140LVT U32 ( .A1(n2), .B1(n81), .ZN(N123) );
  ND2D1BWP30P140LVT U33 ( .A1(n1), .A2(i_data_bus[31]), .ZN(n81) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n83), .A2(i_data_bus[63]), .Z(n2) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n83), .A2(i_data_bus[34]), .Z(n3) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n83), .A2(i_data_bus[35]), .Z(n4) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n83), .A2(i_data_bus[38]), .Z(n5) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n83), .A2(i_data_bus[39]), .Z(n6) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n83), .A2(i_data_bus[42]), .Z(n7) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n83), .A2(i_data_bus[43]), .Z(n8) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n83), .A2(i_data_bus[46]), .Z(n9) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n83), .A2(i_data_bus[47]), .Z(n10) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n83), .A2(i_data_bus[50]), .Z(n11) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n83), .A2(i_data_bus[51]), .Z(n12) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n83), .A2(i_data_bus[54]), .Z(n13) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n83), .A2(i_data_bus[55]), .Z(n14) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n83), .A2(i_data_bus[58]), .Z(n15) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n83), .A2(i_data_bus[59]), .Z(n16) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n83), .A2(i_data_bus[62]), .Z(n17) );
  ND3D1BWP30P140LVT U50 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n18)
         );
  ND2OPTIBD1BWP30P140LVT U51 ( .A1(i_en), .A2(i_valid[0]), .ZN(n19) );
  IND2D1BWP30P140LVT U52 ( .A1(n3), .B1(n20), .ZN(N94) );
  IND2D1BWP30P140LVT U53 ( .A1(n4), .B1(n21), .ZN(N95) );
  IND2D1BWP30P140LVT U54 ( .A1(n5), .B1(n22), .ZN(N98) );
  IND2D1BWP30P140LVT U55 ( .A1(n6), .B1(n23), .ZN(N99) );
  IND2D1BWP30P140LVT U56 ( .A1(n7), .B1(n24), .ZN(N102) );
  IND2D1BWP30P140LVT U57 ( .A1(n8), .B1(n25), .ZN(N103) );
  IND2D1BWP30P140LVT U58 ( .A1(n9), .B1(n26), .ZN(N106) );
  IND2D1BWP30P140LVT U59 ( .A1(n10), .B1(n27), .ZN(N107) );
  IND2D1BWP30P140LVT U60 ( .A1(n11), .B1(n28), .ZN(N110) );
  IND2D1BWP30P140LVT U61 ( .A1(n12), .B1(n29), .ZN(N111) );
  IND2D1BWP30P140LVT U62 ( .A1(n13), .B1(n30), .ZN(N114) );
  IND2D1BWP30P140LVT U63 ( .A1(n14), .B1(n31), .ZN(N115) );
  IND2D1BWP30P140LVT U64 ( .A1(n15), .B1(n32), .ZN(N118) );
  IND2D1BWP30P140LVT U65 ( .A1(n16), .B1(n33), .ZN(N119) );
  IND2D1BWP30P140LVT U66 ( .A1(n17), .B1(n34), .ZN(N122) );
  ND2D1BWP30P140LVT U67 ( .A1(n1), .A2(i_data_bus[0]), .ZN(n37) );
  ND2D1BWP30P140LVT U68 ( .A1(n1), .A2(i_data_bus[1]), .ZN(n39) );
  ND2D1BWP30P140LVT U69 ( .A1(n1), .A2(i_data_bus[4]), .ZN(n41) );
  ND2D1BWP30P140LVT U70 ( .A1(n1), .A2(i_data_bus[5]), .ZN(n43) );
  ND2D1BWP30P140LVT U71 ( .A1(n77), .A2(i_data_bus[40]), .ZN(n44) );
  INVD1BWP30P140LVT U72 ( .I(n44), .ZN(n46) );
  ND2D1BWP30P140LVT U73 ( .A1(n1), .A2(i_data_bus[8]), .ZN(n45) );
  IND2D1BWP30P140LVT U74 ( .A1(n46), .B1(n45), .ZN(N100) );
  ND2D1BWP30P140LVT U75 ( .A1(n77), .A2(i_data_bus[41]), .ZN(n47) );
  INVD1BWP30P140LVT U76 ( .I(n47), .ZN(n49) );
  ND2D1BWP30P140LVT U77 ( .A1(n1), .A2(i_data_bus[9]), .ZN(n48) );
  IND2D1BWP30P140LVT U78 ( .A1(n49), .B1(n48), .ZN(N101) );
  ND2D1BWP30P140LVT U79 ( .A1(n77), .A2(i_data_bus[44]), .ZN(n50) );
  INVD1BWP30P140LVT U80 ( .I(n50), .ZN(n52) );
  ND2D1BWP30P140LVT U81 ( .A1(n1), .A2(i_data_bus[12]), .ZN(n51) );
  IND2D1BWP30P140LVT U82 ( .A1(n52), .B1(n51), .ZN(N104) );
  ND2D1BWP30P140LVT U83 ( .A1(n77), .A2(i_data_bus[45]), .ZN(n53) );
  INVD1BWP30P140LVT U84 ( .I(n53), .ZN(n55) );
  ND2D1BWP30P140LVT U85 ( .A1(n1), .A2(i_data_bus[13]), .ZN(n54) );
  IND2D1BWP30P140LVT U86 ( .A1(n55), .B1(n54), .ZN(N105) );
  ND2D1BWP30P140LVT U87 ( .A1(n77), .A2(i_data_bus[48]), .ZN(n56) );
  INVD1BWP30P140LVT U88 ( .I(n56), .ZN(n58) );
  ND2D1BWP30P140LVT U89 ( .A1(n1), .A2(i_data_bus[16]), .ZN(n57) );
  IND2D1BWP30P140LVT U90 ( .A1(n58), .B1(n57), .ZN(N108) );
  ND2D1BWP30P140LVT U91 ( .A1(n77), .A2(i_data_bus[49]), .ZN(n59) );
  INVD1BWP30P140LVT U92 ( .I(n59), .ZN(n61) );
  ND2D1BWP30P140LVT U93 ( .A1(n1), .A2(i_data_bus[17]), .ZN(n60) );
  IND2D1BWP30P140LVT U94 ( .A1(n61), .B1(n60), .ZN(N109) );
  ND2D1BWP30P140LVT U95 ( .A1(n77), .A2(i_data_bus[52]), .ZN(n62) );
  INVD1BWP30P140LVT U96 ( .I(n62), .ZN(n64) );
  ND2D1BWP30P140LVT U97 ( .A1(n1), .A2(i_data_bus[20]), .ZN(n63) );
  IND2D1BWP30P140LVT U98 ( .A1(n64), .B1(n63), .ZN(N112) );
  ND2D1BWP30P140LVT U99 ( .A1(n77), .A2(i_data_bus[53]), .ZN(n65) );
  INVD1BWP30P140LVT U100 ( .I(n65), .ZN(n67) );
  ND2D1BWP30P140LVT U101 ( .A1(n1), .A2(i_data_bus[21]), .ZN(n66) );
  IND2D1BWP30P140LVT U102 ( .A1(n67), .B1(n66), .ZN(N113) );
  ND2D1BWP30P140LVT U103 ( .A1(n77), .A2(i_data_bus[56]), .ZN(n68) );
  INVD1BWP30P140LVT U104 ( .I(n68), .ZN(n70) );
  ND2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[24]), .ZN(n69) );
  IND2D1BWP30P140LVT U106 ( .A1(n70), .B1(n69), .ZN(N116) );
  ND2D1BWP30P140LVT U107 ( .A1(n77), .A2(i_data_bus[57]), .ZN(n71) );
  INVD1BWP30P140LVT U108 ( .I(n71), .ZN(n73) );
  ND2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[25]), .ZN(n72) );
  IND2D1BWP30P140LVT U110 ( .A1(n73), .B1(n72), .ZN(N117) );
  ND2D1BWP30P140LVT U111 ( .A1(n77), .A2(i_data_bus[60]), .ZN(n74) );
  INVD1BWP30P140LVT U112 ( .I(n74), .ZN(n76) );
  ND2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[28]), .ZN(n75) );
  IND2D1BWP30P140LVT U114 ( .A1(n76), .B1(n75), .ZN(N120) );
  ND2D1BWP30P140LVT U115 ( .A1(n77), .A2(i_data_bus[61]), .ZN(n78) );
  INVD1BWP30P140LVT U116 ( .I(n78), .ZN(n80) );
  ND2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[29]), .ZN(n79) );
  IND2D1BWP30P140LVT U118 ( .A1(n80), .B1(n79), .ZN(N121) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_71 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_71 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_72 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n5), .Z(n1) );
  NR2OPTPAD1BWP30P140LVT U4 ( .A1(i_cmd[0]), .A2(n3), .ZN(n6) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(i_valid[0]), .A2(n2), .ZN(n3) );
  INR2D1BWP30P140LVT U6 ( .A1(i_en), .B1(rst), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n4) );
  NR2D1BWP30P140LVT U8 ( .A1(n4), .A2(rst), .ZN(n5) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_72 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_72 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_12 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_72 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_71 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_70 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_69 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_68 o_data_high ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_67 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_73 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  NR3OPTPAD2BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_73 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_73 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_74 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n33, n34, n35,
         n36, n37;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  ND2OPTIBD1BWP30P140LVT U3 ( .A1(i_en), .A2(i_valid[0]), .ZN(n33) );
  NR2D1BWP30P140LVT U4 ( .A1(n34), .A2(rst), .ZN(n35) );
  NR3D1P5BWP30P140LVT U5 ( .A1(n33), .A2(i_cmd[0]), .A3(rst), .ZN(n37) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n34)
         );
  BUFFD2BWP30P140LVT U7 ( .I(n35), .Z(n36) );
  AO22D1BWP30P140LVT U8 ( .A1(n37), .A2(i_data_bus[0]), .B1(n36), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n37), .A2(i_data_bus[1]), .B1(n36), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n37), .A2(i_data_bus[2]), .B1(n36), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n37), .A2(i_data_bus[3]), .B1(n36), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n37), .A2(i_data_bus[4]), .B1(n36), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n37), .A2(i_data_bus[5]), .B1(n36), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n37), .A2(i_data_bus[6]), .B1(n36), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n37), .A2(i_data_bus[7]), .B1(n36), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n37), .A2(i_data_bus[8]), .B1(n36), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n37), .A2(i_data_bus[9]), .B1(n36), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n37), .A2(i_data_bus[10]), .B1(n36), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n37), .A2(i_data_bus[11]), .B1(n36), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n37), .A2(i_data_bus[12]), .B1(n36), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n37), .A2(i_data_bus[13]), .B1(n36), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n37), .A2(i_data_bus[14]), .B1(n36), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n37), .A2(i_data_bus[15]), .B1(n36), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n37), .A2(i_data_bus[16]), .B1(n36), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n37), .A2(i_data_bus[17]), .B1(n36), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n37), .A2(i_data_bus[18]), .B1(n36), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n37), .A2(i_data_bus[19]), .B1(n36), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n37), .A2(i_data_bus[20]), .B1(n36), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n37), .A2(i_data_bus[21]), .B1(n36), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n37), .A2(i_data_bus[22]), .B1(n36), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n37), .A2(i_data_bus[23]), .B1(n36), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n37), .A2(i_data_bus[24]), .B1(n36), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n37), .A2(i_data_bus[25]), .B1(n36), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n37), .A2(i_data_bus[26]), .B1(n36), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n37), .A2(i_data_bus[27]), .B1(n36), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n37), .A2(i_data_bus[28]), .B1(n36), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n37), .A2(i_data_bus[29]), .B1(n36), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n37), .A2(i_data_bus[30]), .B1(n36), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n37), .A2(i_data_bus[31]), .B1(n36), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n37), .A2(n36), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_74 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_74 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_75 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  ND2D1BWP30P140LVT U9 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3D1P5BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U36 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_75 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_75 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_76 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n5), .Z(n1) );
  NR3D1P5BWP30P140LVT U4 ( .A1(n3), .A2(i_cmd[0]), .A3(rst), .ZN(n2) );
  NR2D1BWP30P140LVT U5 ( .A1(n4), .A2(rst), .ZN(n5) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n3) );
  NR3D1P5BWP30P140LVT U7 ( .A1(n3), .A2(i_cmd[0]), .A3(rst), .ZN(n6) );
  ND3D1BWP30P140LVT U8 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n4) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n2), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n2), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n2), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n2), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n2), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n2), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n2), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n2), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n2), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n2), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n2), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n2), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n2), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n2), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n2), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n2), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_76 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_76 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_77 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n34, n35,
         n36, n37;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n34), .A2(i_cmd[0]), .A3(rst), .ZN(n37) );
  BUFFD2BWP30P140LVT U4 ( .I(n36), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n35), .A2(rst), .ZN(n36) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n34) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n35)
         );
  AO22D1BWP30P140LVT U8 ( .A1(n37), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n37), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n37), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n37), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n37), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n37), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n37), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n37), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n37), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n37), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n37), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n37), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n37), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n37), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n37), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n37), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n37), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n37), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n37), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n37), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n37), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n37), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n37), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n37), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n37), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n37), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n37), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n37), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n37), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n37), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n37), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n37), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n37), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_77 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_77 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_78 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n34, n35,
         n36, n37;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n34), .A2(i_cmd[0]), .A3(rst), .ZN(n37) );
  BUFFD2BWP30P140LVT U4 ( .I(n36), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n35), .A2(rst), .ZN(n36) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n34) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n35)
         );
  AO22D1BWP30P140LVT U8 ( .A1(n37), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n37), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n37), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n37), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n37), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n37), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n37), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n37), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n37), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n37), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n37), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n37), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n37), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n37), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n37), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n37), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n37), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n37), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n37), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n37), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n37), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n37), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n37), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n37), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n37), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n37), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n37), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n37), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n37), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n37), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n37), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n37), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n37), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_78 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_78 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_13 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_78 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_77 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_76 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_75 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_74 o_data_high ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_73 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  CKAN2D1BWP30P140LVT U2 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
  TIELBWP30P140LVT U3 ( .ZN(n_Logic0_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_79 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_79 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_79 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_80 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_80 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_80 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_81 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2OPTIBD1BWP30P140LVT U36 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_81 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_81 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_82 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_82 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_82 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_83 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_83 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_83 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_84 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_84 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_84 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_14 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_84 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_83 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_82 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_81 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_80 o_data_high ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_79 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_85 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n5), .Z(n1) );
  INVD2BWP30P140LVT U4 ( .I(n3), .ZN(n6) );
  OR3D1BWP30P140LVT U5 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .Z(n3) );
  ND2D1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n4) );
  NR2D1BWP30P140LVT U8 ( .A1(n4), .A2(rst), .ZN(n5) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n5), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_85 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_85 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_86 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n5), .Z(n1) );
  INVD2BWP30P140LVT U4 ( .I(n3), .ZN(n6) );
  OR3D1BWP30P140LVT U5 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .Z(n3) );
  ND2D1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n4) );
  NR2D1BWP30P140LVT U8 ( .A1(n4), .A2(rst), .ZN(n5) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n5), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_86 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_86 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_87 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  NR3D1P5BWP30P140LVT U3 ( .A1(i_cmd[0]), .A2(n1), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2D1BWP30P140LVT U24 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U36 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_87 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_87 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_88 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n5), .Z(n1) );
  INVD2BWP30P140LVT U4 ( .I(n3), .ZN(n6) );
  OR3D1BWP30P140LVT U5 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .Z(n3) );
  ND2D1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n4) );
  NR2D1BWP30P140LVT U8 ( .A1(n4), .A2(rst), .ZN(n5) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n5), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_88 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_88 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_89 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n5), .Z(n1) );
  INVD2BWP30P140LVT U4 ( .I(n3), .ZN(n6) );
  OR3D1BWP30P140LVT U5 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .Z(n3) );
  ND2D1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n4) );
  NR2D1BWP30P140LVT U8 ( .A1(n4), .A2(rst), .ZN(n5) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n5), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_89 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_89 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_90 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n5), .Z(n1) );
  INVD2BWP30P140LVT U4 ( .I(n3), .ZN(n6) );
  OR3D1BWP30P140LVT U5 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .Z(n3) );
  ND2D1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n4) );
  NR2D1BWP30P140LVT U8 ( .A1(n4), .A2(rst), .ZN(n5) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n5), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_90 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_90 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_15 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_90 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_89 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_88 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_87 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_86 o_data_high ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_85 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_91 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_91 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_91 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_92 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_92 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_92 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_93 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2D1BWP30P140LVT U36 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_93 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_93 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_94 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n23), .Z(n22) );
  INVD1BWP30P140LVT U4 ( .I(n22), .ZN(n1) );
  INVD1BWP30P140LVT U5 ( .I(n24), .ZN(n2) );
  NR2D1BWP30P140LVT U6 ( .A1(n5), .A2(rst), .ZN(n23) );
  IND2D1BWP30P140LVT U7 ( .A1(n3), .B1(i_valid[0]), .ZN(n4) );
  INVD1BWP30P140LVT U8 ( .I(i_en), .ZN(n3) );
  OAI22D1BWP30P140LVT U9 ( .A1(n2), .A2(n8), .B1(n7), .B2(n6), .ZN(N118) );
  INVD1BWP30P140LVT U10 ( .I(i_data_bus[26]), .ZN(n8) );
  INVD1BWP30P140LVT U11 ( .I(i_data_bus[58]), .ZN(n6) );
  INVD1BWP30P140LVT U12 ( .I(n22), .ZN(n7) );
  OAI22D1BWP30P140LVT U13 ( .A1(n2), .A2(n11), .B1(n10), .B2(n9), .ZN(N119) );
  INVD1BWP30P140LVT U14 ( .I(i_data_bus[27]), .ZN(n11) );
  INVD1BWP30P140LVT U15 ( .I(i_data_bus[59]), .ZN(n9) );
  INVD1BWP30P140LVT U16 ( .I(n22), .ZN(n10) );
  OAI22D1BWP30P140LVT U17 ( .A1(n2), .A2(n14), .B1(n13), .B2(n12), .ZN(N120)
         );
  INVD1BWP30P140LVT U18 ( .I(i_data_bus[28]), .ZN(n14) );
  INVD1BWP30P140LVT U19 ( .I(i_data_bus[60]), .ZN(n12) );
  INVD1BWP30P140LVT U20 ( .I(n22), .ZN(n13) );
  OAI22D1BWP30P140LVT U21 ( .A1(n2), .A2(n16), .B1(n1), .B2(n15), .ZN(N121) );
  INVD1BWP30P140LVT U22 ( .I(i_data_bus[29]), .ZN(n16) );
  INVD1BWP30P140LVT U23 ( .I(i_data_bus[61]), .ZN(n15) );
  OAI22D1BWP30P140LVT U24 ( .A1(n2), .A2(n18), .B1(n1), .B2(n17), .ZN(N122) );
  INVD1BWP30P140LVT U25 ( .I(i_data_bus[30]), .ZN(n18) );
  INVD1BWP30P140LVT U26 ( .I(i_data_bus[62]), .ZN(n17) );
  OAI22D1BWP30P140LVT U27 ( .A1(n2), .A2(n21), .B1(n20), .B2(n19), .ZN(N123)
         );
  INVD1BWP30P140LVT U28 ( .I(i_data_bus[31]), .ZN(n21) );
  INVD1BWP30P140LVT U29 ( .I(i_data_bus[63]), .ZN(n19) );
  INVD1BWP30P140LVT U30 ( .I(n22), .ZN(n20) );
  NR3D1P5BWP30P140LVT U31 ( .A1(n4), .A2(i_cmd[0]), .A3(rst), .ZN(n24) );
  ND3D1BWP30P140LVT U32 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n5)
         );
  AO22D1BWP30P140LVT U33 ( .A1(n24), .A2(i_data_bus[0]), .B1(n22), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U34 ( .A1(n24), .A2(i_data_bus[1]), .B1(n22), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U35 ( .A1(n24), .A2(i_data_bus[2]), .B1(n22), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U36 ( .A1(n24), .A2(i_data_bus[3]), .B1(n22), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U37 ( .A1(n24), .A2(i_data_bus[4]), .B1(n22), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U38 ( .A1(n24), .A2(i_data_bus[5]), .B1(n22), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U39 ( .A1(n24), .A2(i_data_bus[6]), .B1(n22), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U40 ( .A1(n24), .A2(i_data_bus[7]), .B1(n22), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U41 ( .A1(n24), .A2(i_data_bus[8]), .B1(n22), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U42 ( .A1(n24), .A2(i_data_bus[9]), .B1(n22), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U43 ( .A1(n24), .A2(i_data_bus[10]), .B1(n22), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U44 ( .A1(n24), .A2(i_data_bus[11]), .B1(n22), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U45 ( .A1(n24), .A2(i_data_bus[12]), .B1(n22), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U46 ( .A1(n24), .A2(i_data_bus[13]), .B1(n22), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U47 ( .A1(n24), .A2(i_data_bus[14]), .B1(n22), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U48 ( .A1(n24), .A2(i_data_bus[15]), .B1(n22), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U49 ( .A1(n24), .A2(i_data_bus[16]), .B1(n22), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U50 ( .A1(n24), .A2(i_data_bus[17]), .B1(n22), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U51 ( .A1(n24), .A2(i_data_bus[18]), .B1(n22), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U52 ( .A1(n24), .A2(i_data_bus[19]), .B1(n22), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U53 ( .A1(n24), .A2(i_data_bus[20]), .B1(n22), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U54 ( .A1(n24), .A2(i_data_bus[21]), .B1(n22), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U55 ( .A1(n24), .A2(i_data_bus[22]), .B1(n22), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U56 ( .A1(n24), .A2(i_data_bus[23]), .B1(n22), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U57 ( .A1(n24), .A2(i_data_bus[24]), .B1(n22), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U58 ( .A1(n24), .A2(i_data_bus[25]), .B1(n22), .B2(
        i_data_bus[57]), .Z(N117) );
  OR2D1BWP30P140LVT U59 ( .A1(n24), .A2(n23), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_94 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_94 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_95 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  CKBD1BWP30P140LVT U3 ( .I(n5), .Z(n4) );
  NR3OPTPAD2BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n6) );
  CKBD1BWP30P140LVT U5 ( .I(n5), .Z(n3) );
  NR2D1BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n5) );
  AO22D1BWP30P140LVT U7 ( .A1(n6), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  ND2OPTIBD1BWP30P140LVT U8 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U9 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_95 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_95 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_96 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  CKBD1BWP30P140LVT U3 ( .I(n5), .Z(n4) );
  NR3OPTPAD2BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n6) );
  CKBD1BWP30P140LVT U5 ( .I(n5), .Z(n3) );
  NR2D1BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n5) );
  AO22D1BWP30P140LVT U7 ( .A1(n6), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  ND2OPTIBD1BWP30P140LVT U8 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U9 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_96 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_96 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_16 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_96 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_95 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_94 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_93 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_92 o_data_high ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_91 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_97 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_97 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_97 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_98 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_98 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_98 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_99 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U36 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_99 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_99 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_100 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_100 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_100 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_101 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_101 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_101 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_102 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_102 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_102 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_17 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_102 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_101 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_100 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_99 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_98 o_data_high ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_97 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  AN2D2BWP30P140LVT U2 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
  TIELBWP30P140LVT U3 ( .ZN(n_Logic0_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_103 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  NR2OPTPAD1BWP30P140LVT U3 ( .A1(i_cmd[0]), .A2(n3), .ZN(n6) );
  BUFFD2BWP30P140LVT U4 ( .I(n5), .Z(n1) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(i_valid[0]), .A2(n2), .ZN(n3) );
  INR2D1BWP30P140LVT U6 ( .A1(i_en), .B1(rst), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n4) );
  NR2D1BWP30P140LVT U8 ( .A1(n4), .A2(rst), .ZN(n5) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n5), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_103 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_103 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_104 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n2), .Z(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n5), .A2(rst), .ZN(n2) );
  INVD2BWP30P140LVT U5 ( .I(n4), .ZN(n6) );
  OR3D1BWP30P140LVT U6 ( .A1(n3), .A2(i_cmd[0]), .A3(rst), .Z(n4) );
  ND2D1BWP30P140LVT U7 ( .A1(i_en), .A2(i_valid[0]), .ZN(n3) );
  ND3D1BWP30P140LVT U8 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n5) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_104 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_104 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_105 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2D1BWP30P140LVT U24 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U36 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_105 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_105 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_106 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n6) );
  BUFFD2BWP30P140LVT U4 ( .I(n2), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n5), .A2(rst), .ZN(n2) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n3) );
  NR3D0P7BWP30P140LVT U7 ( .A1(n3), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND3D1BWP30P140LVT U8 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n5) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_106 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_106 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_107 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n6) );
  BUFFD2BWP30P140LVT U4 ( .I(n2), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n5), .A2(rst), .ZN(n2) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n3) );
  NR3D0P7BWP30P140LVT U7 ( .A1(n3), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND3D1BWP30P140LVT U8 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n5) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_107 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_107 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_108 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n6) );
  BUFFD2BWP30P140LVT U4 ( .I(n2), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n5), .A2(rst), .ZN(n2) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n3) );
  NR3D0P7BWP30P140LVT U7 ( .A1(n3), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND3D1BWP30P140LVT U8 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n5) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_108 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_108 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_18 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_108 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_107 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_106 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_105 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_104 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_103 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_109 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n35,
         n36, n37;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n35), .A2(i_cmd[0]), .A3(rst), .ZN(n1) );
  BUFFD2BWP30P140LVT U4 ( .I(n37), .Z(n2) );
  NR2D1BWP30P140LVT U5 ( .A1(n36), .A2(rst), .ZN(n37) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n35) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n36)
         );
  AO22D1BWP30P140LVT U8 ( .A1(n1), .A2(i_data_bus[0]), .B1(n2), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n1), .A2(i_data_bus[1]), .B1(n2), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n1), .A2(i_data_bus[2]), .B1(n2), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n1), .A2(i_data_bus[3]), .B1(n2), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n1), .A2(i_data_bus[4]), .B1(n2), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n1), .A2(i_data_bus[5]), .B1(n2), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n1), .A2(i_data_bus[6]), .B1(n2), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n1), .A2(i_data_bus[7]), .B1(n2), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n1), .A2(i_data_bus[8]), .B1(n2), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n1), .A2(i_data_bus[9]), .B1(n2), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n1), .A2(i_data_bus[10]), .B1(n2), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n1), .A2(i_data_bus[11]), .B1(n2), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n1), .A2(i_data_bus[12]), .B1(n2), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n1), .A2(i_data_bus[13]), .B1(n2), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n1), .A2(i_data_bus[14]), .B1(n2), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n1), .A2(i_data_bus[15]), .B1(n2), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n1), .A2(i_data_bus[16]), .B1(n2), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n1), .A2(i_data_bus[17]), .B1(n2), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n1), .A2(i_data_bus[18]), .B1(n2), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n1), .A2(i_data_bus[19]), .B1(n2), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n1), .A2(i_data_bus[20]), .B1(n2), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n1), .A2(i_data_bus[21]), .B1(n2), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n1), .A2(i_data_bus[22]), .B1(n2), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n1), .A2(i_data_bus[23]), .B1(n2), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n1), .A2(i_data_bus[24]), .B1(n2), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n1), .A2(i_data_bus[25]), .B1(n2), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n1), .A2(i_data_bus[26]), .B1(n2), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n1), .A2(i_data_bus[27]), .B1(n2), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n1), .A2(i_data_bus[28]), .B1(n2), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n1), .A2(i_data_bus[29]), .B1(n2), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n1), .A2(i_data_bus[30]), .B1(n2), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n1), .A2(i_data_bus[31]), .B1(n2), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n1), .A2(n37), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_109 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_109 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_110 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n36,
         n37, n38, n39;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n36), .A2(i_cmd[0]), .A3(rst), .ZN(n39) );
  BUFFD2BWP30P140LVT U4 ( .I(n38), .Z(n1) );
  ND2D1BWP30P140LVT U5 ( .A1(n2), .A2(n3), .ZN(N117) );
  ND2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_data_bus[57]), .ZN(n2) );
  ND2D1BWP30P140LVT U7 ( .A1(n39), .A2(i_data_bus[25]), .ZN(n3) );
  NR2D1BWP30P140LVT U8 ( .A1(n37), .A2(rst), .ZN(n38) );
  ND2OPTIBD1BWP30P140LVT U9 ( .A1(i_en), .A2(i_valid[0]), .ZN(n36) );
  ND3D1BWP30P140LVT U10 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n37)
         );
  AO22D1BWP30P140LVT U11 ( .A1(n39), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U12 ( .A1(n39), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U13 ( .A1(n39), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U14 ( .A1(n39), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U15 ( .A1(n39), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U16 ( .A1(n39), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U17 ( .A1(n39), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U18 ( .A1(n39), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U19 ( .A1(n39), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U20 ( .A1(n39), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U21 ( .A1(n39), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U22 ( .A1(n39), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U23 ( .A1(n39), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U24 ( .A1(n39), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U25 ( .A1(n39), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U26 ( .A1(n39), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U27 ( .A1(n39), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U28 ( .A1(n39), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U29 ( .A1(n39), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U30 ( .A1(n39), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U31 ( .A1(n39), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U32 ( .A1(n39), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U33 ( .A1(n39), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U34 ( .A1(n39), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U35 ( .A1(n39), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U36 ( .A1(n39), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U37 ( .A1(n39), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U38 ( .A1(n39), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U39 ( .A1(n39), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U40 ( .A1(n39), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U41 ( .A1(n39), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U42 ( .A1(n39), .A2(n38), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_110 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_110 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_111 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2D1BWP30P140LVT U3 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3D1P5BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U36 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_111 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_111 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_112 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_112 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_112 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_113 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n34, n35,
         n36;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n34), .A2(i_cmd[0]), .A3(rst), .ZN(n1) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n34) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n35)
         );
  NR2D3BWP30P140LVT U6 ( .A1(n35), .A2(rst), .ZN(n36) );
  AO22D1BWP30P140LVT U7 ( .A1(n1), .A2(i_data_bus[0]), .B1(n36), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n1), .A2(i_data_bus[1]), .B1(n36), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n1), .A2(i_data_bus[2]), .B1(n36), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n1), .A2(i_data_bus[3]), .B1(n36), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n1), .A2(i_data_bus[4]), .B1(n36), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n1), .A2(i_data_bus[5]), .B1(n36), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n1), .A2(i_data_bus[6]), .B1(n36), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n1), .A2(i_data_bus[7]), .B1(n36), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n1), .A2(i_data_bus[8]), .B1(n36), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n1), .A2(i_data_bus[9]), .B1(n36), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n1), .A2(i_data_bus[10]), .B1(n36), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n1), .A2(i_data_bus[11]), .B1(n36), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n1), .A2(i_data_bus[12]), .B1(n36), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n1), .A2(i_data_bus[13]), .B1(n36), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n1), .A2(i_data_bus[14]), .B1(n36), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n1), .A2(i_data_bus[15]), .B1(n36), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n1), .A2(i_data_bus[16]), .B1(n36), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n1), .A2(i_data_bus[17]), .B1(n36), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n1), .A2(i_data_bus[18]), .B1(n36), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n1), .A2(i_data_bus[19]), .B1(n36), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n1), .A2(i_data_bus[20]), .B1(n36), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n1), .A2(i_data_bus[21]), .B1(n36), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n1), .A2(i_data_bus[22]), .B1(n36), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n1), .A2(i_data_bus[23]), .B1(n36), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n1), .A2(i_data_bus[24]), .B1(n36), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n1), .A2(i_data_bus[25]), .B1(n36), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n1), .A2(i_data_bus[26]), .B1(n36), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n1), .A2(i_data_bus[27]), .B1(n36), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n1), .A2(i_data_bus[28]), .B1(n36), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n1), .A2(i_data_bus[29]), .B1(n36), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n1), .A2(i_data_bus[30]), .B1(n36), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n1), .A2(i_data_bus[31]), .B1(n36), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n1), .A2(n36), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_113 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_113 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_114 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n33, n34, n35,
         n36;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFD2BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n33), .A2(i_cmd[0]), .A3(rst), .ZN(n36) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n33) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n34)
         );
  NR2D3BWP30P140LVT U6 ( .A1(n34), .A2(rst), .ZN(n35) );
  AO22D1BWP30P140LVT U7 ( .A1(n36), .A2(i_data_bus[0]), .B1(n35), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n36), .A2(i_data_bus[1]), .B1(n35), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n36), .A2(i_data_bus[2]), .B1(n35), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n36), .A2(i_data_bus[3]), .B1(n35), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n36), .A2(i_data_bus[4]), .B1(n35), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n36), .A2(i_data_bus[5]), .B1(n35), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n36), .A2(i_data_bus[6]), .B1(n35), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n36), .A2(i_data_bus[7]), .B1(n35), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n36), .A2(i_data_bus[8]), .B1(n35), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n36), .A2(i_data_bus[9]), .B1(n35), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n36), .A2(i_data_bus[10]), .B1(n35), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n36), .A2(i_data_bus[11]), .B1(n35), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n36), .A2(i_data_bus[12]), .B1(n35), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n36), .A2(i_data_bus[13]), .B1(n35), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n36), .A2(i_data_bus[14]), .B1(n35), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n36), .A2(i_data_bus[15]), .B1(n35), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n36), .A2(i_data_bus[16]), .B1(n35), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n36), .A2(i_data_bus[17]), .B1(n35), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n36), .A2(i_data_bus[18]), .B1(n35), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n36), .A2(i_data_bus[19]), .B1(n35), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n36), .A2(i_data_bus[20]), .B1(n35), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n36), .A2(i_data_bus[21]), .B1(n35), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n36), .A2(i_data_bus[22]), .B1(n35), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n36), .A2(i_data_bus[23]), .B1(n35), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n36), .A2(i_data_bus[24]), .B1(n35), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n36), .A2(i_data_bus[25]), .B1(n35), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n36), .A2(i_data_bus[26]), .B1(n35), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n36), .A2(i_data_bus[27]), .B1(n35), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n36), .A2(i_data_bus[28]), .B1(n35), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n36), .A2(i_data_bus[29]), .B1(n35), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n36), .A2(i_data_bus[30]), .B1(n35), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n36), .A2(i_data_bus[31]), .B1(n35), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n36), .A2(n35), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_114 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_114 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_19 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_114 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_113 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_112 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_111 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_110 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_109 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_115 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_115 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_115 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_116 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D3BWP30P140LVT U3 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_116 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_116 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_117 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2D1BWP30P140LVT U36 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_117 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_117 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_118 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  IND2D1BWP30P140LVT U3 ( .A1(n1), .B1(i_valid[0]), .ZN(n2) );
  INVD1BWP30P140LVT U4 ( .I(i_en), .ZN(n1) );
  NR3D1P5BWP30P140LVT U5 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  NR2D3BWP30P140LVT U7 ( .A1(n3), .A2(rst), .ZN(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_118 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_118 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_119 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D3BWP30P140LVT U3 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_119 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_119 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_120 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2D1BWP30P140LVT U3 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U4 ( .A1(i_cmd[0]), .A2(n1), .A3(rst), .ZN(n4) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_120 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_120 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_20 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_120 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_119 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_118 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_117 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_116 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_115 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_121 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  INVD2BWP30P140LVT U3 ( .I(n3), .ZN(n5) );
  OR3D1BWP30P140LVT U4 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .Z(n3) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  AN3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .Z(n1) );
  INR2D4BWP30P140LVT U7 ( .A1(n1), .B1(rst), .ZN(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_121 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_121 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_122 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  INVD2BWP30P140LVT U3 ( .I(n3), .ZN(n5) );
  OR3D1BWP30P140LVT U4 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .Z(n3) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  AN3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .Z(n1) );
  INR2D4BWP30P140LVT U7 ( .A1(n1), .B1(rst), .ZN(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_122 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_122 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_123 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(i_cmd[0]), .A2(n1), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2D1BWP30P140LVT U24 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U36 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_123 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_123 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_124 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n4), .A2(rst), .ZN(n1) );
  INVD2BWP30P140LVT U4 ( .I(n3), .ZN(n6) );
  OR3D1BWP30P140LVT U5 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .Z(n3) );
  ND2D1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n4) );
  NR2D2BWP30P140LVT U8 ( .A1(n4), .A2(rst), .ZN(n5) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n5), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n5), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n5), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n5), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n5), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n5), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n5), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n5), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n5), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n5), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n5), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n5), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n5), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n5), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n5), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n5), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n5), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n5), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n5), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n5), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n5), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n5), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_124 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_124 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_125 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2OPTPAD2BWP30P140LVT U3 ( .A1(n3), .A2(rst), .ZN(n4) );
  INVD2BWP30P140LVT U4 ( .I(n2), .ZN(n5) );
  OR3D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .Z(n2) );
  ND2D1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_125 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_125 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_126 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2OPTPAD2BWP30P140LVT U3 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND3D1BWP30P140LVT U4 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  INVD2BWP30P140LVT U5 ( .I(n2), .ZN(n5) );
  OR3D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .Z(n2) );
  ND2D1BWP30P140LVT U7 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_126 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_126 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_21 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_126 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_125 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_124 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_123 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_122 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_121 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_127 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D3BWP30P140LVT U3 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_127 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_127 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_128 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2OPTIBD1BWP30P140LVT U3 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_128 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_128 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_129 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2D1BWP30P140LVT U36 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_129 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_129 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_130 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3OPTPAD2BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n1) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n1), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n1), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n1), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n1), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n1), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n1), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n1), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n1), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n1), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n1), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n1), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n1), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n1), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n1), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n1), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n1), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n1), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n1), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n1), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n1), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n1), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n1), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n1), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n1), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n1), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n1), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n1), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n1), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n1), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n1), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n1), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n1), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n1), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_130 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_130 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_131 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  ND2D1BWP30P140LVT U3 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U4 ( .A1(i_cmd[0]), .A2(n1), .A3(rst), .ZN(n4) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_131 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_131 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_132 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2D1BWP30P140LVT U3 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U4 ( .A1(i_cmd[0]), .A2(n1), .A3(rst), .ZN(n4) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_132 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_132 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_22 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_132 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_131 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_130 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_129 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_128 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_127 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_133 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_133 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_133 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_134 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  NR2D1BWP30P140LVT U4 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_134 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_134 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_135 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2D1BWP30P140LVT U36 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_135 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_135 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_136 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  NR2D1BWP30P140LVT U4 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_136 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_136 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_137 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  NR2D1BWP30P140LVT U4 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_137 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_137 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_138 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  NR2D1BWP30P140LVT U4 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_138 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_138 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_23 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_138 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_137 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_136 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_135 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_134 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_133 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_139 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_139 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_139 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_140 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_140 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_140 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_141 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2D1BWP30P140LVT U36 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_141 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_141 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_142 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_142 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_142 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_143 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_143 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_143 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_144 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_144 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_144 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_24 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_144 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_143 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_142 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_141 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_140 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_139 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_145 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_145 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_145 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_146 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  NR2D1BWP30P140LVT U4 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_146 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_146 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_147 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2D1BWP30P140LVT U36 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_147 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_147 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_148 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  NR2D1BWP30P140LVT U4 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_148 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_148 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_149 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  NR2D1BWP30P140LVT U4 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_149 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_149 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_150 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  NR2D1BWP30P140LVT U4 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_150 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_150 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_25 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_150 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_149 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_148 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_147 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_146 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_145 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_151 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_151 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_151 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_152 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_152 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_152 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_153 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2D1BWP30P140LVT U36 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_153 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_153 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_154 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_154 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_154 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_155 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_155 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_155 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_156 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_156 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_156 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_26 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_156 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_155 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_154 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_153 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_152 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_151 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_157 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_157 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_157 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_158 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_158 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_158 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_159 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2OPTIBD1BWP30P140LVT U36 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_159 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_159 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_160 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_160 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_160 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_161 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_161 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_161 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_162 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_162 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_162 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_27 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_162 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_161 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_160 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_159 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_158 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_157 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_163 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_163 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_163 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_164 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_164 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_164 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_165 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2D1BWP30P140LVT U36 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_165 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_165 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_166 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_166 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_166 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_167 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_167 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_167 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_168 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_168 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_168 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_28 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_168 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_167 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_166 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_165 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_164 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_163 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_169 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_169 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_169 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_170 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_170 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_170 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_171 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2D1BWP30P140LVT U36 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_171 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_171 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_172 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_172 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_172 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_173 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_173 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_173 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_174 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_174 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_174 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_29 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_174 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_173 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_172 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_171 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_170 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_169 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_175 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2D1BWP30P140LVT U3 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_175 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_175 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_176 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_176 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_176 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_177 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2D1BWP30P140LVT U36 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_177 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_177 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_178 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_178 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_178 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_179 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_179 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_179 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_180 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_180 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_180 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_30 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_180 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_179 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_178 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_177 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_176 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_175 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_181 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_181 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_181 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_182 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_182 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_182 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_183 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2D1BWP30P140LVT U36 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_183 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_183 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_184 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_184 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_184 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_185 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_185 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_185 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_186 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_186 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_186 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_31 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_186 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_185 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_184 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_183 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_182 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_181 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_187 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2D1BWP30P140LVT U3 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_187 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_187 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_188 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_188 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_188 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_189 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2D1BWP30P140LVT U36 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_189 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_189 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_190 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_190 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_190 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_191 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_191 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_191 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_192 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_192 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_192 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_32 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_192 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_191 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_190 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_189 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_188 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_187 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_193 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D3BWP30P140LVT U3 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_193 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_193 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_194 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2D1BWP30P140LVT U3 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_194 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_194 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_195 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2OPTIBD1BWP30P140LVT U36 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_195 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_195 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_196 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_196 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_196 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_197 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_197 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_197 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_198 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_198 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_198 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_33 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_198 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_197 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_196 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_195 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_194 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_193 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_199 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2D1BWP30P140LVT U3 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_199 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_199 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_200 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_200 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_200 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_201 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2D1BWP30P140LVT U36 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_201 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_201 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_202 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_202 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_202 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_203 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_203 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_203 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_204 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_204 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_204 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_34 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_204 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_203 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_202 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_201 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_200 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_199 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_205 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2D1BWP30P140LVT U3 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U4 ( .A1(i_cmd[0]), .A2(n1), .A3(rst), .ZN(n4) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_205 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_205 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_206 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2D1BWP30P140LVT U3 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_206 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_206 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_207 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U36 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_207 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_207 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_208 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_208 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_208 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_209 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_209 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_209 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_210 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_210 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_210 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_35 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_210 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_209 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_208 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_207 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_206 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_205 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  CKAN2D1BWP30P140LVT U2 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
  TIELBWP30P140LVT U3 ( .ZN(n_Logic0_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_211 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2D1BWP30P140LVT U3 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_211 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_211 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_212 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_212 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_212 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_213 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2D1BWP30P140LVT U36 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_213 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_213 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_214 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_214 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_214 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_215 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_215 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_215 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_216 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_216 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_216 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_36 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_216 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_215 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_214 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_213 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_212 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_211 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_217 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2D1BWP30P140LVT U3 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U4 ( .A1(i_cmd[0]), .A2(n1), .A3(rst), .ZN(n4) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_217 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_217 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_218 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2D1BWP30P140LVT U3 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_218 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_218 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_219 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U36 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_219 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_219 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_220 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_220 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_220 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_221 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_221 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_221 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_222 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  NR2D3BWP30P140LVT U6 ( .A1(n2), .A2(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[0]), .B1(n3), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[1]), .B1(n3), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[2]), .B1(n3), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[3]), .B1(n3), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[4]), .B1(n3), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[5]), .B1(n3), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[6]), .B1(n3), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[7]), .B1(n3), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[8]), .B1(n3), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[9]), .B1(n3), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[10]), .B1(n3), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[11]), .B1(n3), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[12]), .B1(n3), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[13]), .B1(n3), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[14]), .B1(n3), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[15]), .B1(n3), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[16]), .B1(n3), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[17]), .B1(n3), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[18]), .B1(n3), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[19]), .B1(n3), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[20]), .B1(n3), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[21]), .B1(n3), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[22]), .B1(n3), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[23]), .B1(n3), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[24]), .B1(n3), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[25]), .B1(n3), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[26]), .B1(n3), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[27]), .B1(n3), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[28]), .B1(n3), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[29]), .B1(n3), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n4), .A2(i_data_bus[30]), .B1(n3), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n4), .A2(i_data_bus[31]), .B1(n3), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n4), .A2(n3), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_222 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_222 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_37 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_222 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_221 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_220 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_219 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_218 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_217 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  CKAN2D1BWP30P140LVT U2 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
  TIELBWP30P140LVT U3 ( .ZN(n_Logic0_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_223 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_223 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_223 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_224 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_224 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_224 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_225 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2D1BWP30P140LVT U36 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_225 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_225 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_226 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_226 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_226 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_227 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(n2), .A2(rst), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  BUFFD2BWP30P140LVT U7 ( .I(n3), .Z(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_227 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_227 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_228 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_228 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_228 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_38 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_228 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_227 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_226 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_225 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_224 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_223 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_229 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_229 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_229 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_230 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_230 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_230 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_231 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2D1BWP30P140LVT U36 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_231 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_231 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_232 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_232 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_232 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_233 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_233 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_233 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_234 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_234 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_234 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_39 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_234 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_233 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_232 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_231 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_230 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_229 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_235 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_235 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_235 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_236 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n1), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_236 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_236 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_237 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(N91) );
  CKAN2D1BWP30P140LVT U4 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  ND2D1BWP30P140LVT U36 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_237 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_237 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_238 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_238 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_238 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_239 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_239 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_239 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_240 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  BUFFD2BWP30P140LVT U4 ( .I(n4), .Z(n1) );
  NR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .ZN(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n1), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n1), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n1), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n1), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n1), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n1), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n1), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n1), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n1), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n1), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n1), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n1), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n1), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n1), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n1), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n1), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_240 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_240 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_40 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_240 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_239 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_238 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_237 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_236 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_235 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_241 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n33, n34, n35,
         n36;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  NR2OPTIBD6BWP30P140LVT U3 ( .A1(n34), .A2(rst), .ZN(n35) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n33) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n33), .A2(i_cmd[0]), .A3(rst), .ZN(n36) );
  ND3OPTPAD2BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(
        n34) );
  AO22D1BWP30P140LVT U7 ( .A1(n36), .A2(i_data_bus[0]), .B1(n35), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U8 ( .A1(n36), .A2(i_data_bus[1]), .B1(n35), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U9 ( .A1(n36), .A2(i_data_bus[2]), .B1(n35), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U10 ( .A1(n36), .A2(i_data_bus[3]), .B1(n35), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U11 ( .A1(n36), .A2(i_data_bus[4]), .B1(n35), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U12 ( .A1(n36), .A2(i_data_bus[5]), .B1(n35), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U13 ( .A1(n36), .A2(i_data_bus[6]), .B1(n35), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U14 ( .A1(n36), .A2(i_data_bus[7]), .B1(n35), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U15 ( .A1(n36), .A2(i_data_bus[8]), .B1(n35), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U16 ( .A1(n36), .A2(i_data_bus[9]), .B1(n35), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U17 ( .A1(n36), .A2(i_data_bus[10]), .B1(n35), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U18 ( .A1(n36), .A2(i_data_bus[11]), .B1(n35), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U19 ( .A1(n36), .A2(i_data_bus[12]), .B1(n35), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U20 ( .A1(n36), .A2(i_data_bus[13]), .B1(n35), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U21 ( .A1(n36), .A2(i_data_bus[14]), .B1(n35), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U22 ( .A1(n36), .A2(i_data_bus[15]), .B1(n35), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U23 ( .A1(n36), .A2(i_data_bus[16]), .B1(n35), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U24 ( .A1(n36), .A2(i_data_bus[17]), .B1(n35), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U25 ( .A1(n36), .A2(i_data_bus[18]), .B1(n35), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U26 ( .A1(n36), .A2(i_data_bus[19]), .B1(n35), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U27 ( .A1(n36), .A2(i_data_bus[20]), .B1(n35), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U28 ( .A1(n36), .A2(i_data_bus[21]), .B1(n35), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U29 ( .A1(n36), .A2(i_data_bus[22]), .B1(n35), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U30 ( .A1(n36), .A2(i_data_bus[23]), .B1(n35), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U31 ( .A1(n36), .A2(i_data_bus[24]), .B1(n35), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U32 ( .A1(n36), .A2(i_data_bus[25]), .B1(n35), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U33 ( .A1(n36), .A2(i_data_bus[26]), .B1(n35), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U34 ( .A1(n36), .A2(i_data_bus[27]), .B1(n35), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U35 ( .A1(n36), .A2(i_data_bus[28]), .B1(n35), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U36 ( .A1(n36), .A2(i_data_bus[29]), .B1(n35), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U37 ( .A1(n36), .A2(i_data_bus[30]), .B1(n35), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U38 ( .A1(n36), .A2(i_data_bus[31]), .B1(n35), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U39 ( .A1(n36), .A2(n35), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_241 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_241 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_242 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2D1BWP30P140LVT U3 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND2D1BWP30P140LVT U4 ( .A1(i_valid[1]), .A2(n2), .ZN(n3) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  INR2D1BWP30P140LVT U6 ( .A1(i_en), .B1(rst), .ZN(n2) );
  INR2D4BWP30P140LVT U7 ( .A1(i_cmd[0]), .B1(n3), .ZN(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_242 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_242 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_243 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D2BWP30P140LVT U3 ( .A1(i_cmd[0]), .A2(n3), .ZN(N91) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  IND2D1BWP30P140LVT U7 ( .A1(n2), .B1(n1), .ZN(n3) );
  INVD1BWP30P140LVT U8 ( .I(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U36 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U37 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U38 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_243 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_243 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_244 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2D1BWP30P140LVT U3 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND2D1BWP30P140LVT U4 ( .A1(i_valid[1]), .A2(n2), .ZN(n3) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  INR2D1BWP30P140LVT U6 ( .A1(i_en), .B1(rst), .ZN(n2) );
  INR2D4BWP30P140LVT U7 ( .A1(i_cmd[0]), .B1(n3), .ZN(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_244 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_244 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_245 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  INVD6BWP30P140LVT U3 ( .I(n4), .ZN(n5) );
  NR3D1P5BWP30P140LVT U4 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n6) );
  BUFFD4BWP30P140LVT U5 ( .I(n6), .Z(n1) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  ND3D1BWP30P140LVT U7 ( .A1(i_cmd[0]), .A2(i_valid[1]), .A3(i_en), .ZN(n3) );
  OR2D4BWP30P140LVT U8 ( .A1(n3), .A2(rst), .Z(n4) );
  AO22D1BWP30P140LVT U9 ( .A1(n1), .A2(i_data_bus[0]), .B1(n5), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n1), .A2(i_data_bus[1]), .B1(n5), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n1), .A2(i_data_bus[2]), .B1(n5), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n1), .A2(i_data_bus[3]), .B1(n5), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n1), .A2(i_data_bus[4]), .B1(n5), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n1), .A2(i_data_bus[5]), .B1(n5), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n1), .A2(i_data_bus[6]), .B1(n5), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n1), .A2(i_data_bus[7]), .B1(n5), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n1), .A2(i_data_bus[8]), .B1(n5), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n1), .A2(i_data_bus[9]), .B1(n5), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n1), .A2(i_data_bus[10]), .B1(n5), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n1), .A2(i_data_bus[11]), .B1(n5), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n1), .A2(i_data_bus[12]), .B1(n5), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n1), .A2(i_data_bus[13]), .B1(n5), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n1), .A2(i_data_bus[14]), .B1(n5), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n1), .A2(i_data_bus[15]), .B1(n5), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n1), .A2(i_data_bus[16]), .B1(n5), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n1), .A2(i_data_bus[17]), .B1(n5), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n1), .A2(i_data_bus[18]), .B1(n5), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n1), .A2(i_data_bus[19]), .B1(n5), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n1), .A2(i_data_bus[20]), .B1(n5), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n1), .A2(i_data_bus[21]), .B1(n5), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n1), .A2(i_data_bus[22]), .B1(n5), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n1), .A2(i_data_bus[23]), .B1(n5), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n1), .A2(i_data_bus[24]), .B1(n5), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n1), .A2(i_data_bus[25]), .B1(n5), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n1), .A2(i_data_bus[26]), .B1(n5), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n1), .A2(i_data_bus[27]), .B1(n5), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n1), .A2(i_data_bus[28]), .B1(n5), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n1), .A2(i_data_bus[29]), .B1(n5), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n1), .A2(i_data_bus[30]), .B1(n5), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n1), .A2(i_data_bus[31]), .B1(n5), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n1), .A2(n5), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_245 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_245 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_246 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  INVD6BWP30P140LVT U3 ( .I(n4), .ZN(n5) );
  OR3D2BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .Z(n2) );
  OR2D1BWP30P140LVT U5 ( .A1(n3), .A2(rst), .Z(n4) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  INVD8BWP30P140LVT U7 ( .I(n2), .ZN(n6) );
  ND3OPTPAD2BWP30P140LVT U8 ( .A1(i_cmd[0]), .A2(i_valid[1]), .A3(i_en), .ZN(
        n3) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n5), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n5), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n5), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n5), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n5), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n5), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n5), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n5), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n5), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n5), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n5), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n5), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n5), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n5), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n5), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n5), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n5), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n5), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n5), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n5), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n5), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n5), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n5), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n5), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n5), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n5), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n5), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n5), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n5), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n5), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n5), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n5), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n5), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_246 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_246 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_41 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_246 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_245 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_244 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_243 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_242 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_241 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_247 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2D1BWP30P140LVT U3 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  AN2D2BWP30P140LVT U4 ( .A1(i_cmd[0]), .A2(n1), .Z(n4) );
  CKAN2D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(n3), .Z(n1) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  INR2D1BWP30P140LVT U7 ( .A1(i_en), .B1(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_247 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_247 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_248 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n33, n34, n35,
         n36, n37;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  INVD6BWP30P140LVT U3 ( .I(n35), .ZN(n36) );
  OR2D2BWP30P140LVT U4 ( .A1(n34), .A2(rst), .Z(n35) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n33) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n33), .A2(i_cmd[0]), .A3(rst), .ZN(n37) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n34)
         );
  AO22D1BWP30P140LVT U8 ( .A1(n37), .A2(i_data_bus[0]), .B1(n36), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n37), .A2(i_data_bus[1]), .B1(n36), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n37), .A2(i_data_bus[2]), .B1(n36), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n37), .A2(i_data_bus[3]), .B1(n36), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n37), .A2(i_data_bus[4]), .B1(n36), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n37), .A2(i_data_bus[5]), .B1(n36), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n37), .A2(i_data_bus[6]), .B1(n36), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n37), .A2(i_data_bus[7]), .B1(n36), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n37), .A2(i_data_bus[8]), .B1(n36), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n37), .A2(i_data_bus[9]), .B1(n36), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n37), .A2(i_data_bus[10]), .B1(n36), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n37), .A2(i_data_bus[11]), .B1(n36), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n37), .A2(i_data_bus[12]), .B1(n36), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n37), .A2(i_data_bus[13]), .B1(n36), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n37), .A2(i_data_bus[14]), .B1(n36), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n37), .A2(i_data_bus[15]), .B1(n36), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n37), .A2(i_data_bus[16]), .B1(n36), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n37), .A2(i_data_bus[17]), .B1(n36), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n37), .A2(i_data_bus[18]), .B1(n36), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n37), .A2(i_data_bus[19]), .B1(n36), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n37), .A2(i_data_bus[20]), .B1(n36), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n37), .A2(i_data_bus[21]), .B1(n36), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n37), .A2(i_data_bus[22]), .B1(n36), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n37), .A2(i_data_bus[23]), .B1(n36), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n37), .A2(i_data_bus[24]), .B1(n36), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n37), .A2(i_data_bus[25]), .B1(n36), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n37), .A2(i_data_bus[26]), .B1(n36), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n37), .A2(i_data_bus[27]), .B1(n36), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n37), .A2(i_data_bus[28]), .B1(n36), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n37), .A2(i_data_bus[29]), .B1(n36), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n37), .A2(i_data_bus[30]), .B1(n36), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n37), .A2(i_data_bus[31]), .B1(n36), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n37), .A2(n36), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_248 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_248 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_249 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104,
         N105, N106, N107, N108, N109, N110, N111, N112, N113, N114, N115,
         N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(n4), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D2BWP30P140LVT U3 ( .A1(i_cmd[0]), .A2(n3), .ZN(n4) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n4), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n4), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n4), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n4), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n4), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n4), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n4), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n4), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n4), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n4), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n4), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n4), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n4), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n4), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n4), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n4), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n4), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n4), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n4), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n4), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n4), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n4), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n4), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n4), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n4), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n4), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n4), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n4), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n4), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n4), .A2(i_data_bus[31]), .Z(N123) );
  IND2D1BWP30P140LVT U37 ( .A1(n2), .B1(n1), .ZN(n3) );
  INVD1BWP30P140LVT U38 ( .I(rst), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_249 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_249 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_250 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  INVD6BWP30P140LVT U3 ( .I(n3), .ZN(n4) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  OR2D4BWP30P140LVT U7 ( .A1(n2), .A2(rst), .Z(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_250 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_250 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_251 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2OPTPAD4BWP30P140LVT U3 ( .A1(n3), .A2(rst), .ZN(n4) );
  NR3D0P7BWP30P140LVT U4 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D2BWP30P140LVT U5 ( .A1(i_cmd[0]), .A2(i_valid[1]), .A3(i_en), .ZN(n3) );
  BUFFD4BWP30P140LVT U6 ( .I(n5), .Z(n1) );
  ND2OPTIBD1BWP30P140LVT U7 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  AO22D1BWP30P140LVT U8 ( .A1(n1), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n1), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n1), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n1), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n1), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n1), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n1), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n1), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n1), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n1), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n1), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n1), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n1), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n1), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n1), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n1), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n1), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n1), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n1), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n1), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n1), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n1), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n1), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n1), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n1), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n1), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n1), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n1), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n1), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n1), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n1), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n1), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n1), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_251 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_251 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_252 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D0P7BWP30P140LVT U3 ( .A1(n3), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D2BWP30P140LVT U4 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n4) );
  NR2OPTPAD6BWP30P140LVT U5 ( .A1(n4), .A2(rst), .ZN(n2) );
  BUFFD4BWP30P140LVT U6 ( .I(n5), .Z(n1) );
  ND2OPTIBD1BWP30P140LVT U7 ( .A1(i_en), .A2(i_valid[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n1), .A2(i_data_bus[0]), .B1(n2), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n1), .A2(i_data_bus[1]), .B1(n2), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n1), .A2(i_data_bus[2]), .B1(n2), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n1), .A2(i_data_bus[3]), .B1(n2), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n1), .A2(i_data_bus[4]), .B1(n2), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n1), .A2(i_data_bus[5]), .B1(n2), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n1), .A2(i_data_bus[6]), .B1(n2), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n1), .A2(i_data_bus[7]), .B1(n2), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n1), .A2(i_data_bus[8]), .B1(n2), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n1), .A2(i_data_bus[9]), .B1(n2), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n1), .A2(i_data_bus[10]), .B1(n2), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n1), .A2(i_data_bus[11]), .B1(n2), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n1), .A2(i_data_bus[12]), .B1(n2), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n1), .A2(i_data_bus[13]), .B1(n2), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n1), .A2(i_data_bus[14]), .B1(n2), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n1), .A2(i_data_bus[15]), .B1(n2), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n1), .A2(i_data_bus[16]), .B1(n2), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n1), .A2(i_data_bus[17]), .B1(n2), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n1), .A2(i_data_bus[18]), .B1(n2), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n1), .A2(i_data_bus[19]), .B1(n2), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n1), .A2(i_data_bus[20]), .B1(n2), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n1), .A2(i_data_bus[21]), .B1(n2), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n1), .A2(i_data_bus[22]), .B1(n2), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n1), .A2(i_data_bus[23]), .B1(n2), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n1), .A2(i_data_bus[24]), .B1(n2), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n1), .A2(i_data_bus[25]), .B1(n2), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n1), .A2(i_data_bus[26]), .B1(n2), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n1), .A2(i_data_bus[27]), .B1(n2), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n1), .A2(i_data_bus[28]), .B1(n2), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n1), .A2(i_data_bus[29]), .B1(n2), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n1), .A2(i_data_bus[30]), .B1(n2), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n1), .A2(i_data_bus[31]), .B1(n2), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n1), .A2(n2), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_252 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_252 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_42 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_252 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_251 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_250 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_249 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_248 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_247 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_253 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  INVD8BWP30P140LVT U3 ( .I(n4), .ZN(n5) );
  NR3D1P5BWP30P140LVT U4 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n1) );
  ND3OPTPAD1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(
        n3) );
  ND2D1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3D1P5BWP30P140LVT U7 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n6) );
  OR2D4BWP30P140LVT U8 ( .A1(n3), .A2(rst), .Z(n4) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n5), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n1), .A2(i_data_bus[1]), .B1(n5), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n5), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n1), .A2(i_data_bus[3]), .B1(n5), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n5), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n1), .A2(i_data_bus[5]), .B1(n5), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n5), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n1), .A2(i_data_bus[7]), .B1(n5), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n5), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n1), .A2(i_data_bus[9]), .B1(n5), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n5), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n1), .A2(i_data_bus[11]), .B1(n5), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n5), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n1), .A2(i_data_bus[13]), .B1(n5), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n5), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n1), .A2(i_data_bus[15]), .B1(n5), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n5), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n1), .A2(i_data_bus[17]), .B1(n5), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n5), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n1), .A2(i_data_bus[19]), .B1(n5), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n5), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n1), .A2(i_data_bus[21]), .B1(n5), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n5), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n1), .A2(i_data_bus[23]), .B1(n5), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n5), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n1), .A2(i_data_bus[25]), .B1(n5), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n5), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n1), .A2(i_data_bus[27]), .B1(n5), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n5), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n1), .A2(i_data_bus[29]), .B1(n5), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n5), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n1), .A2(i_data_bus[31]), .B1(n5), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n5), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_253 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_253 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_254 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  INVD8BWP30P140LVT U3 ( .I(n4), .ZN(n5) );
  NR3D1P5BWP30P140LVT U4 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n1) );
  ND3OPTPAD1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(
        n3) );
  ND2D1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  NR3D1P5BWP30P140LVT U7 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n6) );
  OR2D4BWP30P140LVT U8 ( .A1(n3), .A2(rst), .Z(n4) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n5), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n1), .A2(i_data_bus[1]), .B1(n5), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n5), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n1), .A2(i_data_bus[3]), .B1(n5), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n5), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n1), .A2(i_data_bus[5]), .B1(n5), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n5), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n1), .A2(i_data_bus[7]), .B1(n5), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n5), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n1), .A2(i_data_bus[9]), .B1(n5), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n5), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n1), .A2(i_data_bus[11]), .B1(n5), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n5), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n1), .A2(i_data_bus[13]), .B1(n5), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n5), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n1), .A2(i_data_bus[15]), .B1(n5), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n5), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n1), .A2(i_data_bus[17]), .B1(n5), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n5), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n1), .A2(i_data_bus[19]), .B1(n5), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n5), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n1), .A2(i_data_bus[21]), .B1(n5), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n5), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n1), .A2(i_data_bus[23]), .B1(n5), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n5), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n1), .A2(i_data_bus[25]), .B1(n5), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n5), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n1), .A2(i_data_bus[27]), .B1(n5), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n5), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n1), .A2(i_data_bus[29]), .B1(n5), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n5), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n1), .A2(i_data_bus[31]), .B1(n5), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n5), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_254 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_254 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_255 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104,
         N105, N106, N107, N108, N109, N110, N111, N112, N113, N114, N115,
         N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4, n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(n5), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(i_cmd[0]), .A2(n4), .ZN(n5) );
  NR2D1BWP30P140LVT U4 ( .A1(i_cmd[0]), .A2(n4), .ZN(n1) );
  IND2D1BWP30P140LVT U5 ( .A1(n3), .B1(n2), .ZN(n4) );
  INVD1BWP30P140LVT U6 ( .I(rst), .ZN(n2) );
  ND2D1BWP30P140LVT U7 ( .A1(i_en), .A2(i_valid[0]), .ZN(n3) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(i_data_bus[31]), .Z(N123) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_255 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_255 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_256 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  INVD8BWP30P140LVT U3 ( .I(n3), .ZN(n4) );
  ND3D1BWP30P140LVT U4 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  OR2D4BWP30P140LVT U7 ( .A1(n2), .A2(rst), .Z(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_256 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_256 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_257 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  INVD6BWP30P140LVT U3 ( .I(n4), .ZN(n5) );
  OR3D2BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .Z(n2) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  INVD8BWP30P140LVT U7 ( .I(n2), .ZN(n6) );
  OR2D4BWP30P140LVT U8 ( .A1(n3), .A2(rst), .Z(n4) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n5), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n5), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n5), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n5), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n5), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n5), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n5), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n5), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n5), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n5), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n5), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n5), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n5), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n5), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n5), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n5), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n5), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n5), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n5), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n5), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n5), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n5), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n5), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n5), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n5), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n5), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n5), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n5), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n5), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n5), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n5), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n5), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n5), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_257 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_257 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_258 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  INVD6BWP30P140LVT U3 ( .I(n4), .ZN(n5) );
  OR3D2BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .Z(n2) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  INVD8BWP30P140LVT U7 ( .I(n2), .ZN(n6) );
  OR2D4BWP30P140LVT U8 ( .A1(n3), .A2(rst), .Z(n4) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n5), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n5), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n5), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n5), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n5), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n5), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n5), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n5), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n5), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n5), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n5), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n5), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n5), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n5), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n5), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n5), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n5), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n5), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n5), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n5), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n5), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n5), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n5), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n5), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n5), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n5), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n5), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n5), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n5), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n5), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n5), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n5), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n5), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_258 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_258 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_43 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_258 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_257 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_256 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_255 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_254 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_253 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_259 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  INVD1BWP30P140LVT U3 ( .I(rst), .ZN(n4) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n3) );
  AN2D4BWP30P140LVT U5 ( .A1(n5), .A2(n4), .Z(n1) );
  AN2D4BWP30P140LVT U6 ( .A1(n5), .A2(n4), .Z(n2) );
  NR3OPTPAD2BWP30P140LVT U7 ( .A1(n3), .A2(i_cmd[0]), .A3(rst), .ZN(n6) );
  AN3D2BWP30P140LVT U8 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .Z(n5) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n2), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n1), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n2), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n1), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n2), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n1), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n2), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n1), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n2), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n1), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n2), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n1), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n2), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n1), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n2), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n1), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n2), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n1), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n2), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n1), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n2), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n1), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n2), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n1), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n2), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n1), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n2), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n1), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n2), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n1), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n2), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n1), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n2), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_259 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_259 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_260 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n32, n33, n34,
         n35, n36;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  INVD6BWP30P140LVT U3 ( .I(n34), .ZN(n35) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n32) );
  AO22D1BWP30P140LVT U5 ( .A1(n36), .A2(i_data_bus[0]), .B1(n35), .B2(
        i_data_bus[32]), .Z(N92) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(i_cmd[0]), .A2(n32), .A3(rst), .ZN(n36) );
  ND3D1BWP30P140LVT U7 ( .A1(i_cmd[0]), .A2(i_en), .A3(i_valid[1]), .ZN(n33)
         );
  OR2D4BWP30P140LVT U8 ( .A1(n33), .A2(rst), .Z(n34) );
  AO22D1BWP30P140LVT U9 ( .A1(n36), .A2(i_data_bus[1]), .B1(n35), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n36), .A2(i_data_bus[2]), .B1(n35), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n36), .A2(i_data_bus[3]), .B1(n35), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n36), .A2(i_data_bus[4]), .B1(n35), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n36), .A2(i_data_bus[5]), .B1(n35), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n36), .A2(i_data_bus[6]), .B1(n35), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n36), .A2(i_data_bus[7]), .B1(n35), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n36), .A2(i_data_bus[8]), .B1(n35), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n36), .A2(i_data_bus[9]), .B1(n35), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n36), .A2(i_data_bus[10]), .B1(n35), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n36), .A2(i_data_bus[11]), .B1(n35), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n36), .A2(i_data_bus[12]), .B1(n35), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n36), .A2(i_data_bus[13]), .B1(n35), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n36), .A2(i_data_bus[14]), .B1(n35), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n36), .A2(i_data_bus[15]), .B1(n35), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n36), .A2(i_data_bus[16]), .B1(n35), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n36), .A2(i_data_bus[17]), .B1(n35), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n36), .A2(i_data_bus[18]), .B1(n35), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n36), .A2(i_data_bus[19]), .B1(n35), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n36), .A2(i_data_bus[20]), .B1(n35), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n36), .A2(i_data_bus[21]), .B1(n35), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n36), .A2(i_data_bus[22]), .B1(n35), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n36), .A2(i_data_bus[23]), .B1(n35), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n36), .A2(i_data_bus[24]), .B1(n35), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n36), .A2(i_data_bus[25]), .B1(n35), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n36), .A2(i_data_bus[26]), .B1(n35), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n36), .A2(i_data_bus[27]), .B1(n35), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n36), .A2(i_data_bus[28]), .B1(n35), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n36), .A2(i_data_bus[29]), .B1(n35), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n36), .A2(i_data_bus[30]), .B1(n35), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n36), .A2(i_data_bus[31]), .B1(n35), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n36), .A2(n35), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_260 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_260 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_261 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D2BWP30P140LVT U3 ( .A1(i_cmd[0]), .A2(n3), .ZN(N91) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U36 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  IND2D1BWP30P140LVT U37 ( .A1(n2), .B1(n1), .ZN(n3) );
  INVD1BWP30P140LVT U38 ( .I(rst), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_261 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_261 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_262 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n33, n34, n35,
         n36, n37;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  INVD6BWP30P140LVT U3 ( .I(n35), .ZN(n36) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n33) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n33), .A2(i_cmd[0]), .A3(rst), .ZN(n37) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n34)
         );
  OR2D4BWP30P140LVT U7 ( .A1(n34), .A2(rst), .Z(n35) );
  AO22D1BWP30P140LVT U8 ( .A1(n37), .A2(i_data_bus[0]), .B1(n36), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n37), .A2(i_data_bus[1]), .B1(n36), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n37), .A2(i_data_bus[2]), .B1(n36), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n37), .A2(i_data_bus[3]), .B1(n36), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n37), .A2(i_data_bus[4]), .B1(n36), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n37), .A2(i_data_bus[5]), .B1(n36), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n37), .A2(i_data_bus[6]), .B1(n36), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n37), .A2(i_data_bus[7]), .B1(n36), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n37), .A2(i_data_bus[8]), .B1(n36), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n37), .A2(i_data_bus[9]), .B1(n36), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n37), .A2(i_data_bus[10]), .B1(n36), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n37), .A2(i_data_bus[11]), .B1(n36), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n37), .A2(i_data_bus[12]), .B1(n36), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n37), .A2(i_data_bus[13]), .B1(n36), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n37), .A2(i_data_bus[14]), .B1(n36), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n37), .A2(i_data_bus[15]), .B1(n36), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n37), .A2(i_data_bus[16]), .B1(n36), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n37), .A2(i_data_bus[17]), .B1(n36), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n37), .A2(i_data_bus[18]), .B1(n36), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n37), .A2(i_data_bus[19]), .B1(n36), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n37), .A2(i_data_bus[20]), .B1(n36), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n37), .A2(i_data_bus[21]), .B1(n36), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n37), .A2(i_data_bus[22]), .B1(n36), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n37), .A2(i_data_bus[23]), .B1(n36), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n37), .A2(i_data_bus[24]), .B1(n36), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n37), .A2(i_data_bus[25]), .B1(n36), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n37), .A2(i_data_bus[26]), .B1(n36), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n37), .A2(i_data_bus[27]), .B1(n36), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n37), .A2(i_data_bus[28]), .B1(n36), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n37), .A2(i_data_bus[29]), .B1(n36), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n37), .A2(i_data_bus[30]), .B1(n36), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n37), .A2(i_data_bus[31]), .B1(n36), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n37), .A2(n36), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_262 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_262 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_263 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2OPTIBD1BWP30P140LVT U3 ( .A1(i_cmd[0]), .A2(n1), .ZN(n3) );
  INR2D1BWP30P140LVT U4 ( .A1(i_en), .B1(rst), .ZN(n2) );
  INVD2BWP30P140LVT U5 ( .I(n3), .ZN(n9) );
  AN3D2BWP30P140LVT U6 ( .A1(i_valid[0]), .A2(n6), .A3(n5), .Z(n10) );
  INVD1BWP30P140LVT U7 ( .I(n4), .ZN(n5) );
  ND2D1BWP30P140LVT U8 ( .A1(n8), .A2(n7), .ZN(N123) );
  ND2D1BWP30P140LVT U9 ( .A1(n10), .A2(i_data_bus[31]), .ZN(n7) );
  ND2D1BWP30P140LVT U10 ( .A1(n9), .A2(i_data_bus[63]), .ZN(n8) );
  CKAN2D1BWP30P140LVT U11 ( .A1(i_valid[1]), .A2(n2), .Z(n1) );
  INVD1BWP30P140LVT U12 ( .I(i_cmd[0]), .ZN(n6) );
  IND2D1BWP30P140LVT U13 ( .A1(rst), .B1(i_en), .ZN(n4) );
  AO22D1BWP30P140LVT U14 ( .A1(n10), .A2(i_data_bus[0]), .B1(n9), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U15 ( .A1(n10), .A2(i_data_bus[1]), .B1(n9), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U16 ( .A1(n10), .A2(i_data_bus[2]), .B1(n9), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U17 ( .A1(n10), .A2(i_data_bus[3]), .B1(n9), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U18 ( .A1(n10), .A2(i_data_bus[4]), .B1(n9), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U19 ( .A1(n10), .A2(i_data_bus[5]), .B1(n9), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U20 ( .A1(n10), .A2(i_data_bus[6]), .B1(n9), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U21 ( .A1(n10), .A2(i_data_bus[7]), .B1(n9), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U22 ( .A1(n10), .A2(i_data_bus[8]), .B1(n9), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U23 ( .A1(n10), .A2(i_data_bus[9]), .B1(n9), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U24 ( .A1(n10), .A2(i_data_bus[10]), .B1(n9), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U25 ( .A1(n10), .A2(i_data_bus[11]), .B1(n9), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U26 ( .A1(n10), .A2(i_data_bus[12]), .B1(n9), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U27 ( .A1(n10), .A2(i_data_bus[13]), .B1(n9), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U28 ( .A1(n10), .A2(i_data_bus[14]), .B1(n9), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U29 ( .A1(n10), .A2(i_data_bus[15]), .B1(n9), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U30 ( .A1(n10), .A2(i_data_bus[16]), .B1(n9), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U31 ( .A1(n10), .A2(i_data_bus[17]), .B1(n9), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U32 ( .A1(n10), .A2(i_data_bus[18]), .B1(n9), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U33 ( .A1(n10), .A2(i_data_bus[19]), .B1(n9), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U34 ( .A1(n10), .A2(i_data_bus[20]), .B1(n9), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U35 ( .A1(n10), .A2(i_data_bus[21]), .B1(n9), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U36 ( .A1(n10), .A2(i_data_bus[22]), .B1(n9), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U37 ( .A1(n10), .A2(i_data_bus[23]), .B1(n9), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U38 ( .A1(n10), .A2(i_data_bus[24]), .B1(n9), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U39 ( .A1(n10), .A2(i_data_bus[25]), .B1(n9), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U40 ( .A1(n10), .A2(i_data_bus[26]), .B1(n9), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U41 ( .A1(n10), .A2(i_data_bus[27]), .B1(n9), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U42 ( .A1(n10), .A2(i_data_bus[28]), .B1(n9), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U43 ( .A1(n10), .A2(i_data_bus[29]), .B1(n9), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U44 ( .A1(n10), .A2(i_data_bus[30]), .B1(n9), .B2(
        i_data_bus[62]), .Z(N122) );
  OR2D1BWP30P140LVT U45 ( .A1(n10), .A2(n9), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_263 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_263 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_264 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  INVD6BWP30P140LVT U3 ( .I(n2), .ZN(n7) );
  INVD1BWP30P140LVT U4 ( .I(i_valid[1]), .ZN(n5) );
  ND2OPTIBD1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  OR3D4BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .Z(n2) );
  INR2D1BWP30P140LVT U7 ( .A1(i_en), .B1(rst), .ZN(n3) );
  ND2OPTIBD2BWP30P140LVT U8 ( .A1(i_cmd[0]), .A2(n3), .ZN(n4) );
  NR2OPTPAD2BWP30P140LVT U9 ( .A1(n5), .A2(n4), .ZN(n6) );
  AO22D1BWP30P140LVT U10 ( .A1(n7), .A2(i_data_bus[0]), .B1(n6), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U11 ( .A1(n7), .A2(i_data_bus[1]), .B1(n6), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U12 ( .A1(n7), .A2(i_data_bus[2]), .B1(n6), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U13 ( .A1(n7), .A2(i_data_bus[3]), .B1(n6), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U14 ( .A1(n7), .A2(i_data_bus[4]), .B1(n6), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U15 ( .A1(n7), .A2(i_data_bus[5]), .B1(n6), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U16 ( .A1(n7), .A2(i_data_bus[6]), .B1(n6), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U17 ( .A1(n7), .A2(i_data_bus[7]), .B1(n6), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U18 ( .A1(n7), .A2(i_data_bus[8]), .B1(n6), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U19 ( .A1(n7), .A2(i_data_bus[9]), .B1(n6), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U20 ( .A1(n7), .A2(i_data_bus[10]), .B1(n6), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U21 ( .A1(n7), .A2(i_data_bus[11]), .B1(n6), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U22 ( .A1(n7), .A2(i_data_bus[12]), .B1(n6), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U23 ( .A1(n7), .A2(i_data_bus[13]), .B1(n6), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U24 ( .A1(n7), .A2(i_data_bus[14]), .B1(n6), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U25 ( .A1(n7), .A2(i_data_bus[15]), .B1(n6), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U26 ( .A1(n7), .A2(i_data_bus[16]), .B1(n6), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U27 ( .A1(n7), .A2(i_data_bus[17]), .B1(n6), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U28 ( .A1(n7), .A2(i_data_bus[18]), .B1(n6), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U29 ( .A1(n7), .A2(i_data_bus[19]), .B1(n6), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U30 ( .A1(n7), .A2(i_data_bus[20]), .B1(n6), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U31 ( .A1(n7), .A2(i_data_bus[21]), .B1(n6), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U32 ( .A1(n7), .A2(i_data_bus[22]), .B1(n6), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U33 ( .A1(n7), .A2(i_data_bus[23]), .B1(n6), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U34 ( .A1(n7), .A2(i_data_bus[24]), .B1(n6), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U35 ( .A1(n7), .A2(i_data_bus[25]), .B1(n6), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U36 ( .A1(n7), .A2(i_data_bus[26]), .B1(n6), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U37 ( .A1(n7), .A2(i_data_bus[27]), .B1(n6), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U38 ( .A1(n7), .A2(i_data_bus[28]), .B1(n6), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U39 ( .A1(n7), .A2(i_data_bus[29]), .B1(n6), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U40 ( .A1(n7), .A2(i_data_bus[30]), .B1(n6), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U41 ( .A1(n7), .A2(i_data_bus[31]), .B1(n6), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U42 ( .A1(n7), .A2(n6), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_264 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_264 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_44 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_264 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_263 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_262 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_261 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_260 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_259 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_265 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n32, n33, n34,
         n35, n36;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  INVD6BWP30P140LVT U3 ( .I(n34), .ZN(n35) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n32) );
  AO22D1BWP30P140LVT U5 ( .A1(n36), .A2(i_data_bus[0]), .B1(n35), .B2(
        i_data_bus[32]), .Z(N92) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(i_cmd[0]), .A2(n32), .A3(rst), .ZN(n36) );
  ND3D1BWP30P140LVT U7 ( .A1(i_cmd[0]), .A2(i_en), .A3(i_valid[1]), .ZN(n33)
         );
  OR2D4BWP30P140LVT U8 ( .A1(n33), .A2(rst), .Z(n34) );
  AO22D1BWP30P140LVT U9 ( .A1(n36), .A2(i_data_bus[1]), .B1(n35), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n36), .A2(i_data_bus[2]), .B1(n35), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n36), .A2(i_data_bus[3]), .B1(n35), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n36), .A2(i_data_bus[4]), .B1(n35), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n36), .A2(i_data_bus[5]), .B1(n35), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n36), .A2(i_data_bus[6]), .B1(n35), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n36), .A2(i_data_bus[7]), .B1(n35), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n36), .A2(i_data_bus[8]), .B1(n35), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n36), .A2(i_data_bus[9]), .B1(n35), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n36), .A2(i_data_bus[10]), .B1(n35), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n36), .A2(i_data_bus[11]), .B1(n35), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n36), .A2(i_data_bus[12]), .B1(n35), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n36), .A2(i_data_bus[13]), .B1(n35), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n36), .A2(i_data_bus[14]), .B1(n35), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n36), .A2(i_data_bus[15]), .B1(n35), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n36), .A2(i_data_bus[16]), .B1(n35), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n36), .A2(i_data_bus[17]), .B1(n35), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n36), .A2(i_data_bus[18]), .B1(n35), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n36), .A2(i_data_bus[19]), .B1(n35), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n36), .A2(i_data_bus[20]), .B1(n35), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n36), .A2(i_data_bus[21]), .B1(n35), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n36), .A2(i_data_bus[22]), .B1(n35), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n36), .A2(i_data_bus[23]), .B1(n35), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n36), .A2(i_data_bus[24]), .B1(n35), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n36), .A2(i_data_bus[25]), .B1(n35), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n36), .A2(i_data_bus[26]), .B1(n35), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n36), .A2(i_data_bus[27]), .B1(n35), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n36), .A2(i_data_bus[28]), .B1(n35), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n36), .A2(i_data_bus[29]), .B1(n35), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n36), .A2(i_data_bus[30]), .B1(n35), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n36), .A2(i_data_bus[31]), .B1(n35), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n36), .A2(n35), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_265 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_265 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_266 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2D1BWP30P140LVT U3 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  ND2D1BWP30P140LVT U4 ( .A1(i_valid[1]), .A2(n2), .ZN(n3) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  INR2D1BWP30P140LVT U6 ( .A1(i_en), .B1(rst), .ZN(n2) );
  INR2D4BWP30P140LVT U7 ( .A1(i_cmd[0]), .B1(n3), .ZN(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_266 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_266 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_267 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D2BWP30P140LVT U3 ( .A1(i_cmd[0]), .A2(n3), .ZN(N91) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U36 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  IND2D1BWP30P140LVT U37 ( .A1(n2), .B1(n1), .ZN(n3) );
  INVD1BWP30P140LVT U38 ( .I(rst), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_267 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_267 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_268 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n33, n34, n35,
         n36, n37;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  INVD6BWP30P140LVT U3 ( .I(n35), .ZN(n36) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n33) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n33), .A2(i_cmd[0]), .A3(rst), .ZN(n37) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n34)
         );
  OR2D4BWP30P140LVT U7 ( .A1(n34), .A2(rst), .Z(n35) );
  AO22D1BWP30P140LVT U8 ( .A1(n37), .A2(i_data_bus[0]), .B1(n36), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n37), .A2(i_data_bus[1]), .B1(n36), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n37), .A2(i_data_bus[2]), .B1(n36), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n37), .A2(i_data_bus[3]), .B1(n36), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n37), .A2(i_data_bus[4]), .B1(n36), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n37), .A2(i_data_bus[5]), .B1(n36), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n37), .A2(i_data_bus[6]), .B1(n36), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n37), .A2(i_data_bus[7]), .B1(n36), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n37), .A2(i_data_bus[8]), .B1(n36), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n37), .A2(i_data_bus[9]), .B1(n36), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n37), .A2(i_data_bus[10]), .B1(n36), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n37), .A2(i_data_bus[11]), .B1(n36), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n37), .A2(i_data_bus[12]), .B1(n36), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n37), .A2(i_data_bus[13]), .B1(n36), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n37), .A2(i_data_bus[14]), .B1(n36), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n37), .A2(i_data_bus[15]), .B1(n36), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n37), .A2(i_data_bus[16]), .B1(n36), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n37), .A2(i_data_bus[17]), .B1(n36), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n37), .A2(i_data_bus[18]), .B1(n36), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n37), .A2(i_data_bus[19]), .B1(n36), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n37), .A2(i_data_bus[20]), .B1(n36), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n37), .A2(i_data_bus[21]), .B1(n36), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n37), .A2(i_data_bus[22]), .B1(n36), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n37), .A2(i_data_bus[23]), .B1(n36), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n37), .A2(i_data_bus[24]), .B1(n36), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n37), .A2(i_data_bus[25]), .B1(n36), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n37), .A2(i_data_bus[26]), .B1(n36), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n37), .A2(i_data_bus[27]), .B1(n36), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n37), .A2(i_data_bus[28]), .B1(n36), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n37), .A2(i_data_bus[29]), .B1(n36), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n37), .A2(i_data_bus[30]), .B1(n36), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n37), .A2(i_data_bus[31]), .B1(n36), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n37), .A2(n36), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_268 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_268 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_269 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  INVD6BWP30P140LVT U3 ( .I(n4), .ZN(n5) );
  OR3D2BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .Z(n2) );
  ND3D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  INVD8BWP30P140LVT U7 ( .I(n2), .ZN(n6) );
  OR2D4BWP30P140LVT U8 ( .A1(n3), .A2(rst), .Z(n4) );
  AO22D1BWP30P140LVT U9 ( .A1(n6), .A2(i_data_bus[0]), .B1(n5), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U10 ( .A1(n6), .A2(i_data_bus[1]), .B1(n5), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U11 ( .A1(n6), .A2(i_data_bus[2]), .B1(n5), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U12 ( .A1(n6), .A2(i_data_bus[3]), .B1(n5), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U13 ( .A1(n6), .A2(i_data_bus[4]), .B1(n5), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U14 ( .A1(n6), .A2(i_data_bus[5]), .B1(n5), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U15 ( .A1(n6), .A2(i_data_bus[6]), .B1(n5), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U16 ( .A1(n6), .A2(i_data_bus[7]), .B1(n5), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U17 ( .A1(n6), .A2(i_data_bus[8]), .B1(n5), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U18 ( .A1(n6), .A2(i_data_bus[9]), .B1(n5), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U19 ( .A1(n6), .A2(i_data_bus[10]), .B1(n5), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U20 ( .A1(n6), .A2(i_data_bus[11]), .B1(n5), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U21 ( .A1(n6), .A2(i_data_bus[12]), .B1(n5), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U22 ( .A1(n6), .A2(i_data_bus[13]), .B1(n5), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U23 ( .A1(n6), .A2(i_data_bus[14]), .B1(n5), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U24 ( .A1(n6), .A2(i_data_bus[15]), .B1(n5), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U25 ( .A1(n6), .A2(i_data_bus[16]), .B1(n5), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U26 ( .A1(n6), .A2(i_data_bus[17]), .B1(n5), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U27 ( .A1(n6), .A2(i_data_bus[18]), .B1(n5), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U28 ( .A1(n6), .A2(i_data_bus[19]), .B1(n5), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U29 ( .A1(n6), .A2(i_data_bus[20]), .B1(n5), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U30 ( .A1(n6), .A2(i_data_bus[21]), .B1(n5), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U31 ( .A1(n6), .A2(i_data_bus[22]), .B1(n5), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U32 ( .A1(n6), .A2(i_data_bus[23]), .B1(n5), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U33 ( .A1(n6), .A2(i_data_bus[24]), .B1(n5), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U34 ( .A1(n6), .A2(i_data_bus[25]), .B1(n5), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U35 ( .A1(n6), .A2(i_data_bus[26]), .B1(n5), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U36 ( .A1(n6), .A2(i_data_bus[27]), .B1(n5), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U37 ( .A1(n6), .A2(i_data_bus[28]), .B1(n5), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U38 ( .A1(n6), .A2(i_data_bus[29]), .B1(n5), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U39 ( .A1(n6), .A2(i_data_bus[30]), .B1(n5), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U40 ( .A1(n6), .A2(i_data_bus[31]), .B1(n5), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U41 ( .A1(n6), .A2(n5), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_269 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_269 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_270 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  INVD6BWP30P140LVT U3 ( .I(n2), .ZN(n7) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  OR3D4BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .Z(n2) );
  INVD1BWP30P140LVT U6 ( .I(i_valid[1]), .ZN(n5) );
  INR2D1BWP30P140LVT U7 ( .A1(i_en), .B1(rst), .ZN(n3) );
  ND2OPTIBD2BWP30P140LVT U8 ( .A1(i_cmd[0]), .A2(n3), .ZN(n4) );
  NR2OPTPAD2BWP30P140LVT U9 ( .A1(n5), .A2(n4), .ZN(n6) );
  AO22D1BWP30P140LVT U10 ( .A1(n7), .A2(i_data_bus[0]), .B1(n6), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U11 ( .A1(n7), .A2(i_data_bus[1]), .B1(n6), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U12 ( .A1(n7), .A2(i_data_bus[2]), .B1(n6), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U13 ( .A1(n7), .A2(i_data_bus[3]), .B1(n6), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U14 ( .A1(n7), .A2(i_data_bus[4]), .B1(n6), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U15 ( .A1(n7), .A2(i_data_bus[5]), .B1(n6), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U16 ( .A1(n7), .A2(i_data_bus[6]), .B1(n6), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U17 ( .A1(n7), .A2(i_data_bus[7]), .B1(n6), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U18 ( .A1(n7), .A2(i_data_bus[8]), .B1(n6), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U19 ( .A1(n7), .A2(i_data_bus[9]), .B1(n6), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U20 ( .A1(n7), .A2(i_data_bus[10]), .B1(n6), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U21 ( .A1(n7), .A2(i_data_bus[11]), .B1(n6), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U22 ( .A1(n7), .A2(i_data_bus[12]), .B1(n6), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U23 ( .A1(n7), .A2(i_data_bus[13]), .B1(n6), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U24 ( .A1(n7), .A2(i_data_bus[14]), .B1(n6), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U25 ( .A1(n7), .A2(i_data_bus[15]), .B1(n6), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U26 ( .A1(n7), .A2(i_data_bus[16]), .B1(n6), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U27 ( .A1(n7), .A2(i_data_bus[17]), .B1(n6), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U28 ( .A1(n7), .A2(i_data_bus[18]), .B1(n6), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U29 ( .A1(n7), .A2(i_data_bus[19]), .B1(n6), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U30 ( .A1(n7), .A2(i_data_bus[20]), .B1(n6), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U31 ( .A1(n7), .A2(i_data_bus[21]), .B1(n6), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U32 ( .A1(n7), .A2(i_data_bus[22]), .B1(n6), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U33 ( .A1(n7), .A2(i_data_bus[23]), .B1(n6), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U34 ( .A1(n7), .A2(i_data_bus[24]), .B1(n6), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U35 ( .A1(n7), .A2(i_data_bus[25]), .B1(n6), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U36 ( .A1(n7), .A2(i_data_bus[26]), .B1(n6), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U37 ( .A1(n7), .A2(i_data_bus[27]), .B1(n6), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U38 ( .A1(n7), .A2(i_data_bus[28]), .B1(n6), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U39 ( .A1(n7), .A2(i_data_bus[29]), .B1(n6), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U40 ( .A1(n7), .A2(i_data_bus[30]), .B1(n6), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U41 ( .A1(n7), .A2(i_data_bus[31]), .B1(n6), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U42 ( .A1(n7), .A2(n6), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_270 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_270 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_45 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_270 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_269 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_268 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_267 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_266 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_265 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[0]), .A2(i_cmd[1]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_271 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  INVD6BWP30P140LVT U3 ( .I(n3), .ZN(n4) );
  ND3D1BWP30P140LVT U4 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  OR2D4BWP30P140LVT U7 ( .A1(n2), .A2(rst), .Z(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_271 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_271 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_272 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n33, n34, n35,
         n36, n37;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  INVD6BWP30P140LVT U3 ( .I(n35), .ZN(n36) );
  OR2D2BWP30P140LVT U4 ( .A1(n34), .A2(rst), .Z(n35) );
  ND2D1BWP30P140LVT U5 ( .A1(i_en), .A2(i_valid[0]), .ZN(n33) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n33), .A2(i_cmd[0]), .A3(rst), .ZN(n37) );
  ND3D1BWP30P140LVT U7 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n34)
         );
  AO22D1BWP30P140LVT U8 ( .A1(n37), .A2(i_data_bus[0]), .B1(n36), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n37), .A2(i_data_bus[1]), .B1(n36), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n37), .A2(i_data_bus[2]), .B1(n36), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n37), .A2(i_data_bus[3]), .B1(n36), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n37), .A2(i_data_bus[4]), .B1(n36), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n37), .A2(i_data_bus[5]), .B1(n36), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n37), .A2(i_data_bus[6]), .B1(n36), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n37), .A2(i_data_bus[7]), .B1(n36), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n37), .A2(i_data_bus[8]), .B1(n36), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n37), .A2(i_data_bus[9]), .B1(n36), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n37), .A2(i_data_bus[10]), .B1(n36), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n37), .A2(i_data_bus[11]), .B1(n36), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n37), .A2(i_data_bus[12]), .B1(n36), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n37), .A2(i_data_bus[13]), .B1(n36), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n37), .A2(i_data_bus[14]), .B1(n36), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n37), .A2(i_data_bus[15]), .B1(n36), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n37), .A2(i_data_bus[16]), .B1(n36), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n37), .A2(i_data_bus[17]), .B1(n36), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n37), .A2(i_data_bus[18]), .B1(n36), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n37), .A2(i_data_bus[19]), .B1(n36), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n37), .A2(i_data_bus[20]), .B1(n36), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n37), .A2(i_data_bus[21]), .B1(n36), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n37), .A2(i_data_bus[22]), .B1(n36), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n37), .A2(i_data_bus[23]), .B1(n36), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n37), .A2(i_data_bus[24]), .B1(n36), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n37), .A2(i_data_bus[25]), .B1(n36), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n37), .A2(i_data_bus[26]), .B1(n36), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n37), .A2(i_data_bus[27]), .B1(n36), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n37), .A2(i_data_bus[28]), .B1(n36), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n37), .A2(i_data_bus[29]), .B1(n36), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n37), .A2(i_data_bus[30]), .B1(n36), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n37), .A2(i_data_bus[31]), .B1(n36), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n37), .A2(n36), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_272 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_272 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_273 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D2BWP30P140LVT U3 ( .A1(i_cmd[0]), .A2(n3), .ZN(N91) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U36 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  IND2D1BWP30P140LVT U37 ( .A1(n2), .B1(n1), .ZN(n3) );
  INVD1BWP30P140LVT U38 ( .I(rst), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_273 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_273 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_274 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  INVD6BWP30P140LVT U3 ( .I(n3), .ZN(n4) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  NR3OPTPAD2BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D1BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n2) );
  OR2D4BWP30P140LVT U7 ( .A1(n2), .A2(rst), .Z(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_274 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_274 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_275 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D8BWP30P140LVT U3 ( .A1(n4), .A2(rst), .ZN(n2) );
  BUFFD4BWP30P140LVT U4 ( .I(n5), .Z(n1) );
  NR3D0P7BWP30P140LVT U5 ( .A1(n3), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  ND3D3BWP30P140LVT U6 ( .A1(i_valid[1]), .A2(i_en), .A3(i_cmd[0]), .ZN(n4) );
  ND2D1BWP30P140LVT U7 ( .A1(i_en), .A2(i_valid[0]), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n1), .A2(i_data_bus[0]), .B1(n2), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n1), .A2(i_data_bus[1]), .B1(n2), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n1), .A2(i_data_bus[2]), .B1(n2), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n1), .A2(i_data_bus[3]), .B1(n2), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n1), .A2(i_data_bus[4]), .B1(n2), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n1), .A2(i_data_bus[5]), .B1(n2), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n1), .A2(i_data_bus[6]), .B1(n2), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n1), .A2(i_data_bus[7]), .B1(n2), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n1), .A2(i_data_bus[8]), .B1(n2), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n1), .A2(i_data_bus[9]), .B1(n2), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n1), .A2(i_data_bus[10]), .B1(n2), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n1), .A2(i_data_bus[11]), .B1(n2), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n1), .A2(i_data_bus[12]), .B1(n2), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n1), .A2(i_data_bus[13]), .B1(n2), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n1), .A2(i_data_bus[14]), .B1(n2), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n1), .A2(i_data_bus[15]), .B1(n2), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n1), .A2(i_data_bus[16]), .B1(n2), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n1), .A2(i_data_bus[17]), .B1(n2), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n1), .A2(i_data_bus[18]), .B1(n2), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n1), .A2(i_data_bus[19]), .B1(n2), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n1), .A2(i_data_bus[20]), .B1(n2), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n1), .A2(i_data_bus[21]), .B1(n2), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n1), .A2(i_data_bus[22]), .B1(n2), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n1), .A2(i_data_bus[23]), .B1(n2), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n1), .A2(i_data_bus[24]), .B1(n2), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n1), .A2(i_data_bus[25]), .B1(n2), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n1), .A2(i_data_bus[26]), .B1(n2), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n1), .A2(i_data_bus[27]), .B1(n2), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n1), .A2(i_data_bus[28]), .B1(n2), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n1), .A2(i_data_bus[29]), .B1(n2), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n1), .A2(i_data_bus[30]), .B1(n2), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n1), .A2(i_data_bus[31]), .B1(n2), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n1), .A2(n2), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_275 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_275 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_276 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U3 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n43) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_valid[0]), .A2(i_en), .ZN(n2) );
  INVD1BWP30P140LVT U5 ( .I(n43), .ZN(n1) );
  ND2OPTIBD1BWP30P140LVT U6 ( .A1(i_cmd[0]), .A2(n3), .ZN(n4) );
  INVD1BWP30P140LVT U7 ( .I(i_data_bus[0]), .ZN(n5) );
  INVD1BWP30P140LVT U8 ( .I(i_data_bus[1]), .ZN(n6) );
  INVD1BWP30P140LVT U9 ( .I(i_data_bus[2]), .ZN(n7) );
  INVD1BWP30P140LVT U10 ( .I(i_data_bus[3]), .ZN(n8) );
  INVD1BWP30P140LVT U11 ( .I(i_data_bus[4]), .ZN(n10) );
  INVD1BWP30P140LVT U12 ( .I(i_data_bus[5]), .ZN(n11) );
  INVD1BWP30P140LVT U13 ( .I(i_data_bus[6]), .ZN(n12) );
  INVD1BWP30P140LVT U14 ( .I(i_data_bus[7]), .ZN(n14) );
  INVD1BWP30P140LVT U15 ( .I(i_data_bus[8]), .ZN(n16) );
  INVD1BWP30P140LVT U16 ( .I(i_data_bus[9]), .ZN(n18) );
  INVD1BWP30P140LVT U17 ( .I(i_data_bus[10]), .ZN(n20) );
  INVD1BWP30P140LVT U18 ( .I(i_data_bus[11]), .ZN(n21) );
  INVD1BWP30P140LVT U19 ( .I(i_data_bus[12]), .ZN(n22) );
  INVD1BWP30P140LVT U20 ( .I(i_data_bus[13]), .ZN(n23) );
  INVD1BWP30P140LVT U21 ( .I(i_data_bus[14]), .ZN(n24) );
  INVD1BWP30P140LVT U22 ( .I(i_data_bus[15]), .ZN(n25) );
  INVD1BWP30P140LVT U23 ( .I(i_data_bus[16]), .ZN(n26) );
  INVD1BWP30P140LVT U24 ( .I(i_data_bus[17]), .ZN(n27) );
  INVD1BWP30P140LVT U25 ( .I(i_data_bus[18]), .ZN(n28) );
  INVD1BWP30P140LVT U26 ( .I(i_data_bus[19]), .ZN(n29) );
  INVD1BWP30P140LVT U27 ( .I(i_data_bus[20]), .ZN(n30) );
  INVD1BWP30P140LVT U28 ( .I(i_data_bus[21]), .ZN(n31) );
  INVD1BWP30P140LVT U29 ( .I(i_data_bus[22]), .ZN(n32) );
  INVD1BWP30P140LVT U30 ( .I(i_data_bus[23]), .ZN(n33) );
  INVD1BWP30P140LVT U31 ( .I(i_data_bus[24]), .ZN(n34) );
  INVD1BWP30P140LVT U32 ( .I(i_data_bus[25]), .ZN(n35) );
  INVD1BWP30P140LVT U33 ( .I(i_data_bus[26]), .ZN(n36) );
  INVD1BWP30P140LVT U34 ( .I(i_data_bus[27]), .ZN(n37) );
  INVD1BWP30P140LVT U35 ( .I(i_data_bus[28]), .ZN(n38) );
  INVD1BWP30P140LVT U36 ( .I(i_data_bus[29]), .ZN(n39) );
  INVD1BWP30P140LVT U37 ( .I(i_data_bus[30]), .ZN(n40) );
  INVD1BWP30P140LVT U38 ( .I(i_data_bus[31]), .ZN(n41) );
  INR2D1BWP30P140LVT U39 ( .A1(i_en), .B1(rst), .ZN(n3) );
  INR2D2BWP30P140LVT U40 ( .A1(i_valid[1]), .B1(n4), .ZN(n42) );
  MOAI22D1BWP30P140LVT U41 ( .A1(n13), .A2(n5), .B1(n42), .B2(i_data_bus[32]), 
        .ZN(N92) );
  MOAI22D1BWP30P140LVT U42 ( .A1(n9), .A2(n6), .B1(n42), .B2(i_data_bus[33]), 
        .ZN(N93) );
  MOAI22D1BWP30P140LVT U43 ( .A1(n17), .A2(n7), .B1(n42), .B2(i_data_bus[34]), 
        .ZN(N94) );
  INVD1BWP30P140LVT U44 ( .I(n43), .ZN(n9) );
  MOAI22D1BWP30P140LVT U45 ( .A1(n9), .A2(n8), .B1(n42), .B2(i_data_bus[35]), 
        .ZN(N95) );
  MOAI22D1BWP30P140LVT U46 ( .A1(n9), .A2(n10), .B1(n42), .B2(i_data_bus[36]), 
        .ZN(N96) );
  MOAI22D1BWP30P140LVT U47 ( .A1(n13), .A2(n11), .B1(n42), .B2(i_data_bus[37]), 
        .ZN(N97) );
  INVD1BWP30P140LVT U48 ( .I(n43), .ZN(n13) );
  MOAI22D1BWP30P140LVT U49 ( .A1(n13), .A2(n12), .B1(n42), .B2(i_data_bus[38]), 
        .ZN(N98) );
  INVD1BWP30P140LVT U50 ( .I(n43), .ZN(n15) );
  MOAI22D1BWP30P140LVT U51 ( .A1(n15), .A2(n14), .B1(n42), .B2(i_data_bus[39]), 
        .ZN(N99) );
  INVD1BWP30P140LVT U52 ( .I(n43), .ZN(n17) );
  MOAI22D1BWP30P140LVT U53 ( .A1(n17), .A2(n16), .B1(n42), .B2(i_data_bus[40]), 
        .ZN(N100) );
  INVD1BWP30P140LVT U54 ( .I(n43), .ZN(n19) );
  MOAI22D1BWP30P140LVT U55 ( .A1(n19), .A2(n18), .B1(n42), .B2(i_data_bus[41]), 
        .ZN(N101) );
  MOAI22D1BWP30P140LVT U56 ( .A1(n1), .A2(n20), .B1(n42), .B2(i_data_bus[42]), 
        .ZN(N102) );
  MOAI22D1BWP30P140LVT U57 ( .A1(n1), .A2(n21), .B1(n42), .B2(i_data_bus[43]), 
        .ZN(N103) );
  MOAI22D1BWP30P140LVT U58 ( .A1(n17), .A2(n22), .B1(n42), .B2(i_data_bus[44]), 
        .ZN(N104) );
  MOAI22D1BWP30P140LVT U59 ( .A1(n9), .A2(n23), .B1(n42), .B2(i_data_bus[45]), 
        .ZN(N105) );
  MOAI22D1BWP30P140LVT U60 ( .A1(n9), .A2(n24), .B1(n42), .B2(i_data_bus[46]), 
        .ZN(N106) );
  MOAI22D1BWP30P140LVT U61 ( .A1(n1), .A2(n25), .B1(n42), .B2(i_data_bus[47]), 
        .ZN(N107) );
  MOAI22D1BWP30P140LVT U62 ( .A1(n13), .A2(n26), .B1(n42), .B2(i_data_bus[48]), 
        .ZN(N108) );
  MOAI22D1BWP30P140LVT U63 ( .A1(n15), .A2(n27), .B1(n42), .B2(i_data_bus[49]), 
        .ZN(N109) );
  MOAI22D1BWP30P140LVT U64 ( .A1(n17), .A2(n28), .B1(n42), .B2(i_data_bus[50]), 
        .ZN(N110) );
  MOAI22D1BWP30P140LVT U65 ( .A1(n19), .A2(n29), .B1(n42), .B2(i_data_bus[51]), 
        .ZN(N111) );
  MOAI22D1BWP30P140LVT U66 ( .A1(n15), .A2(n30), .B1(n42), .B2(i_data_bus[52]), 
        .ZN(N112) );
  MOAI22D1BWP30P140LVT U67 ( .A1(n19), .A2(n31), .B1(n42), .B2(i_data_bus[53]), 
        .ZN(N113) );
  MOAI22D1BWP30P140LVT U68 ( .A1(n1), .A2(n32), .B1(n42), .B2(i_data_bus[54]), 
        .ZN(N114) );
  MOAI22D1BWP30P140LVT U69 ( .A1(n13), .A2(n33), .B1(n42), .B2(i_data_bus[55]), 
        .ZN(N115) );
  MOAI22D1BWP30P140LVT U70 ( .A1(n19), .A2(n34), .B1(n42), .B2(i_data_bus[56]), 
        .ZN(N116) );
  MOAI22D1BWP30P140LVT U71 ( .A1(n15), .A2(n35), .B1(n42), .B2(i_data_bus[57]), 
        .ZN(N117) );
  MOAI22D1BWP30P140LVT U72 ( .A1(n1), .A2(n36), .B1(n42), .B2(i_data_bus[58]), 
        .ZN(N118) );
  MOAI22D1BWP30P140LVT U73 ( .A1(n1), .A2(n37), .B1(n42), .B2(i_data_bus[59]), 
        .ZN(N119) );
  MOAI22D1BWP30P140LVT U74 ( .A1(n19), .A2(n38), .B1(n42), .B2(i_data_bus[60]), 
        .ZN(N120) );
  MOAI22D1BWP30P140LVT U75 ( .A1(n17), .A2(n39), .B1(n42), .B2(i_data_bus[61]), 
        .ZN(N121) );
  MOAI22D1BWP30P140LVT U76 ( .A1(n15), .A2(n40), .B1(n42), .B2(i_data_bus[62]), 
        .ZN(N122) );
  MOAI22D1BWP30P140LVT U77 ( .A1(n13), .A2(n41), .B1(n42), .B2(i_data_bus[63]), 
        .ZN(N123) );
  OR2D1BWP30P140LVT U78 ( .A1(n43), .A2(n42), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_276 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_276 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_46 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_276 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_275 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_274 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_273 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_272 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_271 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_277 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2D1BWP30P140LVT U3 ( .A1(i_en), .A2(i_valid[0]), .ZN(n3) );
  AN2D2BWP30P140LVT U4 ( .A1(i_cmd[0]), .A2(n1), .Z(n5) );
  CKAN2D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(n4), .Z(n1) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n3), .A2(i_cmd[0]), .A3(rst), .ZN(n2) );
  INR2D1BWP30P140LVT U7 ( .A1(i_en), .B1(rst), .ZN(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n2), .A2(i_data_bus[0]), .B1(n5), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n2), .A2(i_data_bus[1]), .B1(n5), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n2), .A2(i_data_bus[2]), .B1(n5), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n2), .A2(i_data_bus[3]), .B1(n5), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n2), .A2(i_data_bus[4]), .B1(n5), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n2), .A2(i_data_bus[5]), .B1(n5), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n2), .A2(i_data_bus[6]), .B1(n5), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n2), .A2(i_data_bus[7]), .B1(n5), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n2), .A2(i_data_bus[8]), .B1(n5), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n2), .A2(i_data_bus[9]), .B1(n5), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n2), .A2(i_data_bus[10]), .B1(n5), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n2), .A2(i_data_bus[11]), .B1(n5), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n2), .A2(i_data_bus[12]), .B1(n5), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n2), .A2(i_data_bus[13]), .B1(n5), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n2), .A2(i_data_bus[14]), .B1(n5), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n2), .A2(i_data_bus[15]), .B1(n5), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n2), .A2(i_data_bus[16]), .B1(n5), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n2), .A2(i_data_bus[17]), .B1(n5), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n2), .A2(i_data_bus[18]), .B1(n5), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n2), .A2(i_data_bus[19]), .B1(n5), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n2), .A2(i_data_bus[20]), .B1(n5), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n2), .A2(i_data_bus[21]), .B1(n5), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n2), .A2(i_data_bus[22]), .B1(n5), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n2), .A2(i_data_bus[23]), .B1(n5), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n2), .A2(i_data_bus[24]), .B1(n5), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n2), .A2(i_data_bus[25]), .B1(n5), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n2), .A2(i_data_bus[26]), .B1(n5), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n2), .A2(i_data_bus[27]), .B1(n5), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n2), .A2(i_data_bus[28]), .B1(n5), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n2), .A2(i_data_bus[29]), .B1(n5), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n2), .A2(i_data_bus[30]), .B1(n5), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n2), .A2(i_data_bus[31]), .B1(n5), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n2), .A2(n5), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_277 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_277 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_278 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2D1BWP30P140LVT U3 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  AN2D2BWP30P140LVT U4 ( .A1(i_cmd[0]), .A2(n1), .Z(n4) );
  CKAN2D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(n3), .Z(n1) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n2), .A2(i_cmd[0]), .A3(rst), .ZN(n5) );
  INR2D1BWP30P140LVT U7 ( .A1(i_en), .B1(rst), .ZN(n3) );
  AO22D1BWP30P140LVT U8 ( .A1(n5), .A2(i_data_bus[0]), .B1(n4), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n5), .A2(i_data_bus[1]), .B1(n4), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n5), .A2(i_data_bus[2]), .B1(n4), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n5), .A2(i_data_bus[3]), .B1(n4), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n5), .A2(i_data_bus[4]), .B1(n4), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n5), .A2(i_data_bus[5]), .B1(n4), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n5), .A2(i_data_bus[6]), .B1(n4), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n5), .A2(i_data_bus[7]), .B1(n4), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n5), .A2(i_data_bus[8]), .B1(n4), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n5), .A2(i_data_bus[9]), .B1(n4), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n5), .A2(i_data_bus[10]), .B1(n4), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n5), .A2(i_data_bus[11]), .B1(n4), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n5), .A2(i_data_bus[12]), .B1(n4), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n5), .A2(i_data_bus[13]), .B1(n4), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n5), .A2(i_data_bus[14]), .B1(n4), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n5), .A2(i_data_bus[15]), .B1(n4), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n5), .A2(i_data_bus[16]), .B1(n4), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n5), .A2(i_data_bus[17]), .B1(n4), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n5), .A2(i_data_bus[18]), .B1(n4), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n5), .A2(i_data_bus[19]), .B1(n4), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n5), .A2(i_data_bus[20]), .B1(n4), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n5), .A2(i_data_bus[21]), .B1(n4), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n5), .A2(i_data_bus[22]), .B1(n4), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n5), .A2(i_data_bus[23]), .B1(n4), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n5), .A2(i_data_bus[24]), .B1(n4), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n5), .A2(i_data_bus[25]), .B1(n4), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n5), .A2(i_data_bus[26]), .B1(n4), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n5), .A2(i_data_bus[27]), .B1(n4), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n5), .A2(i_data_bus[28]), .B1(n4), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n5), .A2(i_data_bus[29]), .B1(n4), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n5), .A2(i_data_bus[30]), .B1(n4), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n5), .A2(i_data_bus[31]), .B1(n4), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n5), .A2(n4), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_278 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_278 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_279 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  NR2D2BWP30P140LVT U3 ( .A1(i_cmd[0]), .A2(n3), .ZN(N91) );
  ND2D1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n2) );
  CKAN2D1BWP30P140LVT U5 ( .A1(N91), .A2(i_data_bus[0]), .Z(N92) );
  CKAN2D1BWP30P140LVT U6 ( .A1(N91), .A2(i_data_bus[1]), .Z(N93) );
  CKAN2D1BWP30P140LVT U7 ( .A1(N91), .A2(i_data_bus[2]), .Z(N94) );
  CKAN2D1BWP30P140LVT U8 ( .A1(N91), .A2(i_data_bus[3]), .Z(N95) );
  CKAN2D1BWP30P140LVT U9 ( .A1(N91), .A2(i_data_bus[4]), .Z(N96) );
  CKAN2D1BWP30P140LVT U10 ( .A1(N91), .A2(i_data_bus[5]), .Z(N97) );
  CKAN2D1BWP30P140LVT U11 ( .A1(N91), .A2(i_data_bus[6]), .Z(N98) );
  CKAN2D1BWP30P140LVT U12 ( .A1(N91), .A2(i_data_bus[7]), .Z(N99) );
  CKAN2D1BWP30P140LVT U13 ( .A1(N91), .A2(i_data_bus[8]), .Z(N100) );
  CKAN2D1BWP30P140LVT U14 ( .A1(N91), .A2(i_data_bus[9]), .Z(N101) );
  CKAN2D1BWP30P140LVT U15 ( .A1(N91), .A2(i_data_bus[10]), .Z(N102) );
  CKAN2D1BWP30P140LVT U16 ( .A1(N91), .A2(i_data_bus[11]), .Z(N103) );
  CKAN2D1BWP30P140LVT U17 ( .A1(N91), .A2(i_data_bus[12]), .Z(N104) );
  CKAN2D1BWP30P140LVT U18 ( .A1(N91), .A2(i_data_bus[13]), .Z(N105) );
  CKAN2D1BWP30P140LVT U19 ( .A1(N91), .A2(i_data_bus[14]), .Z(N106) );
  CKAN2D1BWP30P140LVT U20 ( .A1(N91), .A2(i_data_bus[15]), .Z(N107) );
  CKAN2D1BWP30P140LVT U21 ( .A1(N91), .A2(i_data_bus[16]), .Z(N108) );
  CKAN2D1BWP30P140LVT U22 ( .A1(N91), .A2(i_data_bus[17]), .Z(N109) );
  CKAN2D1BWP30P140LVT U23 ( .A1(N91), .A2(i_data_bus[18]), .Z(N110) );
  CKAN2D1BWP30P140LVT U24 ( .A1(N91), .A2(i_data_bus[19]), .Z(N111) );
  CKAN2D1BWP30P140LVT U25 ( .A1(N91), .A2(i_data_bus[20]), .Z(N112) );
  CKAN2D1BWP30P140LVT U26 ( .A1(N91), .A2(i_data_bus[21]), .Z(N113) );
  CKAN2D1BWP30P140LVT U27 ( .A1(N91), .A2(i_data_bus[22]), .Z(N114) );
  CKAN2D1BWP30P140LVT U28 ( .A1(N91), .A2(i_data_bus[23]), .Z(N115) );
  CKAN2D1BWP30P140LVT U29 ( .A1(N91), .A2(i_data_bus[24]), .Z(N116) );
  CKAN2D1BWP30P140LVT U30 ( .A1(N91), .A2(i_data_bus[25]), .Z(N117) );
  CKAN2D1BWP30P140LVT U31 ( .A1(N91), .A2(i_data_bus[26]), .Z(N118) );
  CKAN2D1BWP30P140LVT U32 ( .A1(N91), .A2(i_data_bus[27]), .Z(N119) );
  CKAN2D1BWP30P140LVT U33 ( .A1(N91), .A2(i_data_bus[28]), .Z(N120) );
  CKAN2D1BWP30P140LVT U34 ( .A1(N91), .A2(i_data_bus[29]), .Z(N121) );
  CKAN2D1BWP30P140LVT U35 ( .A1(N91), .A2(i_data_bus[30]), .Z(N122) );
  CKAN2D1BWP30P140LVT U36 ( .A1(N91), .A2(i_data_bus[31]), .Z(N123) );
  IND2D1BWP30P140LVT U37 ( .A1(n2), .B1(n1), .ZN(n3) );
  INVD1BWP30P140LVT U38 ( .I(rst), .ZN(n1) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_279 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   n1;

  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_279 data_mux ( .clk(clk), 
        .rst(rst), .i_valid({n1, i_valid[0]}), .i_data_bus({n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, i_data_bus[31:0]}), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U1 ( .ZN(n1) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_280 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2D1BWP30P140LVT U3 ( .A1(i_en), .A2(i_valid[0]), .ZN(n3) );
  AN2D2BWP30P140LVT U4 ( .A1(i_cmd[0]), .A2(n1), .Z(n5) );
  CKAN2D1BWP30P140LVT U5 ( .A1(i_valid[1]), .A2(n4), .Z(n1) );
  NR3OPTPAD2BWP30P140LVT U6 ( .A1(n3), .A2(i_cmd[0]), .A3(rst), .ZN(n2) );
  INR2D1BWP30P140LVT U7 ( .A1(i_en), .B1(rst), .ZN(n4) );
  AO22D1BWP30P140LVT U8 ( .A1(n2), .A2(i_data_bus[0]), .B1(n5), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U9 ( .A1(n2), .A2(i_data_bus[1]), .B1(n5), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U10 ( .A1(n2), .A2(i_data_bus[2]), .B1(n5), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U11 ( .A1(n2), .A2(i_data_bus[3]), .B1(n5), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U12 ( .A1(n2), .A2(i_data_bus[4]), .B1(n5), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U13 ( .A1(n2), .A2(i_data_bus[5]), .B1(n5), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U14 ( .A1(n2), .A2(i_data_bus[6]), .B1(n5), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U15 ( .A1(n2), .A2(i_data_bus[7]), .B1(n5), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U16 ( .A1(n2), .A2(i_data_bus[8]), .B1(n5), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U17 ( .A1(n2), .A2(i_data_bus[9]), .B1(n5), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U18 ( .A1(n2), .A2(i_data_bus[10]), .B1(n5), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U19 ( .A1(n2), .A2(i_data_bus[11]), .B1(n5), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U20 ( .A1(n2), .A2(i_data_bus[12]), .B1(n5), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U21 ( .A1(n2), .A2(i_data_bus[13]), .B1(n5), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U22 ( .A1(n2), .A2(i_data_bus[14]), .B1(n5), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U23 ( .A1(n2), .A2(i_data_bus[15]), .B1(n5), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U24 ( .A1(n2), .A2(i_data_bus[16]), .B1(n5), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U25 ( .A1(n2), .A2(i_data_bus[17]), .B1(n5), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U26 ( .A1(n2), .A2(i_data_bus[18]), .B1(n5), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U27 ( .A1(n2), .A2(i_data_bus[19]), .B1(n5), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U28 ( .A1(n2), .A2(i_data_bus[20]), .B1(n5), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U29 ( .A1(n2), .A2(i_data_bus[21]), .B1(n5), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U30 ( .A1(n2), .A2(i_data_bus[22]), .B1(n5), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U31 ( .A1(n2), .A2(i_data_bus[23]), .B1(n5), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U32 ( .A1(n2), .A2(i_data_bus[24]), .B1(n5), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U33 ( .A1(n2), .A2(i_data_bus[25]), .B1(n5), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U34 ( .A1(n2), .A2(i_data_bus[26]), .B1(n5), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U35 ( .A1(n2), .A2(i_data_bus[27]), .B1(n5), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U36 ( .A1(n2), .A2(i_data_bus[28]), .B1(n5), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U37 ( .A1(n2), .A2(i_data_bus[29]), .B1(n5), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U38 ( .A1(n2), .A2(i_data_bus[30]), .B1(n5), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U39 ( .A1(n2), .A2(i_data_bus[31]), .B1(n5), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U40 ( .A1(n2), .A2(n5), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_280 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_280 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_281 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  INVD6BWP30P140LVT U3 ( .I(n2), .ZN(n7) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  OR3D4BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .Z(n2) );
  INVD1BWP30P140LVT U6 ( .I(i_valid[1]), .ZN(n5) );
  INR2D1BWP30P140LVT U7 ( .A1(i_en), .B1(rst), .ZN(n3) );
  ND2OPTIBD2BWP30P140LVT U8 ( .A1(i_cmd[0]), .A2(n3), .ZN(n4) );
  NR2OPTPAD2BWP30P140LVT U9 ( .A1(n5), .A2(n4), .ZN(n6) );
  AO22D1BWP30P140LVT U10 ( .A1(n7), .A2(i_data_bus[0]), .B1(n6), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U11 ( .A1(n7), .A2(i_data_bus[1]), .B1(n6), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U12 ( .A1(n7), .A2(i_data_bus[2]), .B1(n6), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U13 ( .A1(n7), .A2(i_data_bus[3]), .B1(n6), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U14 ( .A1(n7), .A2(i_data_bus[4]), .B1(n6), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U15 ( .A1(n7), .A2(i_data_bus[5]), .B1(n6), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U16 ( .A1(n7), .A2(i_data_bus[6]), .B1(n6), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U17 ( .A1(n7), .A2(i_data_bus[7]), .B1(n6), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U18 ( .A1(n7), .A2(i_data_bus[8]), .B1(n6), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U19 ( .A1(n7), .A2(i_data_bus[9]), .B1(n6), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U20 ( .A1(n7), .A2(i_data_bus[10]), .B1(n6), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U21 ( .A1(n7), .A2(i_data_bus[11]), .B1(n6), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U22 ( .A1(n7), .A2(i_data_bus[12]), .B1(n6), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U23 ( .A1(n7), .A2(i_data_bus[13]), .B1(n6), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U24 ( .A1(n7), .A2(i_data_bus[14]), .B1(n6), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U25 ( .A1(n7), .A2(i_data_bus[15]), .B1(n6), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U26 ( .A1(n7), .A2(i_data_bus[16]), .B1(n6), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U27 ( .A1(n7), .A2(i_data_bus[17]), .B1(n6), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U28 ( .A1(n7), .A2(i_data_bus[18]), .B1(n6), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U29 ( .A1(n7), .A2(i_data_bus[19]), .B1(n6), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U30 ( .A1(n7), .A2(i_data_bus[20]), .B1(n6), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U31 ( .A1(n7), .A2(i_data_bus[21]), .B1(n6), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U32 ( .A1(n7), .A2(i_data_bus[22]), .B1(n6), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U33 ( .A1(n7), .A2(i_data_bus[23]), .B1(n6), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U34 ( .A1(n7), .A2(i_data_bus[24]), .B1(n6), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U35 ( .A1(n7), .A2(i_data_bus[25]), .B1(n6), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U36 ( .A1(n7), .A2(i_data_bus[26]), .B1(n6), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U37 ( .A1(n7), .A2(i_data_bus[27]), .B1(n6), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U38 ( .A1(n7), .A2(i_data_bus[28]), .B1(n6), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U39 ( .A1(n7), .A2(i_data_bus[29]), .B1(n6), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U40 ( .A1(n7), .A2(i_data_bus[30]), .B1(n6), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U41 ( .A1(n7), .A2(i_data_bus[31]), .B1(n6), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U42 ( .A1(n7), .A2(n6), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_281 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_281 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_282 ( clk, rst, i_valid, 
        i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, n1, n2, n3, n4,
         n5, n6, n7;

  DFQD1BWP30P140LVT o_valid_inner_reg ( .D(N91), .CP(clk), .Q(o_valid) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N123), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N122), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N121), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N120), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N119), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N118), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N117), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[0]) );
  INVD6BWP30P140LVT U3 ( .I(n2), .ZN(n7) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(i_en), .A2(i_valid[0]), .ZN(n1) );
  OR3D4BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .A3(rst), .Z(n2) );
  INVD1BWP30P140LVT U6 ( .I(i_valid[1]), .ZN(n5) );
  INR2D1BWP30P140LVT U7 ( .A1(i_en), .B1(rst), .ZN(n3) );
  ND2OPTIBD2BWP30P140LVT U8 ( .A1(i_cmd[0]), .A2(n3), .ZN(n4) );
  NR2OPTPAD2BWP30P140LVT U9 ( .A1(n5), .A2(n4), .ZN(n6) );
  AO22D1BWP30P140LVT U10 ( .A1(n7), .A2(i_data_bus[0]), .B1(n6), .B2(
        i_data_bus[32]), .Z(N92) );
  AO22D1BWP30P140LVT U11 ( .A1(n7), .A2(i_data_bus[1]), .B1(n6), .B2(
        i_data_bus[33]), .Z(N93) );
  AO22D1BWP30P140LVT U12 ( .A1(n7), .A2(i_data_bus[2]), .B1(n6), .B2(
        i_data_bus[34]), .Z(N94) );
  AO22D1BWP30P140LVT U13 ( .A1(n7), .A2(i_data_bus[3]), .B1(n6), .B2(
        i_data_bus[35]), .Z(N95) );
  AO22D1BWP30P140LVT U14 ( .A1(n7), .A2(i_data_bus[4]), .B1(n6), .B2(
        i_data_bus[36]), .Z(N96) );
  AO22D1BWP30P140LVT U15 ( .A1(n7), .A2(i_data_bus[5]), .B1(n6), .B2(
        i_data_bus[37]), .Z(N97) );
  AO22D1BWP30P140LVT U16 ( .A1(n7), .A2(i_data_bus[6]), .B1(n6), .B2(
        i_data_bus[38]), .Z(N98) );
  AO22D1BWP30P140LVT U17 ( .A1(n7), .A2(i_data_bus[7]), .B1(n6), .B2(
        i_data_bus[39]), .Z(N99) );
  AO22D1BWP30P140LVT U18 ( .A1(n7), .A2(i_data_bus[8]), .B1(n6), .B2(
        i_data_bus[40]), .Z(N100) );
  AO22D1BWP30P140LVT U19 ( .A1(n7), .A2(i_data_bus[9]), .B1(n6), .B2(
        i_data_bus[41]), .Z(N101) );
  AO22D1BWP30P140LVT U20 ( .A1(n7), .A2(i_data_bus[10]), .B1(n6), .B2(
        i_data_bus[42]), .Z(N102) );
  AO22D1BWP30P140LVT U21 ( .A1(n7), .A2(i_data_bus[11]), .B1(n6), .B2(
        i_data_bus[43]), .Z(N103) );
  AO22D1BWP30P140LVT U22 ( .A1(n7), .A2(i_data_bus[12]), .B1(n6), .B2(
        i_data_bus[44]), .Z(N104) );
  AO22D1BWP30P140LVT U23 ( .A1(n7), .A2(i_data_bus[13]), .B1(n6), .B2(
        i_data_bus[45]), .Z(N105) );
  AO22D1BWP30P140LVT U24 ( .A1(n7), .A2(i_data_bus[14]), .B1(n6), .B2(
        i_data_bus[46]), .Z(N106) );
  AO22D1BWP30P140LVT U25 ( .A1(n7), .A2(i_data_bus[15]), .B1(n6), .B2(
        i_data_bus[47]), .Z(N107) );
  AO22D1BWP30P140LVT U26 ( .A1(n7), .A2(i_data_bus[16]), .B1(n6), .B2(
        i_data_bus[48]), .Z(N108) );
  AO22D1BWP30P140LVT U27 ( .A1(n7), .A2(i_data_bus[17]), .B1(n6), .B2(
        i_data_bus[49]), .Z(N109) );
  AO22D1BWP30P140LVT U28 ( .A1(n7), .A2(i_data_bus[18]), .B1(n6), .B2(
        i_data_bus[50]), .Z(N110) );
  AO22D1BWP30P140LVT U29 ( .A1(n7), .A2(i_data_bus[19]), .B1(n6), .B2(
        i_data_bus[51]), .Z(N111) );
  AO22D1BWP30P140LVT U30 ( .A1(n7), .A2(i_data_bus[20]), .B1(n6), .B2(
        i_data_bus[52]), .Z(N112) );
  AO22D1BWP30P140LVT U31 ( .A1(n7), .A2(i_data_bus[21]), .B1(n6), .B2(
        i_data_bus[53]), .Z(N113) );
  AO22D1BWP30P140LVT U32 ( .A1(n7), .A2(i_data_bus[22]), .B1(n6), .B2(
        i_data_bus[54]), .Z(N114) );
  AO22D1BWP30P140LVT U33 ( .A1(n7), .A2(i_data_bus[23]), .B1(n6), .B2(
        i_data_bus[55]), .Z(N115) );
  AO22D1BWP30P140LVT U34 ( .A1(n7), .A2(i_data_bus[24]), .B1(n6), .B2(
        i_data_bus[56]), .Z(N116) );
  AO22D1BWP30P140LVT U35 ( .A1(n7), .A2(i_data_bus[25]), .B1(n6), .B2(
        i_data_bus[57]), .Z(N117) );
  AO22D1BWP30P140LVT U36 ( .A1(n7), .A2(i_data_bus[26]), .B1(n6), .B2(
        i_data_bus[58]), .Z(N118) );
  AO22D1BWP30P140LVT U37 ( .A1(n7), .A2(i_data_bus[27]), .B1(n6), .B2(
        i_data_bus[59]), .Z(N119) );
  AO22D1BWP30P140LVT U38 ( .A1(n7), .A2(i_data_bus[28]), .B1(n6), .B2(
        i_data_bus[60]), .Z(N120) );
  AO22D1BWP30P140LVT U39 ( .A1(n7), .A2(i_data_bus[29]), .B1(n6), .B2(
        i_data_bus[61]), .Z(N121) );
  AO22D1BWP30P140LVT U40 ( .A1(n7), .A2(i_data_bus[30]), .B1(n6), .B2(
        i_data_bus[62]), .Z(N122) );
  AO22D1BWP30P140LVT U41 ( .A1(n7), .A2(i_data_bus[31]), .B1(n6), .B2(
        i_data_bus[63]), .Z(N123) );
  OR2D1BWP30P140LVT U42 ( .A1(n7), .A2(n6), .Z(N91) );
endmodule


module merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_282 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input [0:0] i_cmd;
  input clk, rst, i_en;
  output o_valid;


  mux_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_282 data_mux ( .clk(clk), 
        .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), .o_valid(
        o_valid), .o_data_bus(o_data_bus), .i_en(i_en), .i_cmd(i_cmd[0]) );
endmodule


module distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_47 ( clk, rst, 
        i_valid, i_data_bus, o_valid, o_data_bus, i_fwd_valid, i_fwd_data_bus, 
        o_fwd_valid, o_fwd_data_bus, i_en, i_cmd );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [1:0] o_valid;
  output [63:0] o_data_bus;
  input [31:0] i_fwd_data_bus;
  output [31:0] o_fwd_data_bus;
  input [4:0] i_cmd;
  input clk, rst, i_fwd_valid, i_en;
  output o_fwd_valid;
  wire   n_Logic0_, inner_fwd_valid, n_3_net_;
  wire   [1:0] inner_valid;
  wire   [63:0] inner_data_bus;
  wire   [31:0] inner_fwd_data_bus;

  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_282 merge_i_data_high ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[1]), .o_data_bus(inner_data_bus[63:32]), .i_en(
        i_en), .i_cmd(i_cmd[4]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_281 merge_i_data_low ( 
        .clk(clk), .rst(rst), .i_valid(i_valid), .i_data_bus(i_data_bus), 
        .o_valid(inner_valid[0]), .o_data_bus(inner_data_bus[31:0]), .i_en(
        i_en), .i_cmd(i_cmd[3]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_280 o_fwd ( .clk(clk), 
        .rst(rst), .i_valid(inner_valid), .i_data_bus(inner_data_bus), 
        .o_valid(inner_fwd_valid), .o_data_bus(inner_fwd_data_bus), .i_en(i_en), .i_cmd(i_cmd[2]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_279 o_fwd_en ( .clk(clk), 
        .rst(rst), .i_valid({n_Logic0_, inner_fwd_valid}), .i_data_bus({
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, inner_fwd_data_bus}), .o_valid(o_fwd_valid), 
        .o_data_bus(o_fwd_data_bus), .i_en(i_en), .i_cmd(n_3_net_) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_278 o_data_high ( .clk(clk), .rst(rst), .i_valid({inner_valid[1], i_fwd_valid}), .i_data_bus({
        inner_data_bus[63:32], i_fwd_data_bus}), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(i_cmd[1]) );
  merge_2x1_simple_seq_DATA_WIDTH32_COMMAND_WIDTH1_277 o_data_low ( .clk(clk), 
        .rst(rst), .i_valid({inner_valid[0], i_fwd_valid}), .i_data_bus({
        inner_data_bus[31:0], i_fwd_data_bus}), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(i_cmd[0]) );
  TIELBWP30P140LVT U2 ( .ZN(n_Logic0_) );
  CKAN2D1BWP30P140LVT U3 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n_3_net_) );
endmodule


module flatten_benes_simple_seq ( clk, rst, i_valid, i_data_bus, o_valid, 
        o_data_bus, i_en, i_cmd );
  input [15:0] i_valid;
  input [511:0] i_data_bus;
  output [15:0] o_valid;
  output [511:0] o_data_bus;
  input [279:0] i_cmd;
  input clk, rst, i_en;
  wire   n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__0__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__0__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__0__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__0__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__0__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__1__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__1__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__1__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__1__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__1__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__2__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__2__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__2__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__2__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__2__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__3__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__3__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__3__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__3__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__3__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__4__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__4__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__4__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__4__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__4__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__5__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__5__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__5__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__5__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__5__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__6__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__6__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__6__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__6__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__6__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__7__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__7__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__7__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__7__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__7__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__0__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__0__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__0__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__0__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__0__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__1__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__1__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__1__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__1__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__1__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__2__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__2__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__2__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__2__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__2__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__3__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__3__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__3__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__3__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__3__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__4__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__4__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__4__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__4__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__4__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__5__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__5__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__5__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__5__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__5__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__6__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__6__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__6__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__6__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__6__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__7__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__7__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__7__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__7__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__7__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__0__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__0__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__1__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__1__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__2__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__2__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__3__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__3__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__4__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__4__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__5__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__5__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__6__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__6__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__7__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__7__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__0__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__0__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__0__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__0__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__0__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__1__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__1__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__1__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__1__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__1__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__2__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__2__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__2__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__2__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__2__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__3__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__3__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__3__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__3__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__3__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__4__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__4__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__4__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__4__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__4__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__5__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__5__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__5__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__5__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__5__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__6__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__6__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__6__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__6__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__6__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__7__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__7__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__7__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__7__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__7__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__0__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__0__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__0__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__0__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__0__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__1__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__1__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__1__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__1__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__1__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__2__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__2__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__2__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__2__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__2__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__3__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__3__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__3__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__3__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__3__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__4__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__4__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__4__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__4__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__4__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__5__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__5__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__5__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__5__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__5__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__6__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__6__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__6__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__6__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__6__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__7__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__7__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__7__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__7__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__7__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__0__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__0__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__0__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__0__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__0__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__1__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__1__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__1__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__1__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__1__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__2__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__2__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__2__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__2__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__2__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__3__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__3__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__3__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__3__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__3__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__4__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__4__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__4__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__4__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__4__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__5__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__5__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__5__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__5__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__5__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__6__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__6__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__6__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__6__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__6__0_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__7__4_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__7__3_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__7__2_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__7__1_,
         cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__7__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__0__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__0__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__0__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__0__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__0__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__1__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__1__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__1__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__1__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__1__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__2__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__2__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__2__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__2__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__2__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__3__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__3__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__3__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__3__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__3__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__4__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__4__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__4__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__4__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__4__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__5__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__5__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__5__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__5__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__5__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__6__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__6__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__6__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__6__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__6__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__7__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__7__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__7__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__7__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__7__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__0__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__0__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__1__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__1__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__2__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__2__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__3__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__3__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__4__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__4__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__5__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__5__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__6__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__6__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__7__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__7__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__0__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__0__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__0__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__0__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__0__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__1__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__1__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__1__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__1__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__1__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__2__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__2__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__2__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__2__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__2__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__3__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__3__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__3__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__3__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__3__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__4__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__4__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__4__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__4__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__4__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__5__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__5__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__5__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__5__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__5__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__6__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__6__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__6__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__6__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__6__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__7__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__7__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__7__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__7__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__7__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__0__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__0__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__0__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__0__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__0__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__1__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__1__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__1__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__1__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__1__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__2__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__2__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__2__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__2__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__2__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__3__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__3__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__3__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__3__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__3__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__4__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__4__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__4__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__4__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__4__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__5__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__5__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__5__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__5__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__5__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__6__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__6__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__6__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__6__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__6__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__7__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__7__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__7__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__7__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__7__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__0__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__0__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__0__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__0__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__0__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__1__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__1__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__1__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__1__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__1__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__2__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__2__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__2__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__2__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__2__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__3__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__3__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__3__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__3__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__3__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__4__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__4__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__4__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__4__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__4__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__5__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__5__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__5__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__5__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__5__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__6__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__6__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__6__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__6__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__6__0_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__7__4_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__7__3_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__7__2_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__7__1_,
         cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__7__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__0__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__0__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__1__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__1__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__2__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__2__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__3__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__3__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__4__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__4__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__5__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__5__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__6__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__6__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__7__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__7__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__0__4_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__0__3_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__0__2_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__0__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__0__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__1__4_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__1__3_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__1__2_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__1__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__1__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__2__4_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__2__3_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__2__2_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__2__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__2__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__3__4_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__3__3_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__3__2_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__3__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__3__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__4__4_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__4__3_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__4__2_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__4__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__4__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__5__4_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__5__3_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__5__2_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__5__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__5__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__6__4_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__6__3_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__6__2_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__6__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__6__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__7__4_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__7__3_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__7__2_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__7__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__7__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__0__4_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__0__3_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__0__2_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__0__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__0__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__1__4_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__1__3_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__1__2_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__1__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__1__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__2__4_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__2__3_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__2__2_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__2__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__2__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__3__4_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__3__3_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__3__2_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__3__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__3__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__4__4_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__4__3_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__4__2_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__4__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__4__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__5__4_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__5__3_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__5__2_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__5__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__5__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__6__4_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__6__3_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__6__2_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__6__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__6__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__7__4_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__7__3_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__7__2_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__7__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__7__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__0__4_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__0__3_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__0__2_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__0__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__0__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__1__4_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__1__3_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__1__2_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__1__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__1__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__2__4_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__2__3_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__2__2_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__2__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__2__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__3__4_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__3__3_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__3__2_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__3__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__3__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__4__4_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__4__3_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__4__2_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__4__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__4__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__5__4_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__5__3_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__5__2_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__5__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__5__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__6__4_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__6__3_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__6__2_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__6__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__6__0_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__7__4_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__7__3_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__7__2_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__7__1_,
         cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__7__0_,
         connection_0__0__31_, connection_0__0__30_, connection_0__0__29_,
         connection_0__0__28_, connection_0__0__27_, connection_0__0__26_,
         connection_0__0__25_, connection_0__0__24_, connection_0__0__23_,
         connection_0__0__22_, connection_0__0__21_, connection_0__0__20_,
         connection_0__0__19_, connection_0__0__18_, connection_0__0__17_,
         connection_0__0__16_, connection_0__0__15_, connection_0__0__14_,
         connection_0__0__13_, connection_0__0__12_, connection_0__0__11_,
         connection_0__0__10_, connection_0__0__9_, connection_0__0__8_,
         connection_0__0__7_, connection_0__0__6_, connection_0__0__5_,
         connection_0__0__4_, connection_0__0__3_, connection_0__0__2_,
         connection_0__0__1_, connection_0__0__0_, connection_0__1__31_,
         connection_0__1__30_, connection_0__1__29_, connection_0__1__28_,
         connection_0__1__27_, connection_0__1__26_, connection_0__1__25_,
         connection_0__1__24_, connection_0__1__23_, connection_0__1__22_,
         connection_0__1__21_, connection_0__1__20_, connection_0__1__19_,
         connection_0__1__18_, connection_0__1__17_, connection_0__1__16_,
         connection_0__1__15_, connection_0__1__14_, connection_0__1__13_,
         connection_0__1__12_, connection_0__1__11_, connection_0__1__10_,
         connection_0__1__9_, connection_0__1__8_, connection_0__1__7_,
         connection_0__1__6_, connection_0__1__5_, connection_0__1__4_,
         connection_0__1__3_, connection_0__1__2_, connection_0__1__1_,
         connection_0__1__0_, connection_0__2__31_, connection_0__2__30_,
         connection_0__2__29_, connection_0__2__28_, connection_0__2__27_,
         connection_0__2__26_, connection_0__2__25_, connection_0__2__24_,
         connection_0__2__23_, connection_0__2__22_, connection_0__2__21_,
         connection_0__2__20_, connection_0__2__19_, connection_0__2__18_,
         connection_0__2__17_, connection_0__2__16_, connection_0__2__15_,
         connection_0__2__14_, connection_0__2__13_, connection_0__2__12_,
         connection_0__2__11_, connection_0__2__10_, connection_0__2__9_,
         connection_0__2__8_, connection_0__2__7_, connection_0__2__6_,
         connection_0__2__5_, connection_0__2__4_, connection_0__2__3_,
         connection_0__2__2_, connection_0__2__1_, connection_0__2__0_,
         connection_0__3__31_, connection_0__3__30_, connection_0__3__29_,
         connection_0__3__28_, connection_0__3__27_, connection_0__3__26_,
         connection_0__3__25_, connection_0__3__24_, connection_0__3__23_,
         connection_0__3__22_, connection_0__3__21_, connection_0__3__20_,
         connection_0__3__19_, connection_0__3__18_, connection_0__3__17_,
         connection_0__3__16_, connection_0__3__15_, connection_0__3__14_,
         connection_0__3__13_, connection_0__3__12_, connection_0__3__11_,
         connection_0__3__10_, connection_0__3__9_, connection_0__3__8_,
         connection_0__3__7_, connection_0__3__6_, connection_0__3__5_,
         connection_0__3__4_, connection_0__3__3_, connection_0__3__2_,
         connection_0__3__1_, connection_0__3__0_, connection_0__4__31_,
         connection_0__4__30_, connection_0__4__29_, connection_0__4__28_,
         connection_0__4__27_, connection_0__4__26_, connection_0__4__25_,
         connection_0__4__24_, connection_0__4__23_, connection_0__4__22_,
         connection_0__4__21_, connection_0__4__20_, connection_0__4__19_,
         connection_0__4__18_, connection_0__4__17_, connection_0__4__16_,
         connection_0__4__15_, connection_0__4__14_, connection_0__4__13_,
         connection_0__4__12_, connection_0__4__11_, connection_0__4__10_,
         connection_0__4__9_, connection_0__4__8_, connection_0__4__7_,
         connection_0__4__6_, connection_0__4__5_, connection_0__4__4_,
         connection_0__4__3_, connection_0__4__2_, connection_0__4__1_,
         connection_0__4__0_, connection_0__5__31_, connection_0__5__30_,
         connection_0__5__29_, connection_0__5__28_, connection_0__5__27_,
         connection_0__5__26_, connection_0__5__25_, connection_0__5__24_,
         connection_0__5__23_, connection_0__5__22_, connection_0__5__21_,
         connection_0__5__20_, connection_0__5__19_, connection_0__5__18_,
         connection_0__5__17_, connection_0__5__16_, connection_0__5__15_,
         connection_0__5__14_, connection_0__5__13_, connection_0__5__12_,
         connection_0__5__11_, connection_0__5__10_, connection_0__5__9_,
         connection_0__5__8_, connection_0__5__7_, connection_0__5__6_,
         connection_0__5__5_, connection_0__5__4_, connection_0__5__3_,
         connection_0__5__2_, connection_0__5__1_, connection_0__5__0_,
         connection_0__6__31_, connection_0__6__30_, connection_0__6__29_,
         connection_0__6__28_, connection_0__6__27_, connection_0__6__26_,
         connection_0__6__25_, connection_0__6__24_, connection_0__6__23_,
         connection_0__6__22_, connection_0__6__21_, connection_0__6__20_,
         connection_0__6__19_, connection_0__6__18_, connection_0__6__17_,
         connection_0__6__16_, connection_0__6__15_, connection_0__6__14_,
         connection_0__6__13_, connection_0__6__12_, connection_0__6__11_,
         connection_0__6__10_, connection_0__6__9_, connection_0__6__8_,
         connection_0__6__7_, connection_0__6__6_, connection_0__6__5_,
         connection_0__6__4_, connection_0__6__3_, connection_0__6__2_,
         connection_0__6__1_, connection_0__6__0_, connection_0__7__31_,
         connection_0__7__30_, connection_0__7__29_, connection_0__7__28_,
         connection_0__7__27_, connection_0__7__26_, connection_0__7__25_,
         connection_0__7__24_, connection_0__7__23_, connection_0__7__22_,
         connection_0__7__21_, connection_0__7__20_, connection_0__7__19_,
         connection_0__7__18_, connection_0__7__17_, connection_0__7__16_,
         connection_0__7__15_, connection_0__7__14_, connection_0__7__13_,
         connection_0__7__12_, connection_0__7__11_, connection_0__7__10_,
         connection_0__7__9_, connection_0__7__8_, connection_0__7__7_,
         connection_0__7__6_, connection_0__7__5_, connection_0__7__4_,
         connection_0__7__3_, connection_0__7__2_, connection_0__7__1_,
         connection_0__7__0_, connection_0__8__31_, connection_0__8__30_,
         connection_0__8__29_, connection_0__8__28_, connection_0__8__27_,
         connection_0__8__26_, connection_0__8__25_, connection_0__8__24_,
         connection_0__8__23_, connection_0__8__22_, connection_0__8__21_,
         connection_0__8__20_, connection_0__8__19_, connection_0__8__18_,
         connection_0__8__17_, connection_0__8__16_, connection_0__8__15_,
         connection_0__8__14_, connection_0__8__13_, connection_0__8__12_,
         connection_0__8__11_, connection_0__8__10_, connection_0__8__9_,
         connection_0__8__8_, connection_0__8__7_, connection_0__8__6_,
         connection_0__8__5_, connection_0__8__4_, connection_0__8__3_,
         connection_0__8__2_, connection_0__8__1_, connection_0__8__0_,
         connection_0__9__31_, connection_0__9__30_, connection_0__9__29_,
         connection_0__9__28_, connection_0__9__27_, connection_0__9__26_,
         connection_0__9__25_, connection_0__9__24_, connection_0__9__23_,
         connection_0__9__22_, connection_0__9__21_, connection_0__9__20_,
         connection_0__9__19_, connection_0__9__18_, connection_0__9__17_,
         connection_0__9__16_, connection_0__9__15_, connection_0__9__14_,
         connection_0__9__13_, connection_0__9__12_, connection_0__9__11_,
         connection_0__9__10_, connection_0__9__9_, connection_0__9__8_,
         connection_0__9__7_, connection_0__9__6_, connection_0__9__5_,
         connection_0__9__4_, connection_0__9__3_, connection_0__9__2_,
         connection_0__9__1_, connection_0__9__0_, connection_0__10__31_,
         connection_0__10__30_, connection_0__10__29_, connection_0__10__28_,
         connection_0__10__27_, connection_0__10__26_, connection_0__10__25_,
         connection_0__10__24_, connection_0__10__23_, connection_0__10__22_,
         connection_0__10__21_, connection_0__10__20_, connection_0__10__19_,
         connection_0__10__18_, connection_0__10__17_, connection_0__10__16_,
         connection_0__10__15_, connection_0__10__14_, connection_0__10__13_,
         connection_0__10__12_, connection_0__10__11_, connection_0__10__10_,
         connection_0__10__9_, connection_0__10__8_, connection_0__10__7_,
         connection_0__10__6_, connection_0__10__5_, connection_0__10__4_,
         connection_0__10__3_, connection_0__10__2_, connection_0__10__1_,
         connection_0__10__0_, connection_0__11__31_, connection_0__11__30_,
         connection_0__11__29_, connection_0__11__28_, connection_0__11__27_,
         connection_0__11__26_, connection_0__11__25_, connection_0__11__24_,
         connection_0__11__23_, connection_0__11__22_, connection_0__11__21_,
         connection_0__11__20_, connection_0__11__19_, connection_0__11__18_,
         connection_0__11__17_, connection_0__11__16_, connection_0__11__15_,
         connection_0__11__14_, connection_0__11__13_, connection_0__11__12_,
         connection_0__11__11_, connection_0__11__10_, connection_0__11__9_,
         connection_0__11__8_, connection_0__11__7_, connection_0__11__6_,
         connection_0__11__5_, connection_0__11__4_, connection_0__11__3_,
         connection_0__11__2_, connection_0__11__1_, connection_0__11__0_,
         connection_0__12__31_, connection_0__12__30_, connection_0__12__29_,
         connection_0__12__28_, connection_0__12__27_, connection_0__12__26_,
         connection_0__12__25_, connection_0__12__24_, connection_0__12__23_,
         connection_0__12__22_, connection_0__12__21_, connection_0__12__20_,
         connection_0__12__19_, connection_0__12__18_, connection_0__12__17_,
         connection_0__12__16_, connection_0__12__15_, connection_0__12__14_,
         connection_0__12__13_, connection_0__12__12_, connection_0__12__11_,
         connection_0__12__10_, connection_0__12__9_, connection_0__12__8_,
         connection_0__12__7_, connection_0__12__6_, connection_0__12__5_,
         connection_0__12__4_, connection_0__12__3_, connection_0__12__2_,
         connection_0__12__1_, connection_0__12__0_, connection_0__13__31_,
         connection_0__13__30_, connection_0__13__29_, connection_0__13__28_,
         connection_0__13__27_, connection_0__13__26_, connection_0__13__25_,
         connection_0__13__24_, connection_0__13__23_, connection_0__13__22_,
         connection_0__13__21_, connection_0__13__20_, connection_0__13__19_,
         connection_0__13__18_, connection_0__13__17_, connection_0__13__16_,
         connection_0__13__15_, connection_0__13__14_, connection_0__13__13_,
         connection_0__13__12_, connection_0__13__11_, connection_0__13__10_,
         connection_0__13__9_, connection_0__13__8_, connection_0__13__7_,
         connection_0__13__6_, connection_0__13__5_, connection_0__13__4_,
         connection_0__13__3_, connection_0__13__2_, connection_0__13__1_,
         connection_0__13__0_, connection_0__14__31_, connection_0__14__30_,
         connection_0__14__29_, connection_0__14__28_, connection_0__14__27_,
         connection_0__14__26_, connection_0__14__25_, connection_0__14__24_,
         connection_0__14__23_, connection_0__14__22_, connection_0__14__21_,
         connection_0__14__20_, connection_0__14__19_, connection_0__14__18_,
         connection_0__14__17_, connection_0__14__16_, connection_0__14__15_,
         connection_0__14__14_, connection_0__14__13_, connection_0__14__12_,
         connection_0__14__11_, connection_0__14__10_, connection_0__14__9_,
         connection_0__14__8_, connection_0__14__7_, connection_0__14__6_,
         connection_0__14__5_, connection_0__14__4_, connection_0__14__3_,
         connection_0__14__2_, connection_0__14__1_, connection_0__14__0_,
         connection_0__15__31_, connection_0__15__30_, connection_0__15__29_,
         connection_0__15__28_, connection_0__15__27_, connection_0__15__26_,
         connection_0__15__25_, connection_0__15__24_, connection_0__15__23_,
         connection_0__15__22_, connection_0__15__21_, connection_0__15__20_,
         connection_0__15__19_, connection_0__15__18_, connection_0__15__17_,
         connection_0__15__16_, connection_0__15__15_, connection_0__15__14_,
         connection_0__15__13_, connection_0__15__12_, connection_0__15__11_,
         connection_0__15__10_, connection_0__15__9_, connection_0__15__8_,
         connection_0__15__7_, connection_0__15__6_, connection_0__15__5_,
         connection_0__15__4_, connection_0__15__3_, connection_0__15__2_,
         connection_0__15__1_, connection_0__15__0_, connection_valid_0__0_,
         connection_valid_0__1_, connection_valid_0__2_,
         connection_valid_0__3_, connection_valid_0__4_,
         connection_valid_0__5_, connection_valid_0__6_,
         connection_valid_0__7_, connection_valid_0__8_,
         connection_valid_0__9_, connection_valid_0__10_,
         connection_valid_0__11_, connection_valid_0__12_,
         connection_valid_0__13_, connection_valid_0__14_,
         connection_valid_0__15_, connection_valid_1__0_,
         connection_valid_1__1_, connection_valid_1__2_,
         connection_valid_1__3_, connection_valid_1__4_,
         connection_valid_1__5_, connection_valid_1__6_,
         connection_valid_1__7_, connection_valid_1__8_,
         connection_valid_1__9_, connection_valid_1__10_,
         connection_valid_1__11_, connection_valid_1__12_,
         connection_valid_1__13_, connection_valid_1__14_,
         connection_valid_1__15_, connection_valid_2__0_,
         connection_valid_2__1_, connection_valid_2__2_,
         connection_valid_2__3_, connection_valid_2__4_,
         connection_valid_2__5_, connection_valid_2__6_,
         connection_valid_2__7_, connection_valid_2__8_,
         connection_valid_2__9_, connection_valid_2__10_,
         connection_valid_2__11_, connection_valid_2__12_,
         connection_valid_2__13_, connection_valid_2__14_,
         connection_valid_2__15_, connection_valid_3__0_,
         connection_valid_3__1_, connection_valid_3__2_,
         connection_valid_3__3_, connection_valid_3__4_,
         connection_valid_3__5_, connection_valid_3__6_,
         connection_valid_3__7_, connection_valid_3__8_,
         connection_valid_3__9_, connection_valid_3__10_,
         connection_valid_3__11_, connection_valid_3__12_,
         connection_valid_3__13_, connection_valid_3__14_,
         connection_valid_3__15_, connection_valid_4__0_,
         connection_valid_4__1_, connection_valid_4__2_,
         connection_valid_4__3_, connection_valid_4__4_,
         connection_valid_4__5_, connection_valid_4__6_,
         connection_valid_4__7_, connection_valid_4__8_,
         connection_valid_4__9_, connection_valid_4__10_,
         connection_valid_4__11_, connection_valid_4__12_,
         connection_valid_4__13_, connection_valid_4__14_,
         connection_valid_4__15_, connection_valid_5__0_,
         connection_valid_5__1_, connection_valid_5__2_,
         connection_valid_5__3_, connection_valid_5__4_,
         connection_valid_5__5_, connection_valid_5__6_,
         connection_valid_5__7_, connection_valid_5__8_,
         connection_valid_5__9_, connection_valid_5__10_,
         connection_valid_5__11_, connection_valid_5__12_,
         connection_valid_5__13_, connection_valid_5__14_,
         connection_valid_5__15_, connection_1__0__31_, connection_1__0__30_,
         connection_1__0__29_, connection_1__0__28_, connection_1__0__27_,
         connection_1__0__26_, connection_1__0__25_, connection_1__0__24_,
         connection_1__0__23_, connection_1__0__22_, connection_1__0__21_,
         connection_1__0__20_, connection_1__0__19_, connection_1__0__18_,
         connection_1__0__17_, connection_1__0__16_, connection_1__0__15_,
         connection_1__0__14_, connection_1__0__13_, connection_1__0__12_,
         connection_1__0__11_, connection_1__0__10_, connection_1__0__9_,
         connection_1__0__8_, connection_1__0__7_, connection_1__0__6_,
         connection_1__0__5_, connection_1__0__4_, connection_1__0__3_,
         connection_1__0__2_, connection_1__0__1_, connection_1__0__0_,
         connection_1__1__31_, connection_1__1__30_, connection_1__1__29_,
         connection_1__1__28_, connection_1__1__27_, connection_1__1__26_,
         connection_1__1__25_, connection_1__1__24_, connection_1__1__23_,
         connection_1__1__22_, connection_1__1__21_, connection_1__1__20_,
         connection_1__1__19_, connection_1__1__18_, connection_1__1__17_,
         connection_1__1__16_, connection_1__1__15_, connection_1__1__14_,
         connection_1__1__13_, connection_1__1__12_, connection_1__1__11_,
         connection_1__1__10_, connection_1__1__9_, connection_1__1__8_,
         connection_1__1__7_, connection_1__1__6_, connection_1__1__5_,
         connection_1__1__4_, connection_1__1__3_, connection_1__1__2_,
         connection_1__1__1_, connection_1__1__0_, connection_1__2__31_,
         connection_1__2__30_, connection_1__2__29_, connection_1__2__28_,
         connection_1__2__27_, connection_1__2__26_, connection_1__2__25_,
         connection_1__2__24_, connection_1__2__23_, connection_1__2__22_,
         connection_1__2__21_, connection_1__2__20_, connection_1__2__19_,
         connection_1__2__18_, connection_1__2__17_, connection_1__2__16_,
         connection_1__2__15_, connection_1__2__14_, connection_1__2__13_,
         connection_1__2__12_, connection_1__2__11_, connection_1__2__10_,
         connection_1__2__9_, connection_1__2__8_, connection_1__2__7_,
         connection_1__2__6_, connection_1__2__5_, connection_1__2__4_,
         connection_1__2__3_, connection_1__2__2_, connection_1__2__1_,
         connection_1__2__0_, connection_1__3__31_, connection_1__3__30_,
         connection_1__3__29_, connection_1__3__28_, connection_1__3__27_,
         connection_1__3__26_, connection_1__3__25_, connection_1__3__24_,
         connection_1__3__23_, connection_1__3__22_, connection_1__3__21_,
         connection_1__3__20_, connection_1__3__19_, connection_1__3__18_,
         connection_1__3__17_, connection_1__3__16_, connection_1__3__15_,
         connection_1__3__14_, connection_1__3__13_, connection_1__3__12_,
         connection_1__3__11_, connection_1__3__10_, connection_1__3__9_,
         connection_1__3__8_, connection_1__3__7_, connection_1__3__6_,
         connection_1__3__5_, connection_1__3__4_, connection_1__3__3_,
         connection_1__3__2_, connection_1__3__1_, connection_1__3__0_,
         connection_1__4__31_, connection_1__4__30_, connection_1__4__29_,
         connection_1__4__28_, connection_1__4__27_, connection_1__4__26_,
         connection_1__4__25_, connection_1__4__24_, connection_1__4__23_,
         connection_1__4__22_, connection_1__4__21_, connection_1__4__20_,
         connection_1__4__19_, connection_1__4__18_, connection_1__4__17_,
         connection_1__4__16_, connection_1__4__15_, connection_1__4__14_,
         connection_1__4__13_, connection_1__4__12_, connection_1__4__11_,
         connection_1__4__10_, connection_1__4__9_, connection_1__4__8_,
         connection_1__4__7_, connection_1__4__6_, connection_1__4__5_,
         connection_1__4__4_, connection_1__4__3_, connection_1__4__2_,
         connection_1__4__1_, connection_1__4__0_, connection_1__5__31_,
         connection_1__5__30_, connection_1__5__29_, connection_1__5__28_,
         connection_1__5__27_, connection_1__5__26_, connection_1__5__25_,
         connection_1__5__24_, connection_1__5__23_, connection_1__5__22_,
         connection_1__5__21_, connection_1__5__20_, connection_1__5__19_,
         connection_1__5__18_, connection_1__5__17_, connection_1__5__16_,
         connection_1__5__15_, connection_1__5__14_, connection_1__5__13_,
         connection_1__5__12_, connection_1__5__11_, connection_1__5__10_,
         connection_1__5__9_, connection_1__5__8_, connection_1__5__7_,
         connection_1__5__6_, connection_1__5__5_, connection_1__5__4_,
         connection_1__5__3_, connection_1__5__2_, connection_1__5__1_,
         connection_1__5__0_, connection_1__6__31_, connection_1__6__30_,
         connection_1__6__29_, connection_1__6__28_, connection_1__6__27_,
         connection_1__6__26_, connection_1__6__25_, connection_1__6__24_,
         connection_1__6__23_, connection_1__6__22_, connection_1__6__21_,
         connection_1__6__20_, connection_1__6__19_, connection_1__6__18_,
         connection_1__6__17_, connection_1__6__16_, connection_1__6__15_,
         connection_1__6__14_, connection_1__6__13_, connection_1__6__12_,
         connection_1__6__11_, connection_1__6__10_, connection_1__6__9_,
         connection_1__6__8_, connection_1__6__7_, connection_1__6__6_,
         connection_1__6__5_, connection_1__6__4_, connection_1__6__3_,
         connection_1__6__2_, connection_1__6__1_, connection_1__6__0_,
         connection_1__7__31_, connection_1__7__30_, connection_1__7__29_,
         connection_1__7__28_, connection_1__7__27_, connection_1__7__26_,
         connection_1__7__25_, connection_1__7__24_, connection_1__7__23_,
         connection_1__7__22_, connection_1__7__21_, connection_1__7__20_,
         connection_1__7__19_, connection_1__7__18_, connection_1__7__17_,
         connection_1__7__16_, connection_1__7__15_, connection_1__7__14_,
         connection_1__7__13_, connection_1__7__12_, connection_1__7__11_,
         connection_1__7__10_, connection_1__7__9_, connection_1__7__8_,
         connection_1__7__7_, connection_1__7__6_, connection_1__7__5_,
         connection_1__7__4_, connection_1__7__3_, connection_1__7__2_,
         connection_1__7__1_, connection_1__7__0_, connection_1__8__31_,
         connection_1__8__30_, connection_1__8__29_, connection_1__8__28_,
         connection_1__8__27_, connection_1__8__26_, connection_1__8__25_,
         connection_1__8__24_, connection_1__8__23_, connection_1__8__22_,
         connection_1__8__21_, connection_1__8__20_, connection_1__8__19_,
         connection_1__8__18_, connection_1__8__17_, connection_1__8__16_,
         connection_1__8__15_, connection_1__8__14_, connection_1__8__13_,
         connection_1__8__12_, connection_1__8__11_, connection_1__8__10_,
         connection_1__8__9_, connection_1__8__8_, connection_1__8__7_,
         connection_1__8__6_, connection_1__8__5_, connection_1__8__4_,
         connection_1__8__3_, connection_1__8__2_, connection_1__8__1_,
         connection_1__8__0_, connection_1__9__31_, connection_1__9__30_,
         connection_1__9__29_, connection_1__9__28_, connection_1__9__27_,
         connection_1__9__26_, connection_1__9__25_, connection_1__9__24_,
         connection_1__9__23_, connection_1__9__22_, connection_1__9__21_,
         connection_1__9__20_, connection_1__9__19_, connection_1__9__18_,
         connection_1__9__17_, connection_1__9__16_, connection_1__9__15_,
         connection_1__9__14_, connection_1__9__13_, connection_1__9__12_,
         connection_1__9__11_, connection_1__9__10_, connection_1__9__9_,
         connection_1__9__8_, connection_1__9__7_, connection_1__9__6_,
         connection_1__9__5_, connection_1__9__4_, connection_1__9__3_,
         connection_1__9__2_, connection_1__9__1_, connection_1__9__0_,
         connection_1__10__31_, connection_1__10__30_, connection_1__10__29_,
         connection_1__10__28_, connection_1__10__27_, connection_1__10__26_,
         connection_1__10__25_, connection_1__10__24_, connection_1__10__23_,
         connection_1__10__22_, connection_1__10__21_, connection_1__10__20_,
         connection_1__10__19_, connection_1__10__18_, connection_1__10__17_,
         connection_1__10__16_, connection_1__10__15_, connection_1__10__14_,
         connection_1__10__13_, connection_1__10__12_, connection_1__10__11_,
         connection_1__10__10_, connection_1__10__9_, connection_1__10__8_,
         connection_1__10__7_, connection_1__10__6_, connection_1__10__5_,
         connection_1__10__4_, connection_1__10__3_, connection_1__10__2_,
         connection_1__10__1_, connection_1__10__0_, connection_1__11__31_,
         connection_1__11__30_, connection_1__11__29_, connection_1__11__28_,
         connection_1__11__27_, connection_1__11__26_, connection_1__11__25_,
         connection_1__11__24_, connection_1__11__23_, connection_1__11__22_,
         connection_1__11__21_, connection_1__11__20_, connection_1__11__19_,
         connection_1__11__18_, connection_1__11__17_, connection_1__11__16_,
         connection_1__11__15_, connection_1__11__14_, connection_1__11__13_,
         connection_1__11__12_, connection_1__11__11_, connection_1__11__10_,
         connection_1__11__9_, connection_1__11__8_, connection_1__11__7_,
         connection_1__11__6_, connection_1__11__5_, connection_1__11__4_,
         connection_1__11__3_, connection_1__11__2_, connection_1__11__1_,
         connection_1__11__0_, connection_1__12__31_, connection_1__12__30_,
         connection_1__12__29_, connection_1__12__28_, connection_1__12__27_,
         connection_1__12__26_, connection_1__12__25_, connection_1__12__24_,
         connection_1__12__23_, connection_1__12__22_, connection_1__12__21_,
         connection_1__12__20_, connection_1__12__19_, connection_1__12__18_,
         connection_1__12__17_, connection_1__12__16_, connection_1__12__15_,
         connection_1__12__14_, connection_1__12__13_, connection_1__12__12_,
         connection_1__12__11_, connection_1__12__10_, connection_1__12__9_,
         connection_1__12__8_, connection_1__12__7_, connection_1__12__6_,
         connection_1__12__5_, connection_1__12__4_, connection_1__12__3_,
         connection_1__12__2_, connection_1__12__1_, connection_1__12__0_,
         connection_1__13__31_, connection_1__13__30_, connection_1__13__29_,
         connection_1__13__28_, connection_1__13__27_, connection_1__13__26_,
         connection_1__13__25_, connection_1__13__24_, connection_1__13__23_,
         connection_1__13__22_, connection_1__13__21_, connection_1__13__20_,
         connection_1__13__19_, connection_1__13__18_, connection_1__13__17_,
         connection_1__13__16_, connection_1__13__15_, connection_1__13__14_,
         connection_1__13__13_, connection_1__13__12_, connection_1__13__11_,
         connection_1__13__10_, connection_1__13__9_, connection_1__13__8_,
         connection_1__13__7_, connection_1__13__6_, connection_1__13__5_,
         connection_1__13__4_, connection_1__13__3_, connection_1__13__2_,
         connection_1__13__1_, connection_1__13__0_, connection_1__14__31_,
         connection_1__14__30_, connection_1__14__29_, connection_1__14__28_,
         connection_1__14__27_, connection_1__14__26_, connection_1__14__25_,
         connection_1__14__24_, connection_1__14__23_, connection_1__14__22_,
         connection_1__14__21_, connection_1__14__20_, connection_1__14__19_,
         connection_1__14__18_, connection_1__14__17_, connection_1__14__16_,
         connection_1__14__15_, connection_1__14__14_, connection_1__14__13_,
         connection_1__14__12_, connection_1__14__11_, connection_1__14__10_,
         connection_1__14__9_, connection_1__14__8_, connection_1__14__7_,
         connection_1__14__6_, connection_1__14__5_, connection_1__14__4_,
         connection_1__14__3_, connection_1__14__2_, connection_1__14__1_,
         connection_1__14__0_, connection_1__15__31_, connection_1__15__30_,
         connection_1__15__29_, connection_1__15__28_, connection_1__15__27_,
         connection_1__15__26_, connection_1__15__25_, connection_1__15__24_,
         connection_1__15__23_, connection_1__15__22_, connection_1__15__21_,
         connection_1__15__20_, connection_1__15__19_, connection_1__15__18_,
         connection_1__15__17_, connection_1__15__16_, connection_1__15__15_,
         connection_1__15__14_, connection_1__15__13_, connection_1__15__12_,
         connection_1__15__11_, connection_1__15__10_, connection_1__15__9_,
         connection_1__15__8_, connection_1__15__7_, connection_1__15__6_,
         connection_1__15__5_, connection_1__15__4_, connection_1__15__3_,
         connection_1__15__2_, connection_1__15__1_, connection_1__15__0_,
         connection_2__0__31_, connection_2__0__30_, connection_2__0__29_,
         connection_2__0__28_, connection_2__0__27_, connection_2__0__26_,
         connection_2__0__25_, connection_2__0__24_, connection_2__0__23_,
         connection_2__0__22_, connection_2__0__21_, connection_2__0__20_,
         connection_2__0__19_, connection_2__0__18_, connection_2__0__17_,
         connection_2__0__16_, connection_2__0__15_, connection_2__0__14_,
         connection_2__0__13_, connection_2__0__12_, connection_2__0__11_,
         connection_2__0__10_, connection_2__0__9_, connection_2__0__8_,
         connection_2__0__7_, connection_2__0__6_, connection_2__0__5_,
         connection_2__0__4_, connection_2__0__3_, connection_2__0__2_,
         connection_2__0__1_, connection_2__0__0_, connection_2__1__31_,
         connection_2__1__30_, connection_2__1__29_, connection_2__1__28_,
         connection_2__1__27_, connection_2__1__26_, connection_2__1__25_,
         connection_2__1__24_, connection_2__1__23_, connection_2__1__22_,
         connection_2__1__21_, connection_2__1__20_, connection_2__1__19_,
         connection_2__1__18_, connection_2__1__17_, connection_2__1__16_,
         connection_2__1__15_, connection_2__1__14_, connection_2__1__13_,
         connection_2__1__12_, connection_2__1__11_, connection_2__1__10_,
         connection_2__1__9_, connection_2__1__8_, connection_2__1__7_,
         connection_2__1__6_, connection_2__1__5_, connection_2__1__4_,
         connection_2__1__3_, connection_2__1__2_, connection_2__1__1_,
         connection_2__1__0_, connection_2__2__31_, connection_2__2__30_,
         connection_2__2__29_, connection_2__2__28_, connection_2__2__27_,
         connection_2__2__26_, connection_2__2__25_, connection_2__2__24_,
         connection_2__2__23_, connection_2__2__22_, connection_2__2__21_,
         connection_2__2__20_, connection_2__2__19_, connection_2__2__18_,
         connection_2__2__17_, connection_2__2__16_, connection_2__2__15_,
         connection_2__2__14_, connection_2__2__13_, connection_2__2__12_,
         connection_2__2__11_, connection_2__2__10_, connection_2__2__9_,
         connection_2__2__8_, connection_2__2__7_, connection_2__2__6_,
         connection_2__2__5_, connection_2__2__4_, connection_2__2__3_,
         connection_2__2__2_, connection_2__2__1_, connection_2__2__0_,
         connection_2__3__31_, connection_2__3__30_, connection_2__3__29_,
         connection_2__3__28_, connection_2__3__27_, connection_2__3__26_,
         connection_2__3__25_, connection_2__3__24_, connection_2__3__23_,
         connection_2__3__22_, connection_2__3__21_, connection_2__3__20_,
         connection_2__3__19_, connection_2__3__18_, connection_2__3__17_,
         connection_2__3__16_, connection_2__3__15_, connection_2__3__14_,
         connection_2__3__13_, connection_2__3__12_, connection_2__3__11_,
         connection_2__3__10_, connection_2__3__9_, connection_2__3__8_,
         connection_2__3__7_, connection_2__3__6_, connection_2__3__5_,
         connection_2__3__4_, connection_2__3__3_, connection_2__3__2_,
         connection_2__3__1_, connection_2__3__0_, connection_2__4__31_,
         connection_2__4__30_, connection_2__4__29_, connection_2__4__28_,
         connection_2__4__27_, connection_2__4__26_, connection_2__4__25_,
         connection_2__4__24_, connection_2__4__23_, connection_2__4__22_,
         connection_2__4__21_, connection_2__4__20_, connection_2__4__19_,
         connection_2__4__18_, connection_2__4__17_, connection_2__4__16_,
         connection_2__4__15_, connection_2__4__14_, connection_2__4__13_,
         connection_2__4__12_, connection_2__4__11_, connection_2__4__10_,
         connection_2__4__9_, connection_2__4__8_, connection_2__4__7_,
         connection_2__4__6_, connection_2__4__5_, connection_2__4__4_,
         connection_2__4__3_, connection_2__4__2_, connection_2__4__1_,
         connection_2__4__0_, connection_2__5__31_, connection_2__5__30_,
         connection_2__5__29_, connection_2__5__28_, connection_2__5__27_,
         connection_2__5__26_, connection_2__5__25_, connection_2__5__24_,
         connection_2__5__23_, connection_2__5__22_, connection_2__5__21_,
         connection_2__5__20_, connection_2__5__19_, connection_2__5__18_,
         connection_2__5__17_, connection_2__5__16_, connection_2__5__15_,
         connection_2__5__14_, connection_2__5__13_, connection_2__5__12_,
         connection_2__5__11_, connection_2__5__10_, connection_2__5__9_,
         connection_2__5__8_, connection_2__5__7_, connection_2__5__6_,
         connection_2__5__5_, connection_2__5__4_, connection_2__5__3_,
         connection_2__5__2_, connection_2__5__1_, connection_2__5__0_,
         connection_2__6__31_, connection_2__6__30_, connection_2__6__29_,
         connection_2__6__28_, connection_2__6__27_, connection_2__6__26_,
         connection_2__6__25_, connection_2__6__24_, connection_2__6__23_,
         connection_2__6__22_, connection_2__6__21_, connection_2__6__20_,
         connection_2__6__19_, connection_2__6__18_, connection_2__6__17_,
         connection_2__6__16_, connection_2__6__15_, connection_2__6__14_,
         connection_2__6__13_, connection_2__6__12_, connection_2__6__11_,
         connection_2__6__10_, connection_2__6__9_, connection_2__6__8_,
         connection_2__6__7_, connection_2__6__6_, connection_2__6__5_,
         connection_2__6__4_, connection_2__6__3_, connection_2__6__2_,
         connection_2__6__1_, connection_2__6__0_, connection_2__7__31_,
         connection_2__7__30_, connection_2__7__29_, connection_2__7__28_,
         connection_2__7__27_, connection_2__7__26_, connection_2__7__25_,
         connection_2__7__24_, connection_2__7__23_, connection_2__7__22_,
         connection_2__7__21_, connection_2__7__20_, connection_2__7__19_,
         connection_2__7__18_, connection_2__7__17_, connection_2__7__16_,
         connection_2__7__15_, connection_2__7__14_, connection_2__7__13_,
         connection_2__7__12_, connection_2__7__11_, connection_2__7__10_,
         connection_2__7__9_, connection_2__7__8_, connection_2__7__7_,
         connection_2__7__6_, connection_2__7__5_, connection_2__7__4_,
         connection_2__7__3_, connection_2__7__2_, connection_2__7__1_,
         connection_2__7__0_, connection_2__8__31_, connection_2__8__30_,
         connection_2__8__29_, connection_2__8__28_, connection_2__8__27_,
         connection_2__8__26_, connection_2__8__25_, connection_2__8__24_,
         connection_2__8__23_, connection_2__8__22_, connection_2__8__21_,
         connection_2__8__20_, connection_2__8__19_, connection_2__8__18_,
         connection_2__8__17_, connection_2__8__16_, connection_2__8__15_,
         connection_2__8__14_, connection_2__8__13_, connection_2__8__12_,
         connection_2__8__11_, connection_2__8__10_, connection_2__8__9_,
         connection_2__8__8_, connection_2__8__7_, connection_2__8__6_,
         connection_2__8__5_, connection_2__8__4_, connection_2__8__3_,
         connection_2__8__2_, connection_2__8__1_, connection_2__8__0_,
         connection_2__9__31_, connection_2__9__30_, connection_2__9__29_,
         connection_2__9__28_, connection_2__9__27_, connection_2__9__26_,
         connection_2__9__25_, connection_2__9__24_, connection_2__9__23_,
         connection_2__9__22_, connection_2__9__21_, connection_2__9__20_,
         connection_2__9__19_, connection_2__9__18_, connection_2__9__17_,
         connection_2__9__16_, connection_2__9__15_, connection_2__9__14_,
         connection_2__9__13_, connection_2__9__12_, connection_2__9__11_,
         connection_2__9__10_, connection_2__9__9_, connection_2__9__8_,
         connection_2__9__7_, connection_2__9__6_, connection_2__9__5_,
         connection_2__9__4_, connection_2__9__3_, connection_2__9__2_,
         connection_2__9__1_, connection_2__9__0_, connection_2__10__31_,
         connection_2__10__30_, connection_2__10__29_, connection_2__10__28_,
         connection_2__10__27_, connection_2__10__26_, connection_2__10__25_,
         connection_2__10__24_, connection_2__10__23_, connection_2__10__22_,
         connection_2__10__21_, connection_2__10__20_, connection_2__10__19_,
         connection_2__10__18_, connection_2__10__17_, connection_2__10__16_,
         connection_2__10__15_, connection_2__10__14_, connection_2__10__13_,
         connection_2__10__12_, connection_2__10__11_, connection_2__10__10_,
         connection_2__10__9_, connection_2__10__8_, connection_2__10__7_,
         connection_2__10__6_, connection_2__10__5_, connection_2__10__4_,
         connection_2__10__3_, connection_2__10__2_, connection_2__10__1_,
         connection_2__10__0_, connection_2__11__31_, connection_2__11__30_,
         connection_2__11__29_, connection_2__11__28_, connection_2__11__27_,
         connection_2__11__26_, connection_2__11__25_, connection_2__11__24_,
         connection_2__11__23_, connection_2__11__22_, connection_2__11__21_,
         connection_2__11__20_, connection_2__11__19_, connection_2__11__18_,
         connection_2__11__17_, connection_2__11__16_, connection_2__11__15_,
         connection_2__11__14_, connection_2__11__13_, connection_2__11__12_,
         connection_2__11__11_, connection_2__11__10_, connection_2__11__9_,
         connection_2__11__8_, connection_2__11__7_, connection_2__11__6_,
         connection_2__11__5_, connection_2__11__4_, connection_2__11__3_,
         connection_2__11__2_, connection_2__11__1_, connection_2__11__0_,
         connection_2__12__31_, connection_2__12__30_, connection_2__12__29_,
         connection_2__12__28_, connection_2__12__27_, connection_2__12__26_,
         connection_2__12__25_, connection_2__12__24_, connection_2__12__23_,
         connection_2__12__22_, connection_2__12__21_, connection_2__12__20_,
         connection_2__12__19_, connection_2__12__18_, connection_2__12__17_,
         connection_2__12__16_, connection_2__12__15_, connection_2__12__14_,
         connection_2__12__13_, connection_2__12__12_, connection_2__12__11_,
         connection_2__12__10_, connection_2__12__9_, connection_2__12__8_,
         connection_2__12__7_, connection_2__12__6_, connection_2__12__5_,
         connection_2__12__4_, connection_2__12__3_, connection_2__12__2_,
         connection_2__12__1_, connection_2__12__0_, connection_2__13__31_,
         connection_2__13__30_, connection_2__13__29_, connection_2__13__28_,
         connection_2__13__27_, connection_2__13__26_, connection_2__13__25_,
         connection_2__13__24_, connection_2__13__23_, connection_2__13__22_,
         connection_2__13__21_, connection_2__13__20_, connection_2__13__19_,
         connection_2__13__18_, connection_2__13__17_, connection_2__13__16_,
         connection_2__13__15_, connection_2__13__14_, connection_2__13__13_,
         connection_2__13__12_, connection_2__13__11_, connection_2__13__10_,
         connection_2__13__9_, connection_2__13__8_, connection_2__13__7_,
         connection_2__13__6_, connection_2__13__5_, connection_2__13__4_,
         connection_2__13__3_, connection_2__13__2_, connection_2__13__1_,
         connection_2__13__0_, connection_2__14__31_, connection_2__14__30_,
         connection_2__14__29_, connection_2__14__28_, connection_2__14__27_,
         connection_2__14__26_, connection_2__14__25_, connection_2__14__24_,
         connection_2__14__23_, connection_2__14__22_, connection_2__14__21_,
         connection_2__14__20_, connection_2__14__19_, connection_2__14__18_,
         connection_2__14__17_, connection_2__14__16_, connection_2__14__15_,
         connection_2__14__14_, connection_2__14__13_, connection_2__14__12_,
         connection_2__14__11_, connection_2__14__10_, connection_2__14__9_,
         connection_2__14__8_, connection_2__14__7_, connection_2__14__6_,
         connection_2__14__5_, connection_2__14__4_, connection_2__14__3_,
         connection_2__14__2_, connection_2__14__1_, connection_2__14__0_,
         connection_2__15__31_, connection_2__15__30_, connection_2__15__29_,
         connection_2__15__28_, connection_2__15__27_, connection_2__15__26_,
         connection_2__15__25_, connection_2__15__24_, connection_2__15__23_,
         connection_2__15__22_, connection_2__15__21_, connection_2__15__20_,
         connection_2__15__19_, connection_2__15__18_, connection_2__15__17_,
         connection_2__15__16_, connection_2__15__15_, connection_2__15__14_,
         connection_2__15__13_, connection_2__15__12_, connection_2__15__11_,
         connection_2__15__10_, connection_2__15__9_, connection_2__15__8_,
         connection_2__15__7_, connection_2__15__6_, connection_2__15__5_,
         connection_2__15__4_, connection_2__15__3_, connection_2__15__2_,
         connection_2__15__1_, connection_2__15__0_, connection_3__0__31_,
         connection_3__0__30_, connection_3__0__29_, connection_3__0__28_,
         connection_3__0__27_, connection_3__0__26_, connection_3__0__25_,
         connection_3__0__24_, connection_3__0__23_, connection_3__0__22_,
         connection_3__0__21_, connection_3__0__20_, connection_3__0__19_,
         connection_3__0__18_, connection_3__0__17_, connection_3__0__16_,
         connection_3__0__15_, connection_3__0__14_, connection_3__0__13_,
         connection_3__0__12_, connection_3__0__11_, connection_3__0__10_,
         connection_3__0__9_, connection_3__0__8_, connection_3__0__7_,
         connection_3__0__6_, connection_3__0__5_, connection_3__0__4_,
         connection_3__0__3_, connection_3__0__2_, connection_3__0__1_,
         connection_3__0__0_, connection_3__1__31_, connection_3__1__30_,
         connection_3__1__29_, connection_3__1__28_, connection_3__1__27_,
         connection_3__1__26_, connection_3__1__25_, connection_3__1__24_,
         connection_3__1__23_, connection_3__1__22_, connection_3__1__21_,
         connection_3__1__20_, connection_3__1__19_, connection_3__1__18_,
         connection_3__1__17_, connection_3__1__16_, connection_3__1__15_,
         connection_3__1__14_, connection_3__1__13_, connection_3__1__12_,
         connection_3__1__11_, connection_3__1__10_, connection_3__1__9_,
         connection_3__1__8_, connection_3__1__7_, connection_3__1__6_,
         connection_3__1__5_, connection_3__1__4_, connection_3__1__3_,
         connection_3__1__2_, connection_3__1__1_, connection_3__1__0_,
         connection_3__2__31_, connection_3__2__30_, connection_3__2__29_,
         connection_3__2__28_, connection_3__2__27_, connection_3__2__26_,
         connection_3__2__25_, connection_3__2__24_, connection_3__2__23_,
         connection_3__2__22_, connection_3__2__21_, connection_3__2__20_,
         connection_3__2__19_, connection_3__2__18_, connection_3__2__17_,
         connection_3__2__16_, connection_3__2__15_, connection_3__2__14_,
         connection_3__2__13_, connection_3__2__12_, connection_3__2__11_,
         connection_3__2__10_, connection_3__2__9_, connection_3__2__8_,
         connection_3__2__7_, connection_3__2__6_, connection_3__2__5_,
         connection_3__2__4_, connection_3__2__3_, connection_3__2__2_,
         connection_3__2__1_, connection_3__2__0_, connection_3__3__31_,
         connection_3__3__30_, connection_3__3__29_, connection_3__3__28_,
         connection_3__3__27_, connection_3__3__26_, connection_3__3__25_,
         connection_3__3__24_, connection_3__3__23_, connection_3__3__22_,
         connection_3__3__21_, connection_3__3__20_, connection_3__3__19_,
         connection_3__3__18_, connection_3__3__17_, connection_3__3__16_,
         connection_3__3__15_, connection_3__3__14_, connection_3__3__13_,
         connection_3__3__12_, connection_3__3__11_, connection_3__3__10_,
         connection_3__3__9_, connection_3__3__8_, connection_3__3__7_,
         connection_3__3__6_, connection_3__3__5_, connection_3__3__4_,
         connection_3__3__3_, connection_3__3__2_, connection_3__3__1_,
         connection_3__3__0_, connection_3__4__31_, connection_3__4__30_,
         connection_3__4__29_, connection_3__4__28_, connection_3__4__27_,
         connection_3__4__26_, connection_3__4__25_, connection_3__4__24_,
         connection_3__4__23_, connection_3__4__22_, connection_3__4__21_,
         connection_3__4__20_, connection_3__4__19_, connection_3__4__18_,
         connection_3__4__17_, connection_3__4__16_, connection_3__4__15_,
         connection_3__4__14_, connection_3__4__13_, connection_3__4__12_,
         connection_3__4__11_, connection_3__4__10_, connection_3__4__9_,
         connection_3__4__8_, connection_3__4__7_, connection_3__4__6_,
         connection_3__4__5_, connection_3__4__4_, connection_3__4__3_,
         connection_3__4__2_, connection_3__4__1_, connection_3__4__0_,
         connection_3__5__31_, connection_3__5__30_, connection_3__5__29_,
         connection_3__5__28_, connection_3__5__27_, connection_3__5__26_,
         connection_3__5__25_, connection_3__5__24_, connection_3__5__23_,
         connection_3__5__22_, connection_3__5__21_, connection_3__5__20_,
         connection_3__5__19_, connection_3__5__18_, connection_3__5__17_,
         connection_3__5__16_, connection_3__5__15_, connection_3__5__14_,
         connection_3__5__13_, connection_3__5__12_, connection_3__5__11_,
         connection_3__5__10_, connection_3__5__9_, connection_3__5__8_,
         connection_3__5__7_, connection_3__5__6_, connection_3__5__5_,
         connection_3__5__4_, connection_3__5__3_, connection_3__5__2_,
         connection_3__5__1_, connection_3__5__0_, connection_3__6__31_,
         connection_3__6__30_, connection_3__6__29_, connection_3__6__28_,
         connection_3__6__27_, connection_3__6__26_, connection_3__6__25_,
         connection_3__6__24_, connection_3__6__23_, connection_3__6__22_,
         connection_3__6__21_, connection_3__6__20_, connection_3__6__19_,
         connection_3__6__18_, connection_3__6__17_, connection_3__6__16_,
         connection_3__6__15_, connection_3__6__14_, connection_3__6__13_,
         connection_3__6__12_, connection_3__6__11_, connection_3__6__10_,
         connection_3__6__9_, connection_3__6__8_, connection_3__6__7_,
         connection_3__6__6_, connection_3__6__5_, connection_3__6__4_,
         connection_3__6__3_, connection_3__6__2_, connection_3__6__1_,
         connection_3__6__0_, connection_3__7__31_, connection_3__7__30_,
         connection_3__7__29_, connection_3__7__28_, connection_3__7__27_,
         connection_3__7__26_, connection_3__7__25_, connection_3__7__24_,
         connection_3__7__23_, connection_3__7__22_, connection_3__7__21_,
         connection_3__7__20_, connection_3__7__19_, connection_3__7__18_,
         connection_3__7__17_, connection_3__7__16_, connection_3__7__15_,
         connection_3__7__14_, connection_3__7__13_, connection_3__7__12_,
         connection_3__7__11_, connection_3__7__10_, connection_3__7__9_,
         connection_3__7__8_, connection_3__7__7_, connection_3__7__6_,
         connection_3__7__5_, connection_3__7__4_, connection_3__7__3_,
         connection_3__7__2_, connection_3__7__1_, connection_3__7__0_,
         connection_3__8__31_, connection_3__8__30_, connection_3__8__29_,
         connection_3__8__28_, connection_3__8__27_, connection_3__8__26_,
         connection_3__8__25_, connection_3__8__24_, connection_3__8__23_,
         connection_3__8__22_, connection_3__8__21_, connection_3__8__20_,
         connection_3__8__19_, connection_3__8__18_, connection_3__8__17_,
         connection_3__8__16_, connection_3__8__15_, connection_3__8__14_,
         connection_3__8__13_, connection_3__8__12_, connection_3__8__11_,
         connection_3__8__10_, connection_3__8__9_, connection_3__8__8_,
         connection_3__8__7_, connection_3__8__6_, connection_3__8__5_,
         connection_3__8__4_, connection_3__8__3_, connection_3__8__2_,
         connection_3__8__1_, connection_3__8__0_, connection_3__9__31_,
         connection_3__9__30_, connection_3__9__29_, connection_3__9__28_,
         connection_3__9__27_, connection_3__9__26_, connection_3__9__25_,
         connection_3__9__24_, connection_3__9__23_, connection_3__9__22_,
         connection_3__9__21_, connection_3__9__20_, connection_3__9__19_,
         connection_3__9__18_, connection_3__9__17_, connection_3__9__16_,
         connection_3__9__15_, connection_3__9__14_, connection_3__9__13_,
         connection_3__9__12_, connection_3__9__11_, connection_3__9__10_,
         connection_3__9__9_, connection_3__9__8_, connection_3__9__7_,
         connection_3__9__6_, connection_3__9__5_, connection_3__9__4_,
         connection_3__9__3_, connection_3__9__2_, connection_3__9__1_,
         connection_3__9__0_, connection_3__10__31_, connection_3__10__30_,
         connection_3__10__29_, connection_3__10__28_, connection_3__10__27_,
         connection_3__10__26_, connection_3__10__25_, connection_3__10__24_,
         connection_3__10__23_, connection_3__10__22_, connection_3__10__21_,
         connection_3__10__20_, connection_3__10__19_, connection_3__10__18_,
         connection_3__10__17_, connection_3__10__16_, connection_3__10__15_,
         connection_3__10__14_, connection_3__10__13_, connection_3__10__12_,
         connection_3__10__11_, connection_3__10__10_, connection_3__10__9_,
         connection_3__10__8_, connection_3__10__7_, connection_3__10__6_,
         connection_3__10__5_, connection_3__10__4_, connection_3__10__3_,
         connection_3__10__2_, connection_3__10__1_, connection_3__10__0_,
         connection_3__11__31_, connection_3__11__30_, connection_3__11__29_,
         connection_3__11__28_, connection_3__11__27_, connection_3__11__26_,
         connection_3__11__25_, connection_3__11__24_, connection_3__11__23_,
         connection_3__11__22_, connection_3__11__21_, connection_3__11__20_,
         connection_3__11__19_, connection_3__11__18_, connection_3__11__17_,
         connection_3__11__16_, connection_3__11__15_, connection_3__11__14_,
         connection_3__11__13_, connection_3__11__12_, connection_3__11__11_,
         connection_3__11__10_, connection_3__11__9_, connection_3__11__8_,
         connection_3__11__7_, connection_3__11__6_, connection_3__11__5_,
         connection_3__11__4_, connection_3__11__3_, connection_3__11__2_,
         connection_3__11__1_, connection_3__11__0_, connection_3__12__31_,
         connection_3__12__30_, connection_3__12__29_, connection_3__12__28_,
         connection_3__12__27_, connection_3__12__26_, connection_3__12__25_,
         connection_3__12__24_, connection_3__12__23_, connection_3__12__22_,
         connection_3__12__21_, connection_3__12__20_, connection_3__12__19_,
         connection_3__12__18_, connection_3__12__17_, connection_3__12__16_,
         connection_3__12__15_, connection_3__12__14_, connection_3__12__13_,
         connection_3__12__12_, connection_3__12__11_, connection_3__12__10_,
         connection_3__12__9_, connection_3__12__8_, connection_3__12__7_,
         connection_3__12__6_, connection_3__12__5_, connection_3__12__4_,
         connection_3__12__3_, connection_3__12__2_, connection_3__12__1_,
         connection_3__12__0_, connection_3__13__31_, connection_3__13__30_,
         connection_3__13__29_, connection_3__13__28_, connection_3__13__27_,
         connection_3__13__26_, connection_3__13__25_, connection_3__13__24_,
         connection_3__13__23_, connection_3__13__22_, connection_3__13__21_,
         connection_3__13__20_, connection_3__13__19_, connection_3__13__18_,
         connection_3__13__17_, connection_3__13__16_, connection_3__13__15_,
         connection_3__13__14_, connection_3__13__13_, connection_3__13__12_,
         connection_3__13__11_, connection_3__13__10_, connection_3__13__9_,
         connection_3__13__8_, connection_3__13__7_, connection_3__13__6_,
         connection_3__13__5_, connection_3__13__4_, connection_3__13__3_,
         connection_3__13__2_, connection_3__13__1_, connection_3__13__0_,
         connection_3__14__31_, connection_3__14__30_, connection_3__14__29_,
         connection_3__14__28_, connection_3__14__27_, connection_3__14__26_,
         connection_3__14__25_, connection_3__14__24_, connection_3__14__23_,
         connection_3__14__22_, connection_3__14__21_, connection_3__14__20_,
         connection_3__14__19_, connection_3__14__18_, connection_3__14__17_,
         connection_3__14__16_, connection_3__14__15_, connection_3__14__14_,
         connection_3__14__13_, connection_3__14__12_, connection_3__14__11_,
         connection_3__14__10_, connection_3__14__9_, connection_3__14__8_,
         connection_3__14__7_, connection_3__14__6_, connection_3__14__5_,
         connection_3__14__4_, connection_3__14__3_, connection_3__14__2_,
         connection_3__14__1_, connection_3__14__0_, connection_3__15__31_,
         connection_3__15__30_, connection_3__15__29_, connection_3__15__28_,
         connection_3__15__27_, connection_3__15__26_, connection_3__15__25_,
         connection_3__15__24_, connection_3__15__23_, connection_3__15__22_,
         connection_3__15__21_, connection_3__15__20_, connection_3__15__19_,
         connection_3__15__18_, connection_3__15__17_, connection_3__15__16_,
         connection_3__15__15_, connection_3__15__14_, connection_3__15__13_,
         connection_3__15__12_, connection_3__15__11_, connection_3__15__10_,
         connection_3__15__9_, connection_3__15__8_, connection_3__15__7_,
         connection_3__15__6_, connection_3__15__5_, connection_3__15__4_,
         connection_3__15__3_, connection_3__15__2_, connection_3__15__1_,
         connection_3__15__0_, connection_4__0__31_, connection_4__0__30_,
         connection_4__0__29_, connection_4__0__28_, connection_4__0__27_,
         connection_4__0__26_, connection_4__0__25_, connection_4__0__24_,
         connection_4__0__23_, connection_4__0__22_, connection_4__0__21_,
         connection_4__0__20_, connection_4__0__19_, connection_4__0__18_,
         connection_4__0__17_, connection_4__0__16_, connection_4__0__15_,
         connection_4__0__14_, connection_4__0__13_, connection_4__0__12_,
         connection_4__0__11_, connection_4__0__10_, connection_4__0__9_,
         connection_4__0__8_, connection_4__0__7_, connection_4__0__6_,
         connection_4__0__5_, connection_4__0__4_, connection_4__0__3_,
         connection_4__0__2_, connection_4__0__1_, connection_4__0__0_,
         connection_4__1__31_, connection_4__1__30_, connection_4__1__29_,
         connection_4__1__28_, connection_4__1__27_, connection_4__1__26_,
         connection_4__1__25_, connection_4__1__24_, connection_4__1__23_,
         connection_4__1__22_, connection_4__1__21_, connection_4__1__20_,
         connection_4__1__19_, connection_4__1__18_, connection_4__1__17_,
         connection_4__1__16_, connection_4__1__15_, connection_4__1__14_,
         connection_4__1__13_, connection_4__1__12_, connection_4__1__11_,
         connection_4__1__10_, connection_4__1__9_, connection_4__1__8_,
         connection_4__1__7_, connection_4__1__6_, connection_4__1__5_,
         connection_4__1__4_, connection_4__1__3_, connection_4__1__2_,
         connection_4__1__1_, connection_4__1__0_, connection_4__2__31_,
         connection_4__2__30_, connection_4__2__29_, connection_4__2__28_,
         connection_4__2__27_, connection_4__2__26_, connection_4__2__25_,
         connection_4__2__24_, connection_4__2__23_, connection_4__2__22_,
         connection_4__2__21_, connection_4__2__20_, connection_4__2__19_,
         connection_4__2__18_, connection_4__2__17_, connection_4__2__16_,
         connection_4__2__15_, connection_4__2__14_, connection_4__2__13_,
         connection_4__2__12_, connection_4__2__11_, connection_4__2__10_,
         connection_4__2__9_, connection_4__2__8_, connection_4__2__7_,
         connection_4__2__6_, connection_4__2__5_, connection_4__2__4_,
         connection_4__2__3_, connection_4__2__2_, connection_4__2__1_,
         connection_4__2__0_, connection_4__3__31_, connection_4__3__30_,
         connection_4__3__29_, connection_4__3__28_, connection_4__3__27_,
         connection_4__3__26_, connection_4__3__25_, connection_4__3__24_,
         connection_4__3__23_, connection_4__3__22_, connection_4__3__21_,
         connection_4__3__20_, connection_4__3__19_, connection_4__3__18_,
         connection_4__3__17_, connection_4__3__16_, connection_4__3__15_,
         connection_4__3__14_, connection_4__3__13_, connection_4__3__12_,
         connection_4__3__11_, connection_4__3__10_, connection_4__3__9_,
         connection_4__3__8_, connection_4__3__7_, connection_4__3__6_,
         connection_4__3__5_, connection_4__3__4_, connection_4__3__3_,
         connection_4__3__2_, connection_4__3__1_, connection_4__3__0_,
         connection_4__4__31_, connection_4__4__30_, connection_4__4__29_,
         connection_4__4__28_, connection_4__4__27_, connection_4__4__26_,
         connection_4__4__25_, connection_4__4__24_, connection_4__4__23_,
         connection_4__4__22_, connection_4__4__21_, connection_4__4__20_,
         connection_4__4__19_, connection_4__4__18_, connection_4__4__17_,
         connection_4__4__16_, connection_4__4__15_, connection_4__4__14_,
         connection_4__4__13_, connection_4__4__12_, connection_4__4__11_,
         connection_4__4__10_, connection_4__4__9_, connection_4__4__8_,
         connection_4__4__7_, connection_4__4__6_, connection_4__4__5_,
         connection_4__4__4_, connection_4__4__3_, connection_4__4__2_,
         connection_4__4__1_, connection_4__4__0_, connection_4__5__31_,
         connection_4__5__30_, connection_4__5__29_, connection_4__5__28_,
         connection_4__5__27_, connection_4__5__26_, connection_4__5__25_,
         connection_4__5__24_, connection_4__5__23_, connection_4__5__22_,
         connection_4__5__21_, connection_4__5__20_, connection_4__5__19_,
         connection_4__5__18_, connection_4__5__17_, connection_4__5__16_,
         connection_4__5__15_, connection_4__5__14_, connection_4__5__13_,
         connection_4__5__12_, connection_4__5__11_, connection_4__5__10_,
         connection_4__5__9_, connection_4__5__8_, connection_4__5__7_,
         connection_4__5__6_, connection_4__5__5_, connection_4__5__4_,
         connection_4__5__3_, connection_4__5__2_, connection_4__5__1_,
         connection_4__5__0_, connection_4__6__31_, connection_4__6__30_,
         connection_4__6__29_, connection_4__6__28_, connection_4__6__27_,
         connection_4__6__26_, connection_4__6__25_, connection_4__6__24_,
         connection_4__6__23_, connection_4__6__22_, connection_4__6__21_,
         connection_4__6__20_, connection_4__6__19_, connection_4__6__18_,
         connection_4__6__17_, connection_4__6__16_, connection_4__6__15_,
         connection_4__6__14_, connection_4__6__13_, connection_4__6__12_,
         connection_4__6__11_, connection_4__6__10_, connection_4__6__9_,
         connection_4__6__8_, connection_4__6__7_, connection_4__6__6_,
         connection_4__6__5_, connection_4__6__4_, connection_4__6__3_,
         connection_4__6__2_, connection_4__6__1_, connection_4__6__0_,
         connection_4__7__31_, connection_4__7__30_, connection_4__7__29_,
         connection_4__7__28_, connection_4__7__27_, connection_4__7__26_,
         connection_4__7__25_, connection_4__7__24_, connection_4__7__23_,
         connection_4__7__22_, connection_4__7__21_, connection_4__7__20_,
         connection_4__7__19_, connection_4__7__18_, connection_4__7__17_,
         connection_4__7__16_, connection_4__7__15_, connection_4__7__14_,
         connection_4__7__13_, connection_4__7__12_, connection_4__7__11_,
         connection_4__7__10_, connection_4__7__9_, connection_4__7__8_,
         connection_4__7__7_, connection_4__7__6_, connection_4__7__5_,
         connection_4__7__4_, connection_4__7__3_, connection_4__7__2_,
         connection_4__7__1_, connection_4__7__0_, connection_4__8__31_,
         connection_4__8__30_, connection_4__8__29_, connection_4__8__28_,
         connection_4__8__27_, connection_4__8__26_, connection_4__8__25_,
         connection_4__8__24_, connection_4__8__23_, connection_4__8__22_,
         connection_4__8__21_, connection_4__8__20_, connection_4__8__19_,
         connection_4__8__18_, connection_4__8__17_, connection_4__8__16_,
         connection_4__8__15_, connection_4__8__14_, connection_4__8__13_,
         connection_4__8__12_, connection_4__8__11_, connection_4__8__10_,
         connection_4__8__9_, connection_4__8__8_, connection_4__8__7_,
         connection_4__8__6_, connection_4__8__5_, connection_4__8__4_,
         connection_4__8__3_, connection_4__8__2_, connection_4__8__1_,
         connection_4__8__0_, connection_4__9__31_, connection_4__9__30_,
         connection_4__9__29_, connection_4__9__28_, connection_4__9__27_,
         connection_4__9__26_, connection_4__9__25_, connection_4__9__24_,
         connection_4__9__23_, connection_4__9__22_, connection_4__9__21_,
         connection_4__9__20_, connection_4__9__19_, connection_4__9__18_,
         connection_4__9__17_, connection_4__9__16_, connection_4__9__15_,
         connection_4__9__14_, connection_4__9__13_, connection_4__9__12_,
         connection_4__9__11_, connection_4__9__10_, connection_4__9__9_,
         connection_4__9__8_, connection_4__9__7_, connection_4__9__6_,
         connection_4__9__5_, connection_4__9__4_, connection_4__9__3_,
         connection_4__9__2_, connection_4__9__1_, connection_4__9__0_,
         connection_4__10__31_, connection_4__10__30_, connection_4__10__29_,
         connection_4__10__28_, connection_4__10__27_, connection_4__10__26_,
         connection_4__10__25_, connection_4__10__24_, connection_4__10__23_,
         connection_4__10__22_, connection_4__10__21_, connection_4__10__20_,
         connection_4__10__19_, connection_4__10__18_, connection_4__10__17_,
         connection_4__10__16_, connection_4__10__15_, connection_4__10__14_,
         connection_4__10__13_, connection_4__10__12_, connection_4__10__11_,
         connection_4__10__10_, connection_4__10__9_, connection_4__10__8_,
         connection_4__10__7_, connection_4__10__6_, connection_4__10__5_,
         connection_4__10__4_, connection_4__10__3_, connection_4__10__2_,
         connection_4__10__1_, connection_4__10__0_, connection_4__11__31_,
         connection_4__11__30_, connection_4__11__29_, connection_4__11__28_,
         connection_4__11__27_, connection_4__11__26_, connection_4__11__25_,
         connection_4__11__24_, connection_4__11__23_, connection_4__11__22_,
         connection_4__11__21_, connection_4__11__20_, connection_4__11__19_,
         connection_4__11__18_, connection_4__11__17_, connection_4__11__16_,
         connection_4__11__15_, connection_4__11__14_, connection_4__11__13_,
         connection_4__11__12_, connection_4__11__11_, connection_4__11__10_,
         connection_4__11__9_, connection_4__11__8_, connection_4__11__7_,
         connection_4__11__6_, connection_4__11__5_, connection_4__11__4_,
         connection_4__11__3_, connection_4__11__2_, connection_4__11__1_,
         connection_4__11__0_, connection_4__12__31_, connection_4__12__30_,
         connection_4__12__29_, connection_4__12__28_, connection_4__12__27_,
         connection_4__12__26_, connection_4__12__25_, connection_4__12__24_,
         connection_4__12__23_, connection_4__12__22_, connection_4__12__21_,
         connection_4__12__20_, connection_4__12__19_, connection_4__12__18_,
         connection_4__12__17_, connection_4__12__16_, connection_4__12__15_,
         connection_4__12__14_, connection_4__12__13_, connection_4__12__12_,
         connection_4__12__11_, connection_4__12__10_, connection_4__12__9_,
         connection_4__12__8_, connection_4__12__7_, connection_4__12__6_,
         connection_4__12__5_, connection_4__12__4_, connection_4__12__3_,
         connection_4__12__2_, connection_4__12__1_, connection_4__12__0_,
         connection_4__13__31_, connection_4__13__30_, connection_4__13__29_,
         connection_4__13__28_, connection_4__13__27_, connection_4__13__26_,
         connection_4__13__25_, connection_4__13__24_, connection_4__13__23_,
         connection_4__13__22_, connection_4__13__21_, connection_4__13__20_,
         connection_4__13__19_, connection_4__13__18_, connection_4__13__17_,
         connection_4__13__16_, connection_4__13__15_, connection_4__13__14_,
         connection_4__13__13_, connection_4__13__12_, connection_4__13__11_,
         connection_4__13__10_, connection_4__13__9_, connection_4__13__8_,
         connection_4__13__7_, connection_4__13__6_, connection_4__13__5_,
         connection_4__13__4_, connection_4__13__3_, connection_4__13__2_,
         connection_4__13__1_, connection_4__13__0_, connection_4__14__31_,
         connection_4__14__30_, connection_4__14__29_, connection_4__14__28_,
         connection_4__14__27_, connection_4__14__26_, connection_4__14__25_,
         connection_4__14__24_, connection_4__14__23_, connection_4__14__22_,
         connection_4__14__21_, connection_4__14__20_, connection_4__14__19_,
         connection_4__14__18_, connection_4__14__17_, connection_4__14__16_,
         connection_4__14__15_, connection_4__14__14_, connection_4__14__13_,
         connection_4__14__12_, connection_4__14__11_, connection_4__14__10_,
         connection_4__14__9_, connection_4__14__8_, connection_4__14__7_,
         connection_4__14__6_, connection_4__14__5_, connection_4__14__4_,
         connection_4__14__3_, connection_4__14__2_, connection_4__14__1_,
         connection_4__14__0_, connection_4__15__31_, connection_4__15__30_,
         connection_4__15__29_, connection_4__15__28_, connection_4__15__27_,
         connection_4__15__26_, connection_4__15__25_, connection_4__15__24_,
         connection_4__15__23_, connection_4__15__22_, connection_4__15__21_,
         connection_4__15__20_, connection_4__15__19_, connection_4__15__18_,
         connection_4__15__17_, connection_4__15__16_, connection_4__15__15_,
         connection_4__15__14_, connection_4__15__13_, connection_4__15__12_,
         connection_4__15__11_, connection_4__15__10_, connection_4__15__9_,
         connection_4__15__8_, connection_4__15__7_, connection_4__15__6_,
         connection_4__15__5_, connection_4__15__4_, connection_4__15__3_,
         connection_4__15__2_, connection_4__15__1_, connection_4__15__0_,
         connection_5__0__31_, connection_5__0__30_, connection_5__0__29_,
         connection_5__0__28_, connection_5__0__27_, connection_5__0__26_,
         connection_5__0__25_, connection_5__0__24_, connection_5__0__23_,
         connection_5__0__22_, connection_5__0__21_, connection_5__0__20_,
         connection_5__0__19_, connection_5__0__18_, connection_5__0__17_,
         connection_5__0__16_, connection_5__0__15_, connection_5__0__14_,
         connection_5__0__13_, connection_5__0__12_, connection_5__0__11_,
         connection_5__0__10_, connection_5__0__9_, connection_5__0__8_,
         connection_5__0__7_, connection_5__0__6_, connection_5__0__5_,
         connection_5__0__4_, connection_5__0__3_, connection_5__0__2_,
         connection_5__0__1_, connection_5__0__0_, connection_5__1__31_,
         connection_5__1__30_, connection_5__1__29_, connection_5__1__28_,
         connection_5__1__27_, connection_5__1__26_, connection_5__1__25_,
         connection_5__1__24_, connection_5__1__23_, connection_5__1__22_,
         connection_5__1__21_, connection_5__1__20_, connection_5__1__19_,
         connection_5__1__18_, connection_5__1__17_, connection_5__1__16_,
         connection_5__1__15_, connection_5__1__14_, connection_5__1__13_,
         connection_5__1__12_, connection_5__1__11_, connection_5__1__10_,
         connection_5__1__9_, connection_5__1__8_, connection_5__1__7_,
         connection_5__1__6_, connection_5__1__5_, connection_5__1__4_,
         connection_5__1__3_, connection_5__1__2_, connection_5__1__1_,
         connection_5__1__0_, connection_5__2__31_, connection_5__2__30_,
         connection_5__2__29_, connection_5__2__28_, connection_5__2__27_,
         connection_5__2__26_, connection_5__2__25_, connection_5__2__24_,
         connection_5__2__23_, connection_5__2__22_, connection_5__2__21_,
         connection_5__2__20_, connection_5__2__19_, connection_5__2__18_,
         connection_5__2__17_, connection_5__2__16_, connection_5__2__15_,
         connection_5__2__14_, connection_5__2__13_, connection_5__2__12_,
         connection_5__2__11_, connection_5__2__10_, connection_5__2__9_,
         connection_5__2__8_, connection_5__2__7_, connection_5__2__6_,
         connection_5__2__5_, connection_5__2__4_, connection_5__2__3_,
         connection_5__2__2_, connection_5__2__1_, connection_5__2__0_,
         connection_5__3__31_, connection_5__3__30_, connection_5__3__29_,
         connection_5__3__28_, connection_5__3__27_, connection_5__3__26_,
         connection_5__3__25_, connection_5__3__24_, connection_5__3__23_,
         connection_5__3__22_, connection_5__3__21_, connection_5__3__20_,
         connection_5__3__19_, connection_5__3__18_, connection_5__3__17_,
         connection_5__3__16_, connection_5__3__15_, connection_5__3__14_,
         connection_5__3__13_, connection_5__3__12_, connection_5__3__11_,
         connection_5__3__10_, connection_5__3__9_, connection_5__3__8_,
         connection_5__3__7_, connection_5__3__6_, connection_5__3__5_,
         connection_5__3__4_, connection_5__3__3_, connection_5__3__2_,
         connection_5__3__1_, connection_5__3__0_, connection_5__4__31_,
         connection_5__4__30_, connection_5__4__29_, connection_5__4__28_,
         connection_5__4__27_, connection_5__4__26_, connection_5__4__25_,
         connection_5__4__24_, connection_5__4__23_, connection_5__4__22_,
         connection_5__4__21_, connection_5__4__20_, connection_5__4__19_,
         connection_5__4__18_, connection_5__4__17_, connection_5__4__16_,
         connection_5__4__15_, connection_5__4__14_, connection_5__4__13_,
         connection_5__4__12_, connection_5__4__11_, connection_5__4__10_,
         connection_5__4__9_, connection_5__4__8_, connection_5__4__7_,
         connection_5__4__6_, connection_5__4__5_, connection_5__4__4_,
         connection_5__4__3_, connection_5__4__2_, connection_5__4__1_,
         connection_5__4__0_, connection_5__5__31_, connection_5__5__30_,
         connection_5__5__29_, connection_5__5__28_, connection_5__5__27_,
         connection_5__5__26_, connection_5__5__25_, connection_5__5__24_,
         connection_5__5__23_, connection_5__5__22_, connection_5__5__21_,
         connection_5__5__20_, connection_5__5__19_, connection_5__5__18_,
         connection_5__5__17_, connection_5__5__16_, connection_5__5__15_,
         connection_5__5__14_, connection_5__5__13_, connection_5__5__12_,
         connection_5__5__11_, connection_5__5__10_, connection_5__5__9_,
         connection_5__5__8_, connection_5__5__7_, connection_5__5__6_,
         connection_5__5__5_, connection_5__5__4_, connection_5__5__3_,
         connection_5__5__2_, connection_5__5__1_, connection_5__5__0_,
         connection_5__6__31_, connection_5__6__30_, connection_5__6__29_,
         connection_5__6__28_, connection_5__6__27_, connection_5__6__26_,
         connection_5__6__25_, connection_5__6__24_, connection_5__6__23_,
         connection_5__6__22_, connection_5__6__21_, connection_5__6__20_,
         connection_5__6__19_, connection_5__6__18_, connection_5__6__17_,
         connection_5__6__16_, connection_5__6__15_, connection_5__6__14_,
         connection_5__6__13_, connection_5__6__12_, connection_5__6__11_,
         connection_5__6__10_, connection_5__6__9_, connection_5__6__8_,
         connection_5__6__7_, connection_5__6__6_, connection_5__6__5_,
         connection_5__6__4_, connection_5__6__3_, connection_5__6__2_,
         connection_5__6__1_, connection_5__6__0_, connection_5__7__31_,
         connection_5__7__30_, connection_5__7__29_, connection_5__7__28_,
         connection_5__7__27_, connection_5__7__26_, connection_5__7__25_,
         connection_5__7__24_, connection_5__7__23_, connection_5__7__22_,
         connection_5__7__21_, connection_5__7__20_, connection_5__7__19_,
         connection_5__7__18_, connection_5__7__17_, connection_5__7__16_,
         connection_5__7__15_, connection_5__7__14_, connection_5__7__13_,
         connection_5__7__12_, connection_5__7__11_, connection_5__7__10_,
         connection_5__7__9_, connection_5__7__8_, connection_5__7__7_,
         connection_5__7__6_, connection_5__7__5_, connection_5__7__4_,
         connection_5__7__3_, connection_5__7__2_, connection_5__7__1_,
         connection_5__7__0_, connection_5__8__31_, connection_5__8__30_,
         connection_5__8__29_, connection_5__8__28_, connection_5__8__27_,
         connection_5__8__26_, connection_5__8__25_, connection_5__8__24_,
         connection_5__8__23_, connection_5__8__22_, connection_5__8__21_,
         connection_5__8__20_, connection_5__8__19_, connection_5__8__18_,
         connection_5__8__17_, connection_5__8__16_, connection_5__8__15_,
         connection_5__8__14_, connection_5__8__13_, connection_5__8__12_,
         connection_5__8__11_, connection_5__8__10_, connection_5__8__9_,
         connection_5__8__8_, connection_5__8__7_, connection_5__8__6_,
         connection_5__8__5_, connection_5__8__4_, connection_5__8__3_,
         connection_5__8__2_, connection_5__8__1_, connection_5__8__0_,
         connection_5__9__31_, connection_5__9__30_, connection_5__9__29_,
         connection_5__9__28_, connection_5__9__27_, connection_5__9__26_,
         connection_5__9__25_, connection_5__9__24_, connection_5__9__23_,
         connection_5__9__22_, connection_5__9__21_, connection_5__9__20_,
         connection_5__9__19_, connection_5__9__18_, connection_5__9__17_,
         connection_5__9__16_, connection_5__9__15_, connection_5__9__14_,
         connection_5__9__13_, connection_5__9__12_, connection_5__9__11_,
         connection_5__9__10_, connection_5__9__9_, connection_5__9__8_,
         connection_5__9__7_, connection_5__9__6_, connection_5__9__5_,
         connection_5__9__4_, connection_5__9__3_, connection_5__9__2_,
         connection_5__9__1_, connection_5__9__0_, connection_5__10__31_,
         connection_5__10__30_, connection_5__10__29_, connection_5__10__28_,
         connection_5__10__27_, connection_5__10__26_, connection_5__10__25_,
         connection_5__10__24_, connection_5__10__23_, connection_5__10__22_,
         connection_5__10__21_, connection_5__10__20_, connection_5__10__19_,
         connection_5__10__18_, connection_5__10__17_, connection_5__10__16_,
         connection_5__10__15_, connection_5__10__14_, connection_5__10__13_,
         connection_5__10__12_, connection_5__10__11_, connection_5__10__10_,
         connection_5__10__9_, connection_5__10__8_, connection_5__10__7_,
         connection_5__10__6_, connection_5__10__5_, connection_5__10__4_,
         connection_5__10__3_, connection_5__10__2_, connection_5__10__1_,
         connection_5__10__0_, connection_5__11__31_, connection_5__11__30_,
         connection_5__11__29_, connection_5__11__28_, connection_5__11__27_,
         connection_5__11__26_, connection_5__11__25_, connection_5__11__24_,
         connection_5__11__23_, connection_5__11__22_, connection_5__11__21_,
         connection_5__11__20_, connection_5__11__19_, connection_5__11__18_,
         connection_5__11__17_, connection_5__11__16_, connection_5__11__15_,
         connection_5__11__14_, connection_5__11__13_, connection_5__11__12_,
         connection_5__11__11_, connection_5__11__10_, connection_5__11__9_,
         connection_5__11__8_, connection_5__11__7_, connection_5__11__6_,
         connection_5__11__5_, connection_5__11__4_, connection_5__11__3_,
         connection_5__11__2_, connection_5__11__1_, connection_5__11__0_,
         connection_5__12__31_, connection_5__12__30_, connection_5__12__29_,
         connection_5__12__28_, connection_5__12__27_, connection_5__12__26_,
         connection_5__12__25_, connection_5__12__24_, connection_5__12__23_,
         connection_5__12__22_, connection_5__12__21_, connection_5__12__20_,
         connection_5__12__19_, connection_5__12__18_, connection_5__12__17_,
         connection_5__12__16_, connection_5__12__15_, connection_5__12__14_,
         connection_5__12__13_, connection_5__12__12_, connection_5__12__11_,
         connection_5__12__10_, connection_5__12__9_, connection_5__12__8_,
         connection_5__12__7_, connection_5__12__6_, connection_5__12__5_,
         connection_5__12__4_, connection_5__12__3_, connection_5__12__2_,
         connection_5__12__1_, connection_5__12__0_, connection_5__13__31_,
         connection_5__13__30_, connection_5__13__29_, connection_5__13__28_,
         connection_5__13__27_, connection_5__13__26_, connection_5__13__25_,
         connection_5__13__24_, connection_5__13__23_, connection_5__13__22_,
         connection_5__13__21_, connection_5__13__20_, connection_5__13__19_,
         connection_5__13__18_, connection_5__13__17_, connection_5__13__16_,
         connection_5__13__15_, connection_5__13__14_, connection_5__13__13_,
         connection_5__13__12_, connection_5__13__11_, connection_5__13__10_,
         connection_5__13__9_, connection_5__13__8_, connection_5__13__7_,
         connection_5__13__6_, connection_5__13__5_, connection_5__13__4_,
         connection_5__13__3_, connection_5__13__2_, connection_5__13__1_,
         connection_5__13__0_, connection_5__14__31_, connection_5__14__30_,
         connection_5__14__29_, connection_5__14__28_, connection_5__14__27_,
         connection_5__14__26_, connection_5__14__25_, connection_5__14__24_,
         connection_5__14__23_, connection_5__14__22_, connection_5__14__21_,
         connection_5__14__20_, connection_5__14__19_, connection_5__14__18_,
         connection_5__14__17_, connection_5__14__16_, connection_5__14__15_,
         connection_5__14__14_, connection_5__14__13_, connection_5__14__12_,
         connection_5__14__11_, connection_5__14__10_, connection_5__14__9_,
         connection_5__14__8_, connection_5__14__7_, connection_5__14__6_,
         connection_5__14__5_, connection_5__14__4_, connection_5__14__3_,
         connection_5__14__2_, connection_5__14__1_, connection_5__14__0_,
         connection_5__15__31_, connection_5__15__30_, connection_5__15__29_,
         connection_5__15__28_, connection_5__15__27_, connection_5__15__26_,
         connection_5__15__25_, connection_5__15__24_, connection_5__15__23_,
         connection_5__15__22_, connection_5__15__21_, connection_5__15__20_,
         connection_5__15__19_, connection_5__15__18_, connection_5__15__17_,
         connection_5__15__16_, connection_5__15__15_, connection_5__15__14_,
         connection_5__15__13_, connection_5__15__12_, connection_5__15__11_,
         connection_5__15__10_, connection_5__15__9_, connection_5__15__8_,
         connection_5__15__7_, connection_5__15__6_, connection_5__15__5_,
         connection_5__15__4_, connection_5__15__3_, connection_5__15__2_,
         connection_5__15__1_, connection_5__15__0_, n531, n532, n533, n534;
  wire   [119:0] cmd_pipeline_stage_3__pipeline_i_cmd_reg;
  wire   [79:0] cmd_pipeline_stage_4__pipeline_i_cmd_reg;
  wire   [39:0] cmd_pipeline_stage_5__pipeline_i_cmd_reg;
  wire   [767:0] fwd_connection_frist_half;
  wire   [23:0] fwd_connection_valid_frist_half;
  wire   [767:0] fwd_connection_sec_half;
  wire   [23:0] fwd_connection_valid_sec_half;

  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_0 first_half_stages_0__sw_group_0__upper_group_0__genblk1_upper_sw_first_stage ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[1:0]), .i_data_bus(
        i_data_bus[63:0]), .o_valid({connection_valid_0__1_, 
        connection_valid_0__0_}), .o_data_bus({connection_0__1__31_, 
        connection_0__1__30_, connection_0__1__29_, connection_0__1__28_, 
        connection_0__1__27_, connection_0__1__26_, connection_0__1__25_, 
        connection_0__1__24_, connection_0__1__23_, connection_0__1__22_, 
        connection_0__1__21_, connection_0__1__20_, connection_0__1__19_, 
        connection_0__1__18_, connection_0__1__17_, connection_0__1__16_, 
        connection_0__1__15_, connection_0__1__14_, connection_0__1__13_, 
        connection_0__1__12_, connection_0__1__11_, connection_0__1__10_, 
        connection_0__1__9_, connection_0__1__8_, connection_0__1__7_, 
        connection_0__1__6_, connection_0__1__5_, connection_0__1__4_, 
        connection_0__1__3_, connection_0__1__2_, connection_0__1__1_, 
        connection_0__1__0_, connection_0__0__31_, connection_0__0__30_, 
        connection_0__0__29_, connection_0__0__28_, connection_0__0__27_, 
        connection_0__0__26_, connection_0__0__25_, connection_0__0__24_, 
        connection_0__0__23_, connection_0__0__22_, connection_0__0__21_, 
        connection_0__0__20_, connection_0__0__19_, connection_0__0__18_, 
        connection_0__0__17_, connection_0__0__16_, connection_0__0__15_, 
        connection_0__0__14_, connection_0__0__13_, connection_0__0__12_, 
        connection_0__0__11_, connection_0__0__10_, connection_0__0__9_, 
        connection_0__0__8_, connection_0__0__7_, connection_0__0__6_, 
        connection_0__0__5_, connection_0__0__4_, connection_0__0__3_, 
        connection_0__0__2_, connection_0__0__1_, connection_0__0__0_}), 
        .i_fwd_valid(fwd_connection_valid_frist_half[23]), .i_fwd_data_bus(
        fwd_connection_frist_half[767:736]), .o_fwd_valid(
        fwd_connection_valid_frist_half[19]), .o_fwd_data_bus(
        fwd_connection_frist_half[639:608]), .i_en(n533), .i_cmd(i_cmd[4:0])
         );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_47 first_half_stages_0__sw_group_0__upper_group_1__genblk1_upper_sw_first_stage ( 
        .clk(clk), .rst(n532), .i_valid(i_valid[3:2]), .i_data_bus(
        i_data_bus[127:64]), .o_valid({connection_valid_0__3_, 
        connection_valid_0__2_}), .o_data_bus({connection_0__3__31_, 
        connection_0__3__30_, connection_0__3__29_, connection_0__3__28_, 
        connection_0__3__27_, connection_0__3__26_, connection_0__3__25_, 
        connection_0__3__24_, connection_0__3__23_, connection_0__3__22_, 
        connection_0__3__21_, connection_0__3__20_, connection_0__3__19_, 
        connection_0__3__18_, connection_0__3__17_, connection_0__3__16_, 
        connection_0__3__15_, connection_0__3__14_, connection_0__3__13_, 
        connection_0__3__12_, connection_0__3__11_, connection_0__3__10_, 
        connection_0__3__9_, connection_0__3__8_, connection_0__3__7_, 
        connection_0__3__6_, connection_0__3__5_, connection_0__3__4_, 
        connection_0__3__3_, connection_0__3__2_, connection_0__3__1_, 
        connection_0__3__0_, connection_0__2__31_, connection_0__2__30_, 
        connection_0__2__29_, connection_0__2__28_, connection_0__2__27_, 
        connection_0__2__26_, connection_0__2__25_, connection_0__2__24_, 
        connection_0__2__23_, connection_0__2__22_, connection_0__2__21_, 
        connection_0__2__20_, connection_0__2__19_, connection_0__2__18_, 
        connection_0__2__17_, connection_0__2__16_, connection_0__2__15_, 
        connection_0__2__14_, connection_0__2__13_, connection_0__2__12_, 
        connection_0__2__11_, connection_0__2__10_, connection_0__2__9_, 
        connection_0__2__8_, connection_0__2__7_, connection_0__2__6_, 
        connection_0__2__5_, connection_0__2__4_, connection_0__2__3_, 
        connection_0__2__2_, connection_0__2__1_, connection_0__2__0_}), 
        .i_fwd_valid(fwd_connection_valid_frist_half[22]), .i_fwd_data_bus(
        fwd_connection_frist_half[735:704]), .o_fwd_valid(
        fwd_connection_valid_frist_half[18]), .o_fwd_data_bus(
        fwd_connection_frist_half[607:576]), .i_en(i_en), .i_cmd(i_cmd[9:5])
         );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_46 first_half_stages_0__sw_group_0__upper_group_2__genblk1_upper_sw_first_stage ( 
        .clk(clk), .rst(n532), .i_valid(i_valid[5:4]), .i_data_bus(
        i_data_bus[191:128]), .o_valid({connection_valid_0__5_, 
        connection_valid_0__4_}), .o_data_bus({connection_0__5__31_, 
        connection_0__5__30_, connection_0__5__29_, connection_0__5__28_, 
        connection_0__5__27_, connection_0__5__26_, connection_0__5__25_, 
        connection_0__5__24_, connection_0__5__23_, connection_0__5__22_, 
        connection_0__5__21_, connection_0__5__20_, connection_0__5__19_, 
        connection_0__5__18_, connection_0__5__17_, connection_0__5__16_, 
        connection_0__5__15_, connection_0__5__14_, connection_0__5__13_, 
        connection_0__5__12_, connection_0__5__11_, connection_0__5__10_, 
        connection_0__5__9_, connection_0__5__8_, connection_0__5__7_, 
        connection_0__5__6_, connection_0__5__5_, connection_0__5__4_, 
        connection_0__5__3_, connection_0__5__2_, connection_0__5__1_, 
        connection_0__5__0_, connection_0__4__31_, connection_0__4__30_, 
        connection_0__4__29_, connection_0__4__28_, connection_0__4__27_, 
        connection_0__4__26_, connection_0__4__25_, connection_0__4__24_, 
        connection_0__4__23_, connection_0__4__22_, connection_0__4__21_, 
        connection_0__4__20_, connection_0__4__19_, connection_0__4__18_, 
        connection_0__4__17_, connection_0__4__16_, connection_0__4__15_, 
        connection_0__4__14_, connection_0__4__13_, connection_0__4__12_, 
        connection_0__4__11_, connection_0__4__10_, connection_0__4__9_, 
        connection_0__4__8_, connection_0__4__7_, connection_0__4__6_, 
        connection_0__4__5_, connection_0__4__4_, connection_0__4__3_, 
        connection_0__4__2_, connection_0__4__1_, connection_0__4__0_}), 
        .i_fwd_valid(fwd_connection_valid_frist_half[21]), .i_fwd_data_bus(
        fwd_connection_frist_half[703:672]), .o_fwd_valid(
        fwd_connection_valid_frist_half[17]), .o_fwd_data_bus(
        fwd_connection_frist_half[575:544]), .i_en(n533), .i_cmd(i_cmd[14:10])
         );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_45 first_half_stages_0__sw_group_0__upper_group_3__genblk1_upper_sw_first_stage ( 
        .clk(clk), .rst(n532), .i_valid(i_valid[7:6]), .i_data_bus(
        i_data_bus[255:192]), .o_valid({connection_valid_0__7_, 
        connection_valid_0__6_}), .o_data_bus({connection_0__7__31_, 
        connection_0__7__30_, connection_0__7__29_, connection_0__7__28_, 
        connection_0__7__27_, connection_0__7__26_, connection_0__7__25_, 
        connection_0__7__24_, connection_0__7__23_, connection_0__7__22_, 
        connection_0__7__21_, connection_0__7__20_, connection_0__7__19_, 
        connection_0__7__18_, connection_0__7__17_, connection_0__7__16_, 
        connection_0__7__15_, connection_0__7__14_, connection_0__7__13_, 
        connection_0__7__12_, connection_0__7__11_, connection_0__7__10_, 
        connection_0__7__9_, connection_0__7__8_, connection_0__7__7_, 
        connection_0__7__6_, connection_0__7__5_, connection_0__7__4_, 
        connection_0__7__3_, connection_0__7__2_, connection_0__7__1_, 
        connection_0__7__0_, connection_0__6__31_, connection_0__6__30_, 
        connection_0__6__29_, connection_0__6__28_, connection_0__6__27_, 
        connection_0__6__26_, connection_0__6__25_, connection_0__6__24_, 
        connection_0__6__23_, connection_0__6__22_, connection_0__6__21_, 
        connection_0__6__20_, connection_0__6__19_, connection_0__6__18_, 
        connection_0__6__17_, connection_0__6__16_, connection_0__6__15_, 
        connection_0__6__14_, connection_0__6__13_, connection_0__6__12_, 
        connection_0__6__11_, connection_0__6__10_, connection_0__6__9_, 
        connection_0__6__8_, connection_0__6__7_, connection_0__6__6_, 
        connection_0__6__5_, connection_0__6__4_, connection_0__6__3_, 
        connection_0__6__2_, connection_0__6__1_, connection_0__6__0_}), 
        .i_fwd_valid(fwd_connection_valid_frist_half[20]), .i_fwd_data_bus(
        fwd_connection_frist_half[671:640]), .o_fwd_valid(
        fwd_connection_valid_frist_half[16]), .o_fwd_data_bus(
        fwd_connection_frist_half[543:512]), .i_en(i_en), .i_cmd(i_cmd[19:15])
         );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_44 first_half_stages_0__sw_group_0__bottom_group_0__genblk1_bottom_sw_first_stage ( 
        .clk(clk), .rst(n532), .i_valid(i_valid[9:8]), .i_data_bus(
        i_data_bus[319:256]), .o_valid({connection_valid_0__9_, 
        connection_valid_0__8_}), .o_data_bus({connection_0__9__31_, 
        connection_0__9__30_, connection_0__9__29_, connection_0__9__28_, 
        connection_0__9__27_, connection_0__9__26_, connection_0__9__25_, 
        connection_0__9__24_, connection_0__9__23_, connection_0__9__22_, 
        connection_0__9__21_, connection_0__9__20_, connection_0__9__19_, 
        connection_0__9__18_, connection_0__9__17_, connection_0__9__16_, 
        connection_0__9__15_, connection_0__9__14_, connection_0__9__13_, 
        connection_0__9__12_, connection_0__9__11_, connection_0__9__10_, 
        connection_0__9__9_, connection_0__9__8_, connection_0__9__7_, 
        connection_0__9__6_, connection_0__9__5_, connection_0__9__4_, 
        connection_0__9__3_, connection_0__9__2_, connection_0__9__1_, 
        connection_0__9__0_, connection_0__8__31_, connection_0__8__30_, 
        connection_0__8__29_, connection_0__8__28_, connection_0__8__27_, 
        connection_0__8__26_, connection_0__8__25_, connection_0__8__24_, 
        connection_0__8__23_, connection_0__8__22_, connection_0__8__21_, 
        connection_0__8__20_, connection_0__8__19_, connection_0__8__18_, 
        connection_0__8__17_, connection_0__8__16_, connection_0__8__15_, 
        connection_0__8__14_, connection_0__8__13_, connection_0__8__12_, 
        connection_0__8__11_, connection_0__8__10_, connection_0__8__9_, 
        connection_0__8__8_, connection_0__8__7_, connection_0__8__6_, 
        connection_0__8__5_, connection_0__8__4_, connection_0__8__3_, 
        connection_0__8__2_, connection_0__8__1_, connection_0__8__0_}), 
        .i_fwd_valid(fwd_connection_valid_frist_half[19]), .i_fwd_data_bus(
        fwd_connection_frist_half[639:608]), .o_fwd_valid(
        fwd_connection_valid_frist_half[23]), .o_fwd_data_bus(
        fwd_connection_frist_half[767:736]), .i_en(i_en), .i_cmd(i_cmd[24:20])
         );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_43 first_half_stages_0__sw_group_0__bottom_group_1__genblk1_bottom_sw_first_stage ( 
        .clk(clk), .rst(n532), .i_valid(i_valid[11:10]), .i_data_bus(
        i_data_bus[383:320]), .o_valid({connection_valid_0__11_, 
        connection_valid_0__10_}), .o_data_bus({connection_0__11__31_, 
        connection_0__11__30_, connection_0__11__29_, connection_0__11__28_, 
        connection_0__11__27_, connection_0__11__26_, connection_0__11__25_, 
        connection_0__11__24_, connection_0__11__23_, connection_0__11__22_, 
        connection_0__11__21_, connection_0__11__20_, connection_0__11__19_, 
        connection_0__11__18_, connection_0__11__17_, connection_0__11__16_, 
        connection_0__11__15_, connection_0__11__14_, connection_0__11__13_, 
        connection_0__11__12_, connection_0__11__11_, connection_0__11__10_, 
        connection_0__11__9_, connection_0__11__8_, connection_0__11__7_, 
        connection_0__11__6_, connection_0__11__5_, connection_0__11__4_, 
        connection_0__11__3_, connection_0__11__2_, connection_0__11__1_, 
        connection_0__11__0_, connection_0__10__31_, connection_0__10__30_, 
        connection_0__10__29_, connection_0__10__28_, connection_0__10__27_, 
        connection_0__10__26_, connection_0__10__25_, connection_0__10__24_, 
        connection_0__10__23_, connection_0__10__22_, connection_0__10__21_, 
        connection_0__10__20_, connection_0__10__19_, connection_0__10__18_, 
        connection_0__10__17_, connection_0__10__16_, connection_0__10__15_, 
        connection_0__10__14_, connection_0__10__13_, connection_0__10__12_, 
        connection_0__10__11_, connection_0__10__10_, connection_0__10__9_, 
        connection_0__10__8_, connection_0__10__7_, connection_0__10__6_, 
        connection_0__10__5_, connection_0__10__4_, connection_0__10__3_, 
        connection_0__10__2_, connection_0__10__1_, connection_0__10__0_}), 
        .i_fwd_valid(fwd_connection_valid_frist_half[18]), .i_fwd_data_bus(
        fwd_connection_frist_half[607:576]), .o_fwd_valid(
        fwd_connection_valid_frist_half[22]), .o_fwd_data_bus(
        fwd_connection_frist_half[735:704]), .i_en(i_en), .i_cmd(i_cmd[29:25])
         );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_42 first_half_stages_0__sw_group_0__bottom_group_2__genblk1_bottom_sw_first_stage ( 
        .clk(clk), .rst(n532), .i_valid(i_valid[13:12]), .i_data_bus(
        i_data_bus[447:384]), .o_valid({connection_valid_0__13_, 
        connection_valid_0__12_}), .o_data_bus({connection_0__13__31_, 
        connection_0__13__30_, connection_0__13__29_, connection_0__13__28_, 
        connection_0__13__27_, connection_0__13__26_, connection_0__13__25_, 
        connection_0__13__24_, connection_0__13__23_, connection_0__13__22_, 
        connection_0__13__21_, connection_0__13__20_, connection_0__13__19_, 
        connection_0__13__18_, connection_0__13__17_, connection_0__13__16_, 
        connection_0__13__15_, connection_0__13__14_, connection_0__13__13_, 
        connection_0__13__12_, connection_0__13__11_, connection_0__13__10_, 
        connection_0__13__9_, connection_0__13__8_, connection_0__13__7_, 
        connection_0__13__6_, connection_0__13__5_, connection_0__13__4_, 
        connection_0__13__3_, connection_0__13__2_, connection_0__13__1_, 
        connection_0__13__0_, connection_0__12__31_, connection_0__12__30_, 
        connection_0__12__29_, connection_0__12__28_, connection_0__12__27_, 
        connection_0__12__26_, connection_0__12__25_, connection_0__12__24_, 
        connection_0__12__23_, connection_0__12__22_, connection_0__12__21_, 
        connection_0__12__20_, connection_0__12__19_, connection_0__12__18_, 
        connection_0__12__17_, connection_0__12__16_, connection_0__12__15_, 
        connection_0__12__14_, connection_0__12__13_, connection_0__12__12_, 
        connection_0__12__11_, connection_0__12__10_, connection_0__12__9_, 
        connection_0__12__8_, connection_0__12__7_, connection_0__12__6_, 
        connection_0__12__5_, connection_0__12__4_, connection_0__12__3_, 
        connection_0__12__2_, connection_0__12__1_, connection_0__12__0_}), 
        .i_fwd_valid(fwd_connection_valid_frist_half[17]), .i_fwd_data_bus(
        fwd_connection_frist_half[575:544]), .o_fwd_valid(
        fwd_connection_valid_frist_half[21]), .o_fwd_data_bus(
        fwd_connection_frist_half[703:672]), .i_en(n533), .i_cmd(i_cmd[34:30])
         );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_41 first_half_stages_0__sw_group_0__bottom_group_3__genblk1_bottom_sw_first_stage ( 
        .clk(clk), .rst(n532), .i_valid(i_valid[15:14]), .i_data_bus(
        i_data_bus[511:448]), .o_valid({connection_valid_0__15_, 
        connection_valid_0__14_}), .o_data_bus({connection_0__15__31_, 
        connection_0__15__30_, connection_0__15__29_, connection_0__15__28_, 
        connection_0__15__27_, connection_0__15__26_, connection_0__15__25_, 
        connection_0__15__24_, connection_0__15__23_, connection_0__15__22_, 
        connection_0__15__21_, connection_0__15__20_, connection_0__15__19_, 
        connection_0__15__18_, connection_0__15__17_, connection_0__15__16_, 
        connection_0__15__15_, connection_0__15__14_, connection_0__15__13_, 
        connection_0__15__12_, connection_0__15__11_, connection_0__15__10_, 
        connection_0__15__9_, connection_0__15__8_, connection_0__15__7_, 
        connection_0__15__6_, connection_0__15__5_, connection_0__15__4_, 
        connection_0__15__3_, connection_0__15__2_, connection_0__15__1_, 
        connection_0__15__0_, connection_0__14__31_, connection_0__14__30_, 
        connection_0__14__29_, connection_0__14__28_, connection_0__14__27_, 
        connection_0__14__26_, connection_0__14__25_, connection_0__14__24_, 
        connection_0__14__23_, connection_0__14__22_, connection_0__14__21_, 
        connection_0__14__20_, connection_0__14__19_, connection_0__14__18_, 
        connection_0__14__17_, connection_0__14__16_, connection_0__14__15_, 
        connection_0__14__14_, connection_0__14__13_, connection_0__14__12_, 
        connection_0__14__11_, connection_0__14__10_, connection_0__14__9_, 
        connection_0__14__8_, connection_0__14__7_, connection_0__14__6_, 
        connection_0__14__5_, connection_0__14__4_, connection_0__14__3_, 
        connection_0__14__2_, connection_0__14__1_, connection_0__14__0_}), 
        .i_fwd_valid(fwd_connection_valid_frist_half[16]), .i_fwd_data_bus(
        fwd_connection_frist_half[543:512]), .o_fwd_valid(
        fwd_connection_valid_frist_half[20]), .o_fwd_data_bus(
        fwd_connection_frist_half[671:640]), .i_en(i_en), .i_cmd(i_cmd[39:35])
         );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_40 first_half_stages_1__sw_group_0__upper_group_0__genblk1_upper_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_0__1_, 
        connection_valid_0__0_}), .i_data_bus({connection_0__1__31_, 
        connection_0__1__30_, connection_0__1__29_, connection_0__1__28_, 
        connection_0__1__27_, connection_0__1__26_, connection_0__1__25_, 
        connection_0__1__24_, connection_0__1__23_, connection_0__1__22_, 
        connection_0__1__21_, connection_0__1__20_, connection_0__1__19_, 
        connection_0__1__18_, connection_0__1__17_, connection_0__1__16_, 
        connection_0__1__15_, connection_0__1__14_, connection_0__1__13_, 
        connection_0__1__12_, connection_0__1__11_, connection_0__1__10_, 
        connection_0__1__9_, connection_0__1__8_, connection_0__1__7_, 
        connection_0__1__6_, connection_0__1__5_, connection_0__1__4_, 
        connection_0__1__3_, connection_0__1__2_, connection_0__1__1_, 
        connection_0__1__0_, connection_0__0__31_, connection_0__0__30_, 
        connection_0__0__29_, connection_0__0__28_, connection_0__0__27_, 
        connection_0__0__26_, connection_0__0__25_, connection_0__0__24_, 
        connection_0__0__23_, connection_0__0__22_, connection_0__0__21_, 
        connection_0__0__20_, connection_0__0__19_, connection_0__0__18_, 
        connection_0__0__17_, connection_0__0__16_, connection_0__0__15_, 
        connection_0__0__14_, connection_0__0__13_, connection_0__0__12_, 
        connection_0__0__11_, connection_0__0__10_, connection_0__0__9_, 
        connection_0__0__8_, connection_0__0__7_, connection_0__0__6_, 
        connection_0__0__5_, connection_0__0__4_, connection_0__0__3_, 
        connection_0__0__2_, connection_0__0__1_, connection_0__0__0_}), 
        .o_valid({connection_valid_1__1_, connection_valid_1__0_}), 
        .o_data_bus({connection_1__1__31_, connection_1__1__30_, 
        connection_1__1__29_, connection_1__1__28_, connection_1__1__27_, 
        connection_1__1__26_, connection_1__1__25_, connection_1__1__24_, 
        connection_1__1__23_, connection_1__1__22_, connection_1__1__21_, 
        connection_1__1__20_, connection_1__1__19_, connection_1__1__18_, 
        connection_1__1__17_, connection_1__1__16_, connection_1__1__15_, 
        connection_1__1__14_, connection_1__1__13_, connection_1__1__12_, 
        connection_1__1__11_, connection_1__1__10_, connection_1__1__9_, 
        connection_1__1__8_, connection_1__1__7_, connection_1__1__6_, 
        connection_1__1__5_, connection_1__1__4_, connection_1__1__3_, 
        connection_1__1__2_, connection_1__1__1_, connection_1__1__0_, 
        connection_1__0__31_, connection_1__0__30_, connection_1__0__29_, 
        connection_1__0__28_, connection_1__0__27_, connection_1__0__26_, 
        connection_1__0__25_, connection_1__0__24_, connection_1__0__23_, 
        connection_1__0__22_, connection_1__0__21_, connection_1__0__20_, 
        connection_1__0__19_, connection_1__0__18_, connection_1__0__17_, 
        connection_1__0__16_, connection_1__0__15_, connection_1__0__14_, 
        connection_1__0__13_, connection_1__0__12_, connection_1__0__11_, 
        connection_1__0__10_, connection_1__0__9_, connection_1__0__8_, 
        connection_1__0__7_, connection_1__0__6_, connection_1__0__5_, 
        connection_1__0__4_, connection_1__0__3_, connection_1__0__2_, 
        connection_1__0__1_, connection_1__0__0_}), .i_fwd_valid(
        fwd_connection_valid_frist_half[15]), .i_fwd_data_bus(
        fwd_connection_frist_half[511:480]), .o_fwd_valid(
        fwd_connection_valid_frist_half[13]), .o_fwd_data_bus(
        fwd_connection_frist_half[447:416]), .i_en(n533), .i_cmd({
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__0__4_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__0__3_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__0__2_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__0__1_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__0__0_}) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_39 first_half_stages_1__sw_group_0__upper_group_1__genblk1_upper_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_0__3_, 
        connection_valid_0__2_}), .i_data_bus({connection_0__3__31_, 
        connection_0__3__30_, connection_0__3__29_, connection_0__3__28_, 
        connection_0__3__27_, connection_0__3__26_, connection_0__3__25_, 
        connection_0__3__24_, connection_0__3__23_, connection_0__3__22_, 
        connection_0__3__21_, connection_0__3__20_, connection_0__3__19_, 
        connection_0__3__18_, connection_0__3__17_, connection_0__3__16_, 
        connection_0__3__15_, connection_0__3__14_, connection_0__3__13_, 
        connection_0__3__12_, connection_0__3__11_, connection_0__3__10_, 
        connection_0__3__9_, connection_0__3__8_, connection_0__3__7_, 
        connection_0__3__6_, connection_0__3__5_, connection_0__3__4_, 
        connection_0__3__3_, connection_0__3__2_, connection_0__3__1_, 
        connection_0__3__0_, connection_0__2__31_, connection_0__2__30_, 
        connection_0__2__29_, connection_0__2__28_, connection_0__2__27_, 
        connection_0__2__26_, connection_0__2__25_, connection_0__2__24_, 
        connection_0__2__23_, connection_0__2__22_, connection_0__2__21_, 
        connection_0__2__20_, connection_0__2__19_, connection_0__2__18_, 
        connection_0__2__17_, connection_0__2__16_, connection_0__2__15_, 
        connection_0__2__14_, connection_0__2__13_, connection_0__2__12_, 
        connection_0__2__11_, connection_0__2__10_, connection_0__2__9_, 
        connection_0__2__8_, connection_0__2__7_, connection_0__2__6_, 
        connection_0__2__5_, connection_0__2__4_, connection_0__2__3_, 
        connection_0__2__2_, connection_0__2__1_, connection_0__2__0_}), 
        .o_valid({connection_valid_1__3_, connection_valid_1__2_}), 
        .o_data_bus({connection_1__3__31_, connection_1__3__30_, 
        connection_1__3__29_, connection_1__3__28_, connection_1__3__27_, 
        connection_1__3__26_, connection_1__3__25_, connection_1__3__24_, 
        connection_1__3__23_, connection_1__3__22_, connection_1__3__21_, 
        connection_1__3__20_, connection_1__3__19_, connection_1__3__18_, 
        connection_1__3__17_, connection_1__3__16_, connection_1__3__15_, 
        connection_1__3__14_, connection_1__3__13_, connection_1__3__12_, 
        connection_1__3__11_, connection_1__3__10_, connection_1__3__9_, 
        connection_1__3__8_, connection_1__3__7_, connection_1__3__6_, 
        connection_1__3__5_, connection_1__3__4_, connection_1__3__3_, 
        connection_1__3__2_, connection_1__3__1_, connection_1__3__0_, 
        connection_1__2__31_, connection_1__2__30_, connection_1__2__29_, 
        connection_1__2__28_, connection_1__2__27_, connection_1__2__26_, 
        connection_1__2__25_, connection_1__2__24_, connection_1__2__23_, 
        connection_1__2__22_, connection_1__2__21_, connection_1__2__20_, 
        connection_1__2__19_, connection_1__2__18_, connection_1__2__17_, 
        connection_1__2__16_, connection_1__2__15_, connection_1__2__14_, 
        connection_1__2__13_, connection_1__2__12_, connection_1__2__11_, 
        connection_1__2__10_, connection_1__2__9_, connection_1__2__8_, 
        connection_1__2__7_, connection_1__2__6_, connection_1__2__5_, 
        connection_1__2__4_, connection_1__2__3_, connection_1__2__2_, 
        connection_1__2__1_, connection_1__2__0_}), .i_fwd_valid(
        fwd_connection_valid_frist_half[14]), .i_fwd_data_bus(
        fwd_connection_frist_half[479:448]), .o_fwd_valid(
        fwd_connection_valid_frist_half[12]), .o_fwd_data_bus(
        fwd_connection_frist_half[415:384]), .i_en(n533), .i_cmd({
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__1__4_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__1__3_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__1__2_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__1__1_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__1__0_}) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_38 first_half_stages_1__sw_group_0__bottom_group_0__genblk1_bottom_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_0__5_, 
        connection_valid_0__4_}), .i_data_bus({connection_0__5__31_, 
        connection_0__5__30_, connection_0__5__29_, connection_0__5__28_, 
        connection_0__5__27_, connection_0__5__26_, connection_0__5__25_, 
        connection_0__5__24_, connection_0__5__23_, connection_0__5__22_, 
        connection_0__5__21_, connection_0__5__20_, connection_0__5__19_, 
        connection_0__5__18_, connection_0__5__17_, connection_0__5__16_, 
        connection_0__5__15_, connection_0__5__14_, connection_0__5__13_, 
        connection_0__5__12_, connection_0__5__11_, connection_0__5__10_, 
        connection_0__5__9_, connection_0__5__8_, connection_0__5__7_, 
        connection_0__5__6_, connection_0__5__5_, connection_0__5__4_, 
        connection_0__5__3_, connection_0__5__2_, connection_0__5__1_, 
        connection_0__5__0_, connection_0__4__31_, connection_0__4__30_, 
        connection_0__4__29_, connection_0__4__28_, connection_0__4__27_, 
        connection_0__4__26_, connection_0__4__25_, connection_0__4__24_, 
        connection_0__4__23_, connection_0__4__22_, connection_0__4__21_, 
        connection_0__4__20_, connection_0__4__19_, connection_0__4__18_, 
        connection_0__4__17_, connection_0__4__16_, connection_0__4__15_, 
        connection_0__4__14_, connection_0__4__13_, connection_0__4__12_, 
        connection_0__4__11_, connection_0__4__10_, connection_0__4__9_, 
        connection_0__4__8_, connection_0__4__7_, connection_0__4__6_, 
        connection_0__4__5_, connection_0__4__4_, connection_0__4__3_, 
        connection_0__4__2_, connection_0__4__1_, connection_0__4__0_}), 
        .o_valid({connection_valid_1__5_, connection_valid_1__4_}), 
        .o_data_bus({connection_1__5__31_, connection_1__5__30_, 
        connection_1__5__29_, connection_1__5__28_, connection_1__5__27_, 
        connection_1__5__26_, connection_1__5__25_, connection_1__5__24_, 
        connection_1__5__23_, connection_1__5__22_, connection_1__5__21_, 
        connection_1__5__20_, connection_1__5__19_, connection_1__5__18_, 
        connection_1__5__17_, connection_1__5__16_, connection_1__5__15_, 
        connection_1__5__14_, connection_1__5__13_, connection_1__5__12_, 
        connection_1__5__11_, connection_1__5__10_, connection_1__5__9_, 
        connection_1__5__8_, connection_1__5__7_, connection_1__5__6_, 
        connection_1__5__5_, connection_1__5__4_, connection_1__5__3_, 
        connection_1__5__2_, connection_1__5__1_, connection_1__5__0_, 
        connection_1__4__31_, connection_1__4__30_, connection_1__4__29_, 
        connection_1__4__28_, connection_1__4__27_, connection_1__4__26_, 
        connection_1__4__25_, connection_1__4__24_, connection_1__4__23_, 
        connection_1__4__22_, connection_1__4__21_, connection_1__4__20_, 
        connection_1__4__19_, connection_1__4__18_, connection_1__4__17_, 
        connection_1__4__16_, connection_1__4__15_, connection_1__4__14_, 
        connection_1__4__13_, connection_1__4__12_, connection_1__4__11_, 
        connection_1__4__10_, connection_1__4__9_, connection_1__4__8_, 
        connection_1__4__7_, connection_1__4__6_, connection_1__4__5_, 
        connection_1__4__4_, connection_1__4__3_, connection_1__4__2_, 
        connection_1__4__1_, connection_1__4__0_}), .i_fwd_valid(
        fwd_connection_valid_frist_half[13]), .i_fwd_data_bus(
        fwd_connection_frist_half[447:416]), .o_fwd_valid(
        fwd_connection_valid_frist_half[15]), .o_fwd_data_bus(
        fwd_connection_frist_half[511:480]), .i_en(i_en), .i_cmd({
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__2__4_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__2__3_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__2__2_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__2__1_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__2__0_}) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_37 first_half_stages_1__sw_group_0__bottom_group_1__genblk1_bottom_sw ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__7_, 
        connection_valid_0__6_}), .i_data_bus({connection_0__7__31_, 
        connection_0__7__30_, connection_0__7__29_, connection_0__7__28_, 
        connection_0__7__27_, connection_0__7__26_, connection_0__7__25_, 
        connection_0__7__24_, connection_0__7__23_, connection_0__7__22_, 
        connection_0__7__21_, connection_0__7__20_, connection_0__7__19_, 
        connection_0__7__18_, connection_0__7__17_, connection_0__7__16_, 
        connection_0__7__15_, connection_0__7__14_, connection_0__7__13_, 
        connection_0__7__12_, connection_0__7__11_, connection_0__7__10_, 
        connection_0__7__9_, connection_0__7__8_, connection_0__7__7_, 
        connection_0__7__6_, connection_0__7__5_, connection_0__7__4_, 
        connection_0__7__3_, connection_0__7__2_, connection_0__7__1_, 
        connection_0__7__0_, connection_0__6__31_, connection_0__6__30_, 
        connection_0__6__29_, connection_0__6__28_, connection_0__6__27_, 
        connection_0__6__26_, connection_0__6__25_, connection_0__6__24_, 
        connection_0__6__23_, connection_0__6__22_, connection_0__6__21_, 
        connection_0__6__20_, connection_0__6__19_, connection_0__6__18_, 
        connection_0__6__17_, connection_0__6__16_, connection_0__6__15_, 
        connection_0__6__14_, connection_0__6__13_, connection_0__6__12_, 
        connection_0__6__11_, connection_0__6__10_, connection_0__6__9_, 
        connection_0__6__8_, connection_0__6__7_, connection_0__6__6_, 
        connection_0__6__5_, connection_0__6__4_, connection_0__6__3_, 
        connection_0__6__2_, connection_0__6__1_, connection_0__6__0_}), 
        .o_valid({connection_valid_1__7_, connection_valid_1__6_}), 
        .o_data_bus({connection_1__7__31_, connection_1__7__30_, 
        connection_1__7__29_, connection_1__7__28_, connection_1__7__27_, 
        connection_1__7__26_, connection_1__7__25_, connection_1__7__24_, 
        connection_1__7__23_, connection_1__7__22_, connection_1__7__21_, 
        connection_1__7__20_, connection_1__7__19_, connection_1__7__18_, 
        connection_1__7__17_, connection_1__7__16_, connection_1__7__15_, 
        connection_1__7__14_, connection_1__7__13_, connection_1__7__12_, 
        connection_1__7__11_, connection_1__7__10_, connection_1__7__9_, 
        connection_1__7__8_, connection_1__7__7_, connection_1__7__6_, 
        connection_1__7__5_, connection_1__7__4_, connection_1__7__3_, 
        connection_1__7__2_, connection_1__7__1_, connection_1__7__0_, 
        connection_1__6__31_, connection_1__6__30_, connection_1__6__29_, 
        connection_1__6__28_, connection_1__6__27_, connection_1__6__26_, 
        connection_1__6__25_, connection_1__6__24_, connection_1__6__23_, 
        connection_1__6__22_, connection_1__6__21_, connection_1__6__20_, 
        connection_1__6__19_, connection_1__6__18_, connection_1__6__17_, 
        connection_1__6__16_, connection_1__6__15_, connection_1__6__14_, 
        connection_1__6__13_, connection_1__6__12_, connection_1__6__11_, 
        connection_1__6__10_, connection_1__6__9_, connection_1__6__8_, 
        connection_1__6__7_, connection_1__6__6_, connection_1__6__5_, 
        connection_1__6__4_, connection_1__6__3_, connection_1__6__2_, 
        connection_1__6__1_, connection_1__6__0_}), .i_fwd_valid(
        fwd_connection_valid_frist_half[12]), .i_fwd_data_bus(
        fwd_connection_frist_half[415:384]), .o_fwd_valid(
        fwd_connection_valid_frist_half[14]), .o_fwd_data_bus(
        fwd_connection_frist_half[479:448]), .i_en(n533), .i_cmd({
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__3__4_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__3__3_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__3__2_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__3__1_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__3__0_}) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_36 first_half_stages_1__sw_group_1__upper_group_0__genblk1_upper_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_0__9_, 
        connection_valid_0__8_}), .i_data_bus({connection_0__9__31_, 
        connection_0__9__30_, connection_0__9__29_, connection_0__9__28_, 
        connection_0__9__27_, connection_0__9__26_, connection_0__9__25_, 
        connection_0__9__24_, connection_0__9__23_, connection_0__9__22_, 
        connection_0__9__21_, connection_0__9__20_, connection_0__9__19_, 
        connection_0__9__18_, connection_0__9__17_, connection_0__9__16_, 
        connection_0__9__15_, connection_0__9__14_, connection_0__9__13_, 
        connection_0__9__12_, connection_0__9__11_, connection_0__9__10_, 
        connection_0__9__9_, connection_0__9__8_, connection_0__9__7_, 
        connection_0__9__6_, connection_0__9__5_, connection_0__9__4_, 
        connection_0__9__3_, connection_0__9__2_, connection_0__9__1_, 
        connection_0__9__0_, connection_0__8__31_, connection_0__8__30_, 
        connection_0__8__29_, connection_0__8__28_, connection_0__8__27_, 
        connection_0__8__26_, connection_0__8__25_, connection_0__8__24_, 
        connection_0__8__23_, connection_0__8__22_, connection_0__8__21_, 
        connection_0__8__20_, connection_0__8__19_, connection_0__8__18_, 
        connection_0__8__17_, connection_0__8__16_, connection_0__8__15_, 
        connection_0__8__14_, connection_0__8__13_, connection_0__8__12_, 
        connection_0__8__11_, connection_0__8__10_, connection_0__8__9_, 
        connection_0__8__8_, connection_0__8__7_, connection_0__8__6_, 
        connection_0__8__5_, connection_0__8__4_, connection_0__8__3_, 
        connection_0__8__2_, connection_0__8__1_, connection_0__8__0_}), 
        .o_valid({connection_valid_1__9_, connection_valid_1__8_}), 
        .o_data_bus({connection_1__9__31_, connection_1__9__30_, 
        connection_1__9__29_, connection_1__9__28_, connection_1__9__27_, 
        connection_1__9__26_, connection_1__9__25_, connection_1__9__24_, 
        connection_1__9__23_, connection_1__9__22_, connection_1__9__21_, 
        connection_1__9__20_, connection_1__9__19_, connection_1__9__18_, 
        connection_1__9__17_, connection_1__9__16_, connection_1__9__15_, 
        connection_1__9__14_, connection_1__9__13_, connection_1__9__12_, 
        connection_1__9__11_, connection_1__9__10_, connection_1__9__9_, 
        connection_1__9__8_, connection_1__9__7_, connection_1__9__6_, 
        connection_1__9__5_, connection_1__9__4_, connection_1__9__3_, 
        connection_1__9__2_, connection_1__9__1_, connection_1__9__0_, 
        connection_1__8__31_, connection_1__8__30_, connection_1__8__29_, 
        connection_1__8__28_, connection_1__8__27_, connection_1__8__26_, 
        connection_1__8__25_, connection_1__8__24_, connection_1__8__23_, 
        connection_1__8__22_, connection_1__8__21_, connection_1__8__20_, 
        connection_1__8__19_, connection_1__8__18_, connection_1__8__17_, 
        connection_1__8__16_, connection_1__8__15_, connection_1__8__14_, 
        connection_1__8__13_, connection_1__8__12_, connection_1__8__11_, 
        connection_1__8__10_, connection_1__8__9_, connection_1__8__8_, 
        connection_1__8__7_, connection_1__8__6_, connection_1__8__5_, 
        connection_1__8__4_, connection_1__8__3_, connection_1__8__2_, 
        connection_1__8__1_, connection_1__8__0_}), .i_fwd_valid(
        fwd_connection_valid_frist_half[11]), .i_fwd_data_bus(
        fwd_connection_frist_half[383:352]), .o_fwd_valid(
        fwd_connection_valid_frist_half[9]), .o_fwd_data_bus(
        fwd_connection_frist_half[319:288]), .i_en(n533), .i_cmd({
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__4__4_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__4__3_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__4__2_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__4__1_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__4__0_}) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_35 first_half_stages_1__sw_group_1__upper_group_1__genblk1_upper_sw ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__11_, 
        connection_valid_0__10_}), .i_data_bus({connection_0__11__31_, 
        connection_0__11__30_, connection_0__11__29_, connection_0__11__28_, 
        connection_0__11__27_, connection_0__11__26_, connection_0__11__25_, 
        connection_0__11__24_, connection_0__11__23_, connection_0__11__22_, 
        connection_0__11__21_, connection_0__11__20_, connection_0__11__19_, 
        connection_0__11__18_, connection_0__11__17_, connection_0__11__16_, 
        connection_0__11__15_, connection_0__11__14_, connection_0__11__13_, 
        connection_0__11__12_, connection_0__11__11_, connection_0__11__10_, 
        connection_0__11__9_, connection_0__11__8_, connection_0__11__7_, 
        connection_0__11__6_, connection_0__11__5_, connection_0__11__4_, 
        connection_0__11__3_, connection_0__11__2_, connection_0__11__1_, 
        connection_0__11__0_, connection_0__10__31_, connection_0__10__30_, 
        connection_0__10__29_, connection_0__10__28_, connection_0__10__27_, 
        connection_0__10__26_, connection_0__10__25_, connection_0__10__24_, 
        connection_0__10__23_, connection_0__10__22_, connection_0__10__21_, 
        connection_0__10__20_, connection_0__10__19_, connection_0__10__18_, 
        connection_0__10__17_, connection_0__10__16_, connection_0__10__15_, 
        connection_0__10__14_, connection_0__10__13_, connection_0__10__12_, 
        connection_0__10__11_, connection_0__10__10_, connection_0__10__9_, 
        connection_0__10__8_, connection_0__10__7_, connection_0__10__6_, 
        connection_0__10__5_, connection_0__10__4_, connection_0__10__3_, 
        connection_0__10__2_, connection_0__10__1_, connection_0__10__0_}), 
        .o_valid({connection_valid_1__11_, connection_valid_1__10_}), 
        .o_data_bus({connection_1__11__31_, connection_1__11__30_, 
        connection_1__11__29_, connection_1__11__28_, connection_1__11__27_, 
        connection_1__11__26_, connection_1__11__25_, connection_1__11__24_, 
        connection_1__11__23_, connection_1__11__22_, connection_1__11__21_, 
        connection_1__11__20_, connection_1__11__19_, connection_1__11__18_, 
        connection_1__11__17_, connection_1__11__16_, connection_1__11__15_, 
        connection_1__11__14_, connection_1__11__13_, connection_1__11__12_, 
        connection_1__11__11_, connection_1__11__10_, connection_1__11__9_, 
        connection_1__11__8_, connection_1__11__7_, connection_1__11__6_, 
        connection_1__11__5_, connection_1__11__4_, connection_1__11__3_, 
        connection_1__11__2_, connection_1__11__1_, connection_1__11__0_, 
        connection_1__10__31_, connection_1__10__30_, connection_1__10__29_, 
        connection_1__10__28_, connection_1__10__27_, connection_1__10__26_, 
        connection_1__10__25_, connection_1__10__24_, connection_1__10__23_, 
        connection_1__10__22_, connection_1__10__21_, connection_1__10__20_, 
        connection_1__10__19_, connection_1__10__18_, connection_1__10__17_, 
        connection_1__10__16_, connection_1__10__15_, connection_1__10__14_, 
        connection_1__10__13_, connection_1__10__12_, connection_1__10__11_, 
        connection_1__10__10_, connection_1__10__9_, connection_1__10__8_, 
        connection_1__10__7_, connection_1__10__6_, connection_1__10__5_, 
        connection_1__10__4_, connection_1__10__3_, connection_1__10__2_, 
        connection_1__10__1_, connection_1__10__0_}), .i_fwd_valid(
        fwd_connection_valid_frist_half[10]), .i_fwd_data_bus(
        fwd_connection_frist_half[351:320]), .o_fwd_valid(
        fwd_connection_valid_frist_half[8]), .o_fwd_data_bus(
        fwd_connection_frist_half[287:256]), .i_en(n533), .i_cmd({
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__5__4_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__5__3_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__5__2_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__5__1_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__5__0_}) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_34 first_half_stages_1__sw_group_1__bottom_group_0__genblk1_bottom_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_0__13_, 
        connection_valid_0__12_}), .i_data_bus({connection_0__13__31_, 
        connection_0__13__30_, connection_0__13__29_, connection_0__13__28_, 
        connection_0__13__27_, connection_0__13__26_, connection_0__13__25_, 
        connection_0__13__24_, connection_0__13__23_, connection_0__13__22_, 
        connection_0__13__21_, connection_0__13__20_, connection_0__13__19_, 
        connection_0__13__18_, connection_0__13__17_, connection_0__13__16_, 
        connection_0__13__15_, connection_0__13__14_, connection_0__13__13_, 
        connection_0__13__12_, connection_0__13__11_, connection_0__13__10_, 
        connection_0__13__9_, connection_0__13__8_, connection_0__13__7_, 
        connection_0__13__6_, connection_0__13__5_, connection_0__13__4_, 
        connection_0__13__3_, connection_0__13__2_, connection_0__13__1_, 
        connection_0__13__0_, connection_0__12__31_, connection_0__12__30_, 
        connection_0__12__29_, connection_0__12__28_, connection_0__12__27_, 
        connection_0__12__26_, connection_0__12__25_, connection_0__12__24_, 
        connection_0__12__23_, connection_0__12__22_, connection_0__12__21_, 
        connection_0__12__20_, connection_0__12__19_, connection_0__12__18_, 
        connection_0__12__17_, connection_0__12__16_, connection_0__12__15_, 
        connection_0__12__14_, connection_0__12__13_, connection_0__12__12_, 
        connection_0__12__11_, connection_0__12__10_, connection_0__12__9_, 
        connection_0__12__8_, connection_0__12__7_, connection_0__12__6_, 
        connection_0__12__5_, connection_0__12__4_, connection_0__12__3_, 
        connection_0__12__2_, connection_0__12__1_, connection_0__12__0_}), 
        .o_valid({connection_valid_1__13_, connection_valid_1__12_}), 
        .o_data_bus({connection_1__13__31_, connection_1__13__30_, 
        connection_1__13__29_, connection_1__13__28_, connection_1__13__27_, 
        connection_1__13__26_, connection_1__13__25_, connection_1__13__24_, 
        connection_1__13__23_, connection_1__13__22_, connection_1__13__21_, 
        connection_1__13__20_, connection_1__13__19_, connection_1__13__18_, 
        connection_1__13__17_, connection_1__13__16_, connection_1__13__15_, 
        connection_1__13__14_, connection_1__13__13_, connection_1__13__12_, 
        connection_1__13__11_, connection_1__13__10_, connection_1__13__9_, 
        connection_1__13__8_, connection_1__13__7_, connection_1__13__6_, 
        connection_1__13__5_, connection_1__13__4_, connection_1__13__3_, 
        connection_1__13__2_, connection_1__13__1_, connection_1__13__0_, 
        connection_1__12__31_, connection_1__12__30_, connection_1__12__29_, 
        connection_1__12__28_, connection_1__12__27_, connection_1__12__26_, 
        connection_1__12__25_, connection_1__12__24_, connection_1__12__23_, 
        connection_1__12__22_, connection_1__12__21_, connection_1__12__20_, 
        connection_1__12__19_, connection_1__12__18_, connection_1__12__17_, 
        connection_1__12__16_, connection_1__12__15_, connection_1__12__14_, 
        connection_1__12__13_, connection_1__12__12_, connection_1__12__11_, 
        connection_1__12__10_, connection_1__12__9_, connection_1__12__8_, 
        connection_1__12__7_, connection_1__12__6_, connection_1__12__5_, 
        connection_1__12__4_, connection_1__12__3_, connection_1__12__2_, 
        connection_1__12__1_, connection_1__12__0_}), .i_fwd_valid(
        fwd_connection_valid_frist_half[9]), .i_fwd_data_bus(
        fwd_connection_frist_half[319:288]), .o_fwd_valid(
        fwd_connection_valid_frist_half[11]), .o_fwd_data_bus(
        fwd_connection_frist_half[383:352]), .i_en(n533), .i_cmd({
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__6__4_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__6__3_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__6__2_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__6__1_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__6__0_}) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_33 first_half_stages_1__sw_group_1__bottom_group_1__genblk1_bottom_sw ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_0__15_, 
        connection_valid_0__14_}), .i_data_bus({connection_0__15__31_, 
        connection_0__15__30_, connection_0__15__29_, connection_0__15__28_, 
        connection_0__15__27_, connection_0__15__26_, connection_0__15__25_, 
        connection_0__15__24_, connection_0__15__23_, connection_0__15__22_, 
        connection_0__15__21_, connection_0__15__20_, connection_0__15__19_, 
        connection_0__15__18_, connection_0__15__17_, connection_0__15__16_, 
        connection_0__15__15_, connection_0__15__14_, connection_0__15__13_, 
        connection_0__15__12_, connection_0__15__11_, connection_0__15__10_, 
        connection_0__15__9_, connection_0__15__8_, connection_0__15__7_, 
        connection_0__15__6_, connection_0__15__5_, connection_0__15__4_, 
        connection_0__15__3_, connection_0__15__2_, connection_0__15__1_, 
        connection_0__15__0_, connection_0__14__31_, connection_0__14__30_, 
        connection_0__14__29_, connection_0__14__28_, connection_0__14__27_, 
        connection_0__14__26_, connection_0__14__25_, connection_0__14__24_, 
        connection_0__14__23_, connection_0__14__22_, connection_0__14__21_, 
        connection_0__14__20_, connection_0__14__19_, connection_0__14__18_, 
        connection_0__14__17_, connection_0__14__16_, connection_0__14__15_, 
        connection_0__14__14_, connection_0__14__13_, connection_0__14__12_, 
        connection_0__14__11_, connection_0__14__10_, connection_0__14__9_, 
        connection_0__14__8_, connection_0__14__7_, connection_0__14__6_, 
        connection_0__14__5_, connection_0__14__4_, connection_0__14__3_, 
        connection_0__14__2_, connection_0__14__1_, connection_0__14__0_}), 
        .o_valid({connection_valid_1__15_, connection_valid_1__14_}), 
        .o_data_bus({connection_1__15__31_, connection_1__15__30_, 
        connection_1__15__29_, connection_1__15__28_, connection_1__15__27_, 
        connection_1__15__26_, connection_1__15__25_, connection_1__15__24_, 
        connection_1__15__23_, connection_1__15__22_, connection_1__15__21_, 
        connection_1__15__20_, connection_1__15__19_, connection_1__15__18_, 
        connection_1__15__17_, connection_1__15__16_, connection_1__15__15_, 
        connection_1__15__14_, connection_1__15__13_, connection_1__15__12_, 
        connection_1__15__11_, connection_1__15__10_, connection_1__15__9_, 
        connection_1__15__8_, connection_1__15__7_, connection_1__15__6_, 
        connection_1__15__5_, connection_1__15__4_, connection_1__15__3_, 
        connection_1__15__2_, connection_1__15__1_, connection_1__15__0_, 
        connection_1__14__31_, connection_1__14__30_, connection_1__14__29_, 
        connection_1__14__28_, connection_1__14__27_, connection_1__14__26_, 
        connection_1__14__25_, connection_1__14__24_, connection_1__14__23_, 
        connection_1__14__22_, connection_1__14__21_, connection_1__14__20_, 
        connection_1__14__19_, connection_1__14__18_, connection_1__14__17_, 
        connection_1__14__16_, connection_1__14__15_, connection_1__14__14_, 
        connection_1__14__13_, connection_1__14__12_, connection_1__14__11_, 
        connection_1__14__10_, connection_1__14__9_, connection_1__14__8_, 
        connection_1__14__7_, connection_1__14__6_, connection_1__14__5_, 
        connection_1__14__4_, connection_1__14__3_, connection_1__14__2_, 
        connection_1__14__1_, connection_1__14__0_}), .i_fwd_valid(
        fwd_connection_valid_frist_half[8]), .i_fwd_data_bus(
        fwd_connection_frist_half[287:256]), .o_fwd_valid(
        fwd_connection_valid_frist_half[10]), .o_fwd_data_bus(
        fwd_connection_frist_half[351:320]), .i_en(n533), .i_cmd({
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__7__4_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__7__3_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__7__2_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__7__1_, 
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__7__0_}) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_32 first_half_stages_2__sw_group_0__upper_group_0__genblk1_upper_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_1__1_, 
        connection_valid_1__0_}), .i_data_bus({connection_1__1__31_, 
        connection_1__1__30_, connection_1__1__29_, connection_1__1__28_, 
        connection_1__1__27_, connection_1__1__26_, connection_1__1__25_, 
        connection_1__1__24_, connection_1__1__23_, connection_1__1__22_, 
        connection_1__1__21_, connection_1__1__20_, connection_1__1__19_, 
        connection_1__1__18_, connection_1__1__17_, connection_1__1__16_, 
        connection_1__1__15_, connection_1__1__14_, connection_1__1__13_, 
        connection_1__1__12_, connection_1__1__11_, connection_1__1__10_, 
        connection_1__1__9_, connection_1__1__8_, connection_1__1__7_, 
        connection_1__1__6_, connection_1__1__5_, connection_1__1__4_, 
        connection_1__1__3_, connection_1__1__2_, connection_1__1__1_, 
        connection_1__1__0_, connection_1__0__31_, connection_1__0__30_, 
        connection_1__0__29_, connection_1__0__28_, connection_1__0__27_, 
        connection_1__0__26_, connection_1__0__25_, connection_1__0__24_, 
        connection_1__0__23_, connection_1__0__22_, connection_1__0__21_, 
        connection_1__0__20_, connection_1__0__19_, connection_1__0__18_, 
        connection_1__0__17_, connection_1__0__16_, connection_1__0__15_, 
        connection_1__0__14_, connection_1__0__13_, connection_1__0__12_, 
        connection_1__0__11_, connection_1__0__10_, connection_1__0__9_, 
        connection_1__0__8_, connection_1__0__7_, connection_1__0__6_, 
        connection_1__0__5_, connection_1__0__4_, connection_1__0__3_, 
        connection_1__0__2_, connection_1__0__1_, connection_1__0__0_}), 
        .o_valid({connection_valid_2__1_, connection_valid_2__0_}), 
        .o_data_bus({connection_2__1__31_, connection_2__1__30_, 
        connection_2__1__29_, connection_2__1__28_, connection_2__1__27_, 
        connection_2__1__26_, connection_2__1__25_, connection_2__1__24_, 
        connection_2__1__23_, connection_2__1__22_, connection_2__1__21_, 
        connection_2__1__20_, connection_2__1__19_, connection_2__1__18_, 
        connection_2__1__17_, connection_2__1__16_, connection_2__1__15_, 
        connection_2__1__14_, connection_2__1__13_, connection_2__1__12_, 
        connection_2__1__11_, connection_2__1__10_, connection_2__1__9_, 
        connection_2__1__8_, connection_2__1__7_, connection_2__1__6_, 
        connection_2__1__5_, connection_2__1__4_, connection_2__1__3_, 
        connection_2__1__2_, connection_2__1__1_, connection_2__1__0_, 
        connection_2__0__31_, connection_2__0__30_, connection_2__0__29_, 
        connection_2__0__28_, connection_2__0__27_, connection_2__0__26_, 
        connection_2__0__25_, connection_2__0__24_, connection_2__0__23_, 
        connection_2__0__22_, connection_2__0__21_, connection_2__0__20_, 
        connection_2__0__19_, connection_2__0__18_, connection_2__0__17_, 
        connection_2__0__16_, connection_2__0__15_, connection_2__0__14_, 
        connection_2__0__13_, connection_2__0__12_, connection_2__0__11_, 
        connection_2__0__10_, connection_2__0__9_, connection_2__0__8_, 
        connection_2__0__7_, connection_2__0__6_, connection_2__0__5_, 
        connection_2__0__4_, connection_2__0__3_, connection_2__0__2_, 
        connection_2__0__1_, connection_2__0__0_}), .i_fwd_valid(
        fwd_connection_valid_frist_half[7]), .i_fwd_data_bus(
        fwd_connection_frist_half[255:224]), .o_fwd_valid(
        fwd_connection_valid_frist_half[6]), .o_fwd_data_bus(
        fwd_connection_frist_half[223:192]), .i_en(n533), .i_cmd({
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__0__4_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__0__3_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__0__2_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__0__1_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__0__0_}) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_31 first_half_stages_2__sw_group_0__bottom_group_0__genblk1_bottom_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_1__3_, 
        connection_valid_1__2_}), .i_data_bus({connection_1__3__31_, 
        connection_1__3__30_, connection_1__3__29_, connection_1__3__28_, 
        connection_1__3__27_, connection_1__3__26_, connection_1__3__25_, 
        connection_1__3__24_, connection_1__3__23_, connection_1__3__22_, 
        connection_1__3__21_, connection_1__3__20_, connection_1__3__19_, 
        connection_1__3__18_, connection_1__3__17_, connection_1__3__16_, 
        connection_1__3__15_, connection_1__3__14_, connection_1__3__13_, 
        connection_1__3__12_, connection_1__3__11_, connection_1__3__10_, 
        connection_1__3__9_, connection_1__3__8_, connection_1__3__7_, 
        connection_1__3__6_, connection_1__3__5_, connection_1__3__4_, 
        connection_1__3__3_, connection_1__3__2_, connection_1__3__1_, 
        connection_1__3__0_, connection_1__2__31_, connection_1__2__30_, 
        connection_1__2__29_, connection_1__2__28_, connection_1__2__27_, 
        connection_1__2__26_, connection_1__2__25_, connection_1__2__24_, 
        connection_1__2__23_, connection_1__2__22_, connection_1__2__21_, 
        connection_1__2__20_, connection_1__2__19_, connection_1__2__18_, 
        connection_1__2__17_, connection_1__2__16_, connection_1__2__15_, 
        connection_1__2__14_, connection_1__2__13_, connection_1__2__12_, 
        connection_1__2__11_, connection_1__2__10_, connection_1__2__9_, 
        connection_1__2__8_, connection_1__2__7_, connection_1__2__6_, 
        connection_1__2__5_, connection_1__2__4_, connection_1__2__3_, 
        connection_1__2__2_, connection_1__2__1_, connection_1__2__0_}), 
        .o_valid({connection_valid_2__3_, connection_valid_2__2_}), 
        .o_data_bus({connection_2__3__31_, connection_2__3__30_, 
        connection_2__3__29_, connection_2__3__28_, connection_2__3__27_, 
        connection_2__3__26_, connection_2__3__25_, connection_2__3__24_, 
        connection_2__3__23_, connection_2__3__22_, connection_2__3__21_, 
        connection_2__3__20_, connection_2__3__19_, connection_2__3__18_, 
        connection_2__3__17_, connection_2__3__16_, connection_2__3__15_, 
        connection_2__3__14_, connection_2__3__13_, connection_2__3__12_, 
        connection_2__3__11_, connection_2__3__10_, connection_2__3__9_, 
        connection_2__3__8_, connection_2__3__7_, connection_2__3__6_, 
        connection_2__3__5_, connection_2__3__4_, connection_2__3__3_, 
        connection_2__3__2_, connection_2__3__1_, connection_2__3__0_, 
        connection_2__2__31_, connection_2__2__30_, connection_2__2__29_, 
        connection_2__2__28_, connection_2__2__27_, connection_2__2__26_, 
        connection_2__2__25_, connection_2__2__24_, connection_2__2__23_, 
        connection_2__2__22_, connection_2__2__21_, connection_2__2__20_, 
        connection_2__2__19_, connection_2__2__18_, connection_2__2__17_, 
        connection_2__2__16_, connection_2__2__15_, connection_2__2__14_, 
        connection_2__2__13_, connection_2__2__12_, connection_2__2__11_, 
        connection_2__2__10_, connection_2__2__9_, connection_2__2__8_, 
        connection_2__2__7_, connection_2__2__6_, connection_2__2__5_, 
        connection_2__2__4_, connection_2__2__3_, connection_2__2__2_, 
        connection_2__2__1_, connection_2__2__0_}), .i_fwd_valid(
        fwd_connection_valid_frist_half[6]), .i_fwd_data_bus(
        fwd_connection_frist_half[223:192]), .o_fwd_valid(
        fwd_connection_valid_frist_half[7]), .o_fwd_data_bus(
        fwd_connection_frist_half[255:224]), .i_en(n533), .i_cmd({
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__1__4_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__1__3_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__1__2_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__1__1_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__1__0_}) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_30 first_half_stages_2__sw_group_1__upper_group_0__genblk1_upper_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_1__5_, 
        connection_valid_1__4_}), .i_data_bus({connection_1__5__31_, 
        connection_1__5__30_, connection_1__5__29_, connection_1__5__28_, 
        connection_1__5__27_, connection_1__5__26_, connection_1__5__25_, 
        connection_1__5__24_, connection_1__5__23_, connection_1__5__22_, 
        connection_1__5__21_, connection_1__5__20_, connection_1__5__19_, 
        connection_1__5__18_, connection_1__5__17_, connection_1__5__16_, 
        connection_1__5__15_, connection_1__5__14_, connection_1__5__13_, 
        connection_1__5__12_, connection_1__5__11_, connection_1__5__10_, 
        connection_1__5__9_, connection_1__5__8_, connection_1__5__7_, 
        connection_1__5__6_, connection_1__5__5_, connection_1__5__4_, 
        connection_1__5__3_, connection_1__5__2_, connection_1__5__1_, 
        connection_1__5__0_, connection_1__4__31_, connection_1__4__30_, 
        connection_1__4__29_, connection_1__4__28_, connection_1__4__27_, 
        connection_1__4__26_, connection_1__4__25_, connection_1__4__24_, 
        connection_1__4__23_, connection_1__4__22_, connection_1__4__21_, 
        connection_1__4__20_, connection_1__4__19_, connection_1__4__18_, 
        connection_1__4__17_, connection_1__4__16_, connection_1__4__15_, 
        connection_1__4__14_, connection_1__4__13_, connection_1__4__12_, 
        connection_1__4__11_, connection_1__4__10_, connection_1__4__9_, 
        connection_1__4__8_, connection_1__4__7_, connection_1__4__6_, 
        connection_1__4__5_, connection_1__4__4_, connection_1__4__3_, 
        connection_1__4__2_, connection_1__4__1_, connection_1__4__0_}), 
        .o_valid({connection_valid_2__5_, connection_valid_2__4_}), 
        .o_data_bus({connection_2__5__31_, connection_2__5__30_, 
        connection_2__5__29_, connection_2__5__28_, connection_2__5__27_, 
        connection_2__5__26_, connection_2__5__25_, connection_2__5__24_, 
        connection_2__5__23_, connection_2__5__22_, connection_2__5__21_, 
        connection_2__5__20_, connection_2__5__19_, connection_2__5__18_, 
        connection_2__5__17_, connection_2__5__16_, connection_2__5__15_, 
        connection_2__5__14_, connection_2__5__13_, connection_2__5__12_, 
        connection_2__5__11_, connection_2__5__10_, connection_2__5__9_, 
        connection_2__5__8_, connection_2__5__7_, connection_2__5__6_, 
        connection_2__5__5_, connection_2__5__4_, connection_2__5__3_, 
        connection_2__5__2_, connection_2__5__1_, connection_2__5__0_, 
        connection_2__4__31_, connection_2__4__30_, connection_2__4__29_, 
        connection_2__4__28_, connection_2__4__27_, connection_2__4__26_, 
        connection_2__4__25_, connection_2__4__24_, connection_2__4__23_, 
        connection_2__4__22_, connection_2__4__21_, connection_2__4__20_, 
        connection_2__4__19_, connection_2__4__18_, connection_2__4__17_, 
        connection_2__4__16_, connection_2__4__15_, connection_2__4__14_, 
        connection_2__4__13_, connection_2__4__12_, connection_2__4__11_, 
        connection_2__4__10_, connection_2__4__9_, connection_2__4__8_, 
        connection_2__4__7_, connection_2__4__6_, connection_2__4__5_, 
        connection_2__4__4_, connection_2__4__3_, connection_2__4__2_, 
        connection_2__4__1_, connection_2__4__0_}), .i_fwd_valid(
        fwd_connection_valid_frist_half[5]), .i_fwd_data_bus(
        fwd_connection_frist_half[191:160]), .o_fwd_valid(
        fwd_connection_valid_frist_half[4]), .o_fwd_data_bus(
        fwd_connection_frist_half[159:128]), .i_en(n533), .i_cmd({
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__2__4_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__2__3_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__2__2_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__2__1_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__2__0_}) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_29 first_half_stages_2__sw_group_1__bottom_group_0__genblk1_bottom_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_1__7_, 
        connection_valid_1__6_}), .i_data_bus({connection_1__7__31_, 
        connection_1__7__30_, connection_1__7__29_, connection_1__7__28_, 
        connection_1__7__27_, connection_1__7__26_, connection_1__7__25_, 
        connection_1__7__24_, connection_1__7__23_, connection_1__7__22_, 
        connection_1__7__21_, connection_1__7__20_, connection_1__7__19_, 
        connection_1__7__18_, connection_1__7__17_, connection_1__7__16_, 
        connection_1__7__15_, connection_1__7__14_, connection_1__7__13_, 
        connection_1__7__12_, connection_1__7__11_, connection_1__7__10_, 
        connection_1__7__9_, connection_1__7__8_, connection_1__7__7_, 
        connection_1__7__6_, connection_1__7__5_, connection_1__7__4_, 
        connection_1__7__3_, connection_1__7__2_, connection_1__7__1_, 
        connection_1__7__0_, connection_1__6__31_, connection_1__6__30_, 
        connection_1__6__29_, connection_1__6__28_, connection_1__6__27_, 
        connection_1__6__26_, connection_1__6__25_, connection_1__6__24_, 
        connection_1__6__23_, connection_1__6__22_, connection_1__6__21_, 
        connection_1__6__20_, connection_1__6__19_, connection_1__6__18_, 
        connection_1__6__17_, connection_1__6__16_, connection_1__6__15_, 
        connection_1__6__14_, connection_1__6__13_, connection_1__6__12_, 
        connection_1__6__11_, connection_1__6__10_, connection_1__6__9_, 
        connection_1__6__8_, connection_1__6__7_, connection_1__6__6_, 
        connection_1__6__5_, connection_1__6__4_, connection_1__6__3_, 
        connection_1__6__2_, connection_1__6__1_, connection_1__6__0_}), 
        .o_valid({connection_valid_2__7_, connection_valid_2__6_}), 
        .o_data_bus({connection_2__7__31_, connection_2__7__30_, 
        connection_2__7__29_, connection_2__7__28_, connection_2__7__27_, 
        connection_2__7__26_, connection_2__7__25_, connection_2__7__24_, 
        connection_2__7__23_, connection_2__7__22_, connection_2__7__21_, 
        connection_2__7__20_, connection_2__7__19_, connection_2__7__18_, 
        connection_2__7__17_, connection_2__7__16_, connection_2__7__15_, 
        connection_2__7__14_, connection_2__7__13_, connection_2__7__12_, 
        connection_2__7__11_, connection_2__7__10_, connection_2__7__9_, 
        connection_2__7__8_, connection_2__7__7_, connection_2__7__6_, 
        connection_2__7__5_, connection_2__7__4_, connection_2__7__3_, 
        connection_2__7__2_, connection_2__7__1_, connection_2__7__0_, 
        connection_2__6__31_, connection_2__6__30_, connection_2__6__29_, 
        connection_2__6__28_, connection_2__6__27_, connection_2__6__26_, 
        connection_2__6__25_, connection_2__6__24_, connection_2__6__23_, 
        connection_2__6__22_, connection_2__6__21_, connection_2__6__20_, 
        connection_2__6__19_, connection_2__6__18_, connection_2__6__17_, 
        connection_2__6__16_, connection_2__6__15_, connection_2__6__14_, 
        connection_2__6__13_, connection_2__6__12_, connection_2__6__11_, 
        connection_2__6__10_, connection_2__6__9_, connection_2__6__8_, 
        connection_2__6__7_, connection_2__6__6_, connection_2__6__5_, 
        connection_2__6__4_, connection_2__6__3_, connection_2__6__2_, 
        connection_2__6__1_, connection_2__6__0_}), .i_fwd_valid(
        fwd_connection_valid_frist_half[4]), .i_fwd_data_bus(
        fwd_connection_frist_half[159:128]), .o_fwd_valid(
        fwd_connection_valid_frist_half[5]), .o_fwd_data_bus(
        fwd_connection_frist_half[191:160]), .i_en(n533), .i_cmd({
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__3__4_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__3__3_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__3__2_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__3__1_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__3__0_}) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_28 first_half_stages_2__sw_group_2__upper_group_0__genblk1_upper_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_1__9_, 
        connection_valid_1__8_}), .i_data_bus({connection_1__9__31_, 
        connection_1__9__30_, connection_1__9__29_, connection_1__9__28_, 
        connection_1__9__27_, connection_1__9__26_, connection_1__9__25_, 
        connection_1__9__24_, connection_1__9__23_, connection_1__9__22_, 
        connection_1__9__21_, connection_1__9__20_, connection_1__9__19_, 
        connection_1__9__18_, connection_1__9__17_, connection_1__9__16_, 
        connection_1__9__15_, connection_1__9__14_, connection_1__9__13_, 
        connection_1__9__12_, connection_1__9__11_, connection_1__9__10_, 
        connection_1__9__9_, connection_1__9__8_, connection_1__9__7_, 
        connection_1__9__6_, connection_1__9__5_, connection_1__9__4_, 
        connection_1__9__3_, connection_1__9__2_, connection_1__9__1_, 
        connection_1__9__0_, connection_1__8__31_, connection_1__8__30_, 
        connection_1__8__29_, connection_1__8__28_, connection_1__8__27_, 
        connection_1__8__26_, connection_1__8__25_, connection_1__8__24_, 
        connection_1__8__23_, connection_1__8__22_, connection_1__8__21_, 
        connection_1__8__20_, connection_1__8__19_, connection_1__8__18_, 
        connection_1__8__17_, connection_1__8__16_, connection_1__8__15_, 
        connection_1__8__14_, connection_1__8__13_, connection_1__8__12_, 
        connection_1__8__11_, connection_1__8__10_, connection_1__8__9_, 
        connection_1__8__8_, connection_1__8__7_, connection_1__8__6_, 
        connection_1__8__5_, connection_1__8__4_, connection_1__8__3_, 
        connection_1__8__2_, connection_1__8__1_, connection_1__8__0_}), 
        .o_valid({connection_valid_2__9_, connection_valid_2__8_}), 
        .o_data_bus({connection_2__9__31_, connection_2__9__30_, 
        connection_2__9__29_, connection_2__9__28_, connection_2__9__27_, 
        connection_2__9__26_, connection_2__9__25_, connection_2__9__24_, 
        connection_2__9__23_, connection_2__9__22_, connection_2__9__21_, 
        connection_2__9__20_, connection_2__9__19_, connection_2__9__18_, 
        connection_2__9__17_, connection_2__9__16_, connection_2__9__15_, 
        connection_2__9__14_, connection_2__9__13_, connection_2__9__12_, 
        connection_2__9__11_, connection_2__9__10_, connection_2__9__9_, 
        connection_2__9__8_, connection_2__9__7_, connection_2__9__6_, 
        connection_2__9__5_, connection_2__9__4_, connection_2__9__3_, 
        connection_2__9__2_, connection_2__9__1_, connection_2__9__0_, 
        connection_2__8__31_, connection_2__8__30_, connection_2__8__29_, 
        connection_2__8__28_, connection_2__8__27_, connection_2__8__26_, 
        connection_2__8__25_, connection_2__8__24_, connection_2__8__23_, 
        connection_2__8__22_, connection_2__8__21_, connection_2__8__20_, 
        connection_2__8__19_, connection_2__8__18_, connection_2__8__17_, 
        connection_2__8__16_, connection_2__8__15_, connection_2__8__14_, 
        connection_2__8__13_, connection_2__8__12_, connection_2__8__11_, 
        connection_2__8__10_, connection_2__8__9_, connection_2__8__8_, 
        connection_2__8__7_, connection_2__8__6_, connection_2__8__5_, 
        connection_2__8__4_, connection_2__8__3_, connection_2__8__2_, 
        connection_2__8__1_, connection_2__8__0_}), .i_fwd_valid(
        fwd_connection_valid_frist_half[3]), .i_fwd_data_bus(
        fwd_connection_frist_half[127:96]), .o_fwd_valid(
        fwd_connection_valid_frist_half[2]), .o_fwd_data_bus(
        fwd_connection_frist_half[95:64]), .i_en(n533), .i_cmd({
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__4__4_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__4__3_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__4__2_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__4__1_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__4__0_}) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_27 first_half_stages_2__sw_group_2__bottom_group_0__genblk1_bottom_sw ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_1__11_, 
        connection_valid_1__10_}), .i_data_bus({connection_1__11__31_, 
        connection_1__11__30_, connection_1__11__29_, connection_1__11__28_, 
        connection_1__11__27_, connection_1__11__26_, connection_1__11__25_, 
        connection_1__11__24_, connection_1__11__23_, connection_1__11__22_, 
        connection_1__11__21_, connection_1__11__20_, connection_1__11__19_, 
        connection_1__11__18_, connection_1__11__17_, connection_1__11__16_, 
        connection_1__11__15_, connection_1__11__14_, connection_1__11__13_, 
        connection_1__11__12_, connection_1__11__11_, connection_1__11__10_, 
        connection_1__11__9_, connection_1__11__8_, connection_1__11__7_, 
        connection_1__11__6_, connection_1__11__5_, connection_1__11__4_, 
        connection_1__11__3_, connection_1__11__2_, connection_1__11__1_, 
        connection_1__11__0_, connection_1__10__31_, connection_1__10__30_, 
        connection_1__10__29_, connection_1__10__28_, connection_1__10__27_, 
        connection_1__10__26_, connection_1__10__25_, connection_1__10__24_, 
        connection_1__10__23_, connection_1__10__22_, connection_1__10__21_, 
        connection_1__10__20_, connection_1__10__19_, connection_1__10__18_, 
        connection_1__10__17_, connection_1__10__16_, connection_1__10__15_, 
        connection_1__10__14_, connection_1__10__13_, connection_1__10__12_, 
        connection_1__10__11_, connection_1__10__10_, connection_1__10__9_, 
        connection_1__10__8_, connection_1__10__7_, connection_1__10__6_, 
        connection_1__10__5_, connection_1__10__4_, connection_1__10__3_, 
        connection_1__10__2_, connection_1__10__1_, connection_1__10__0_}), 
        .o_valid({connection_valid_2__11_, connection_valid_2__10_}), 
        .o_data_bus({connection_2__11__31_, connection_2__11__30_, 
        connection_2__11__29_, connection_2__11__28_, connection_2__11__27_, 
        connection_2__11__26_, connection_2__11__25_, connection_2__11__24_, 
        connection_2__11__23_, connection_2__11__22_, connection_2__11__21_, 
        connection_2__11__20_, connection_2__11__19_, connection_2__11__18_, 
        connection_2__11__17_, connection_2__11__16_, connection_2__11__15_, 
        connection_2__11__14_, connection_2__11__13_, connection_2__11__12_, 
        connection_2__11__11_, connection_2__11__10_, connection_2__11__9_, 
        connection_2__11__8_, connection_2__11__7_, connection_2__11__6_, 
        connection_2__11__5_, connection_2__11__4_, connection_2__11__3_, 
        connection_2__11__2_, connection_2__11__1_, connection_2__11__0_, 
        connection_2__10__31_, connection_2__10__30_, connection_2__10__29_, 
        connection_2__10__28_, connection_2__10__27_, connection_2__10__26_, 
        connection_2__10__25_, connection_2__10__24_, connection_2__10__23_, 
        connection_2__10__22_, connection_2__10__21_, connection_2__10__20_, 
        connection_2__10__19_, connection_2__10__18_, connection_2__10__17_, 
        connection_2__10__16_, connection_2__10__15_, connection_2__10__14_, 
        connection_2__10__13_, connection_2__10__12_, connection_2__10__11_, 
        connection_2__10__10_, connection_2__10__9_, connection_2__10__8_, 
        connection_2__10__7_, connection_2__10__6_, connection_2__10__5_, 
        connection_2__10__4_, connection_2__10__3_, connection_2__10__2_, 
        connection_2__10__1_, connection_2__10__0_}), .i_fwd_valid(
        fwd_connection_valid_frist_half[2]), .i_fwd_data_bus(
        fwd_connection_frist_half[95:64]), .o_fwd_valid(
        fwd_connection_valid_frist_half[3]), .o_fwd_data_bus(
        fwd_connection_frist_half[127:96]), .i_en(n533), .i_cmd({
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__5__4_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__5__3_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__5__2_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__5__1_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__5__0_}) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_26 first_half_stages_2__sw_group_3__upper_group_0__genblk1_upper_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_1__13_, 
        connection_valid_1__12_}), .i_data_bus({connection_1__13__31_, 
        connection_1__13__30_, connection_1__13__29_, connection_1__13__28_, 
        connection_1__13__27_, connection_1__13__26_, connection_1__13__25_, 
        connection_1__13__24_, connection_1__13__23_, connection_1__13__22_, 
        connection_1__13__21_, connection_1__13__20_, connection_1__13__19_, 
        connection_1__13__18_, connection_1__13__17_, connection_1__13__16_, 
        connection_1__13__15_, connection_1__13__14_, connection_1__13__13_, 
        connection_1__13__12_, connection_1__13__11_, connection_1__13__10_, 
        connection_1__13__9_, connection_1__13__8_, connection_1__13__7_, 
        connection_1__13__6_, connection_1__13__5_, connection_1__13__4_, 
        connection_1__13__3_, connection_1__13__2_, connection_1__13__1_, 
        connection_1__13__0_, connection_1__12__31_, connection_1__12__30_, 
        connection_1__12__29_, connection_1__12__28_, connection_1__12__27_, 
        connection_1__12__26_, connection_1__12__25_, connection_1__12__24_, 
        connection_1__12__23_, connection_1__12__22_, connection_1__12__21_, 
        connection_1__12__20_, connection_1__12__19_, connection_1__12__18_, 
        connection_1__12__17_, connection_1__12__16_, connection_1__12__15_, 
        connection_1__12__14_, connection_1__12__13_, connection_1__12__12_, 
        connection_1__12__11_, connection_1__12__10_, connection_1__12__9_, 
        connection_1__12__8_, connection_1__12__7_, connection_1__12__6_, 
        connection_1__12__5_, connection_1__12__4_, connection_1__12__3_, 
        connection_1__12__2_, connection_1__12__1_, connection_1__12__0_}), 
        .o_valid({connection_valid_2__13_, connection_valid_2__12_}), 
        .o_data_bus({connection_2__13__31_, connection_2__13__30_, 
        connection_2__13__29_, connection_2__13__28_, connection_2__13__27_, 
        connection_2__13__26_, connection_2__13__25_, connection_2__13__24_, 
        connection_2__13__23_, connection_2__13__22_, connection_2__13__21_, 
        connection_2__13__20_, connection_2__13__19_, connection_2__13__18_, 
        connection_2__13__17_, connection_2__13__16_, connection_2__13__15_, 
        connection_2__13__14_, connection_2__13__13_, connection_2__13__12_, 
        connection_2__13__11_, connection_2__13__10_, connection_2__13__9_, 
        connection_2__13__8_, connection_2__13__7_, connection_2__13__6_, 
        connection_2__13__5_, connection_2__13__4_, connection_2__13__3_, 
        connection_2__13__2_, connection_2__13__1_, connection_2__13__0_, 
        connection_2__12__31_, connection_2__12__30_, connection_2__12__29_, 
        connection_2__12__28_, connection_2__12__27_, connection_2__12__26_, 
        connection_2__12__25_, connection_2__12__24_, connection_2__12__23_, 
        connection_2__12__22_, connection_2__12__21_, connection_2__12__20_, 
        connection_2__12__19_, connection_2__12__18_, connection_2__12__17_, 
        connection_2__12__16_, connection_2__12__15_, connection_2__12__14_, 
        connection_2__12__13_, connection_2__12__12_, connection_2__12__11_, 
        connection_2__12__10_, connection_2__12__9_, connection_2__12__8_, 
        connection_2__12__7_, connection_2__12__6_, connection_2__12__5_, 
        connection_2__12__4_, connection_2__12__3_, connection_2__12__2_, 
        connection_2__12__1_, connection_2__12__0_}), .i_fwd_valid(
        fwd_connection_valid_frist_half[1]), .i_fwd_data_bus(
        fwd_connection_frist_half[63:32]), .o_fwd_valid(
        fwd_connection_valid_frist_half[0]), .o_fwd_data_bus(
        fwd_connection_frist_half[31:0]), .i_en(n533), .i_cmd({
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__6__4_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__6__3_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__6__2_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__6__1_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__6__0_}) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_25 first_half_stages_2__sw_group_3__bottom_group_0__genblk1_bottom_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_1__15_, 
        connection_valid_1__14_}), .i_data_bus({connection_1__15__31_, 
        connection_1__15__30_, connection_1__15__29_, connection_1__15__28_, 
        connection_1__15__27_, connection_1__15__26_, connection_1__15__25_, 
        connection_1__15__24_, connection_1__15__23_, connection_1__15__22_, 
        connection_1__15__21_, connection_1__15__20_, connection_1__15__19_, 
        connection_1__15__18_, connection_1__15__17_, connection_1__15__16_, 
        connection_1__15__15_, connection_1__15__14_, connection_1__15__13_, 
        connection_1__15__12_, connection_1__15__11_, connection_1__15__10_, 
        connection_1__15__9_, connection_1__15__8_, connection_1__15__7_, 
        connection_1__15__6_, connection_1__15__5_, connection_1__15__4_, 
        connection_1__15__3_, connection_1__15__2_, connection_1__15__1_, 
        connection_1__15__0_, connection_1__14__31_, connection_1__14__30_, 
        connection_1__14__29_, connection_1__14__28_, connection_1__14__27_, 
        connection_1__14__26_, connection_1__14__25_, connection_1__14__24_, 
        connection_1__14__23_, connection_1__14__22_, connection_1__14__21_, 
        connection_1__14__20_, connection_1__14__19_, connection_1__14__18_, 
        connection_1__14__17_, connection_1__14__16_, connection_1__14__15_, 
        connection_1__14__14_, connection_1__14__13_, connection_1__14__12_, 
        connection_1__14__11_, connection_1__14__10_, connection_1__14__9_, 
        connection_1__14__8_, connection_1__14__7_, connection_1__14__6_, 
        connection_1__14__5_, connection_1__14__4_, connection_1__14__3_, 
        connection_1__14__2_, connection_1__14__1_, connection_1__14__0_}), 
        .o_valid({connection_valid_2__15_, connection_valid_2__14_}), 
        .o_data_bus({connection_2__15__31_, connection_2__15__30_, 
        connection_2__15__29_, connection_2__15__28_, connection_2__15__27_, 
        connection_2__15__26_, connection_2__15__25_, connection_2__15__24_, 
        connection_2__15__23_, connection_2__15__22_, connection_2__15__21_, 
        connection_2__15__20_, connection_2__15__19_, connection_2__15__18_, 
        connection_2__15__17_, connection_2__15__16_, connection_2__15__15_, 
        connection_2__15__14_, connection_2__15__13_, connection_2__15__12_, 
        connection_2__15__11_, connection_2__15__10_, connection_2__15__9_, 
        connection_2__15__8_, connection_2__15__7_, connection_2__15__6_, 
        connection_2__15__5_, connection_2__15__4_, connection_2__15__3_, 
        connection_2__15__2_, connection_2__15__1_, connection_2__15__0_, 
        connection_2__14__31_, connection_2__14__30_, connection_2__14__29_, 
        connection_2__14__28_, connection_2__14__27_, connection_2__14__26_, 
        connection_2__14__25_, connection_2__14__24_, connection_2__14__23_, 
        connection_2__14__22_, connection_2__14__21_, connection_2__14__20_, 
        connection_2__14__19_, connection_2__14__18_, connection_2__14__17_, 
        connection_2__14__16_, connection_2__14__15_, connection_2__14__14_, 
        connection_2__14__13_, connection_2__14__12_, connection_2__14__11_, 
        connection_2__14__10_, connection_2__14__9_, connection_2__14__8_, 
        connection_2__14__7_, connection_2__14__6_, connection_2__14__5_, 
        connection_2__14__4_, connection_2__14__3_, connection_2__14__2_, 
        connection_2__14__1_, connection_2__14__0_}), .i_fwd_valid(
        fwd_connection_valid_frist_half[0]), .i_fwd_data_bus(
        fwd_connection_frist_half[31:0]), .o_fwd_valid(
        fwd_connection_valid_frist_half[1]), .o_fwd_data_bus(
        fwd_connection_frist_half[63:32]), .i_en(n533), .i_cmd({
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__7__4_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__7__3_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__7__2_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__7__1_, 
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__7__0_}) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_0 middle_stage_0__middle_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__1_, 
        connection_valid_2__0_}), .i_data_bus({connection_2__1__31_, 
        connection_2__1__30_, connection_2__1__29_, connection_2__1__28_, 
        connection_2__1__27_, connection_2__1__26_, connection_2__1__25_, 
        connection_2__1__24_, connection_2__1__23_, connection_2__1__22_, 
        connection_2__1__21_, connection_2__1__20_, connection_2__1__19_, 
        connection_2__1__18_, connection_2__1__17_, connection_2__1__16_, 
        connection_2__1__15_, connection_2__1__14_, connection_2__1__13_, 
        connection_2__1__12_, connection_2__1__11_, connection_2__1__10_, 
        connection_2__1__9_, connection_2__1__8_, connection_2__1__7_, 
        connection_2__1__6_, connection_2__1__5_, connection_2__1__4_, 
        connection_2__1__3_, connection_2__1__2_, connection_2__1__1_, 
        connection_2__1__0_, connection_2__0__31_, connection_2__0__30_, 
        connection_2__0__29_, connection_2__0__28_, connection_2__0__27_, 
        connection_2__0__26_, connection_2__0__25_, connection_2__0__24_, 
        connection_2__0__23_, connection_2__0__22_, connection_2__0__21_, 
        connection_2__0__20_, connection_2__0__19_, connection_2__0__18_, 
        connection_2__0__17_, connection_2__0__16_, connection_2__0__15_, 
        connection_2__0__14_, connection_2__0__13_, connection_2__0__12_, 
        connection_2__0__11_, connection_2__0__10_, connection_2__0__9_, 
        connection_2__0__8_, connection_2__0__7_, connection_2__0__6_, 
        connection_2__0__5_, connection_2__0__4_, connection_2__0__3_, 
        connection_2__0__2_, connection_2__0__1_, connection_2__0__0_}), 
        .o_valid({connection_valid_3__1_, connection_valid_3__0_}), 
        .o_data_bus({connection_3__1__31_, connection_3__1__30_, 
        connection_3__1__29_, connection_3__1__28_, connection_3__1__27_, 
        connection_3__1__26_, connection_3__1__25_, connection_3__1__24_, 
        connection_3__1__23_, connection_3__1__22_, connection_3__1__21_, 
        connection_3__1__20_, connection_3__1__19_, connection_3__1__18_, 
        connection_3__1__17_, connection_3__1__16_, connection_3__1__15_, 
        connection_3__1__14_, connection_3__1__13_, connection_3__1__12_, 
        connection_3__1__11_, connection_3__1__10_, connection_3__1__9_, 
        connection_3__1__8_, connection_3__1__7_, connection_3__1__6_, 
        connection_3__1__5_, connection_3__1__4_, connection_3__1__3_, 
        connection_3__1__2_, connection_3__1__1_, connection_3__1__0_, 
        connection_3__0__31_, connection_3__0__30_, connection_3__0__29_, 
        connection_3__0__28_, connection_3__0__27_, connection_3__0__26_, 
        connection_3__0__25_, connection_3__0__24_, connection_3__0__23_, 
        connection_3__0__22_, connection_3__0__21_, connection_3__0__20_, 
        connection_3__0__19_, connection_3__0__18_, connection_3__0__17_, 
        connection_3__0__16_, connection_3__0__15_, connection_3__0__14_, 
        connection_3__0__13_, connection_3__0__12_, connection_3__0__11_, 
        connection_3__0__10_, connection_3__0__9_, connection_3__0__8_, 
        connection_3__0__7_, connection_3__0__6_, connection_3__0__5_, 
        connection_3__0__4_, connection_3__0__3_, connection_3__0__2_, 
        connection_3__0__1_, connection_3__0__0_}), .i_en(i_en), .i_cmd({
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__0__1_, 
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__0__0_}) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_7 middle_stage_1__middle_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__3_, 
        connection_valid_2__2_}), .i_data_bus({connection_2__3__31_, 
        connection_2__3__30_, connection_2__3__29_, connection_2__3__28_, 
        connection_2__3__27_, connection_2__3__26_, connection_2__3__25_, 
        connection_2__3__24_, connection_2__3__23_, connection_2__3__22_, 
        connection_2__3__21_, connection_2__3__20_, connection_2__3__19_, 
        connection_2__3__18_, connection_2__3__17_, connection_2__3__16_, 
        connection_2__3__15_, connection_2__3__14_, connection_2__3__13_, 
        connection_2__3__12_, connection_2__3__11_, connection_2__3__10_, 
        connection_2__3__9_, connection_2__3__8_, connection_2__3__7_, 
        connection_2__3__6_, connection_2__3__5_, connection_2__3__4_, 
        connection_2__3__3_, connection_2__3__2_, connection_2__3__1_, 
        connection_2__3__0_, connection_2__2__31_, connection_2__2__30_, 
        connection_2__2__29_, connection_2__2__28_, connection_2__2__27_, 
        connection_2__2__26_, connection_2__2__25_, connection_2__2__24_, 
        connection_2__2__23_, connection_2__2__22_, connection_2__2__21_, 
        connection_2__2__20_, connection_2__2__19_, connection_2__2__18_, 
        connection_2__2__17_, connection_2__2__16_, connection_2__2__15_, 
        connection_2__2__14_, connection_2__2__13_, connection_2__2__12_, 
        connection_2__2__11_, connection_2__2__10_, connection_2__2__9_, 
        connection_2__2__8_, connection_2__2__7_, connection_2__2__6_, 
        connection_2__2__5_, connection_2__2__4_, connection_2__2__3_, 
        connection_2__2__2_, connection_2__2__1_, connection_2__2__0_}), 
        .o_valid({connection_valid_3__3_, connection_valid_3__2_}), 
        .o_data_bus({connection_3__3__31_, connection_3__3__30_, 
        connection_3__3__29_, connection_3__3__28_, connection_3__3__27_, 
        connection_3__3__26_, connection_3__3__25_, connection_3__3__24_, 
        connection_3__3__23_, connection_3__3__22_, connection_3__3__21_, 
        connection_3__3__20_, connection_3__3__19_, connection_3__3__18_, 
        connection_3__3__17_, connection_3__3__16_, connection_3__3__15_, 
        connection_3__3__14_, connection_3__3__13_, connection_3__3__12_, 
        connection_3__3__11_, connection_3__3__10_, connection_3__3__9_, 
        connection_3__3__8_, connection_3__3__7_, connection_3__3__6_, 
        connection_3__3__5_, connection_3__3__4_, connection_3__3__3_, 
        connection_3__3__2_, connection_3__3__1_, connection_3__3__0_, 
        connection_3__2__31_, connection_3__2__30_, connection_3__2__29_, 
        connection_3__2__28_, connection_3__2__27_, connection_3__2__26_, 
        connection_3__2__25_, connection_3__2__24_, connection_3__2__23_, 
        connection_3__2__22_, connection_3__2__21_, connection_3__2__20_, 
        connection_3__2__19_, connection_3__2__18_, connection_3__2__17_, 
        connection_3__2__16_, connection_3__2__15_, connection_3__2__14_, 
        connection_3__2__13_, connection_3__2__12_, connection_3__2__11_, 
        connection_3__2__10_, connection_3__2__9_, connection_3__2__8_, 
        connection_3__2__7_, connection_3__2__6_, connection_3__2__5_, 
        connection_3__2__4_, connection_3__2__3_, connection_3__2__2_, 
        connection_3__2__1_, connection_3__2__0_}), .i_en(n533), .i_cmd({
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__1__1_, 
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__1__0_}) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_6 middle_stage_2__middle_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__5_, 
        connection_valid_2__4_}), .i_data_bus({connection_2__5__31_, 
        connection_2__5__30_, connection_2__5__29_, connection_2__5__28_, 
        connection_2__5__27_, connection_2__5__26_, connection_2__5__25_, 
        connection_2__5__24_, connection_2__5__23_, connection_2__5__22_, 
        connection_2__5__21_, connection_2__5__20_, connection_2__5__19_, 
        connection_2__5__18_, connection_2__5__17_, connection_2__5__16_, 
        connection_2__5__15_, connection_2__5__14_, connection_2__5__13_, 
        connection_2__5__12_, connection_2__5__11_, connection_2__5__10_, 
        connection_2__5__9_, connection_2__5__8_, connection_2__5__7_, 
        connection_2__5__6_, connection_2__5__5_, connection_2__5__4_, 
        connection_2__5__3_, connection_2__5__2_, connection_2__5__1_, 
        connection_2__5__0_, connection_2__4__31_, connection_2__4__30_, 
        connection_2__4__29_, connection_2__4__28_, connection_2__4__27_, 
        connection_2__4__26_, connection_2__4__25_, connection_2__4__24_, 
        connection_2__4__23_, connection_2__4__22_, connection_2__4__21_, 
        connection_2__4__20_, connection_2__4__19_, connection_2__4__18_, 
        connection_2__4__17_, connection_2__4__16_, connection_2__4__15_, 
        connection_2__4__14_, connection_2__4__13_, connection_2__4__12_, 
        connection_2__4__11_, connection_2__4__10_, connection_2__4__9_, 
        connection_2__4__8_, connection_2__4__7_, connection_2__4__6_, 
        connection_2__4__5_, connection_2__4__4_, connection_2__4__3_, 
        connection_2__4__2_, connection_2__4__1_, connection_2__4__0_}), 
        .o_valid({connection_valid_3__5_, connection_valid_3__4_}), 
        .o_data_bus({connection_3__5__31_, connection_3__5__30_, 
        connection_3__5__29_, connection_3__5__28_, connection_3__5__27_, 
        connection_3__5__26_, connection_3__5__25_, connection_3__5__24_, 
        connection_3__5__23_, connection_3__5__22_, connection_3__5__21_, 
        connection_3__5__20_, connection_3__5__19_, connection_3__5__18_, 
        connection_3__5__17_, connection_3__5__16_, connection_3__5__15_, 
        connection_3__5__14_, connection_3__5__13_, connection_3__5__12_, 
        connection_3__5__11_, connection_3__5__10_, connection_3__5__9_, 
        connection_3__5__8_, connection_3__5__7_, connection_3__5__6_, 
        connection_3__5__5_, connection_3__5__4_, connection_3__5__3_, 
        connection_3__5__2_, connection_3__5__1_, connection_3__5__0_, 
        connection_3__4__31_, connection_3__4__30_, connection_3__4__29_, 
        connection_3__4__28_, connection_3__4__27_, connection_3__4__26_, 
        connection_3__4__25_, connection_3__4__24_, connection_3__4__23_, 
        connection_3__4__22_, connection_3__4__21_, connection_3__4__20_, 
        connection_3__4__19_, connection_3__4__18_, connection_3__4__17_, 
        connection_3__4__16_, connection_3__4__15_, connection_3__4__14_, 
        connection_3__4__13_, connection_3__4__12_, connection_3__4__11_, 
        connection_3__4__10_, connection_3__4__9_, connection_3__4__8_, 
        connection_3__4__7_, connection_3__4__6_, connection_3__4__5_, 
        connection_3__4__4_, connection_3__4__3_, connection_3__4__2_, 
        connection_3__4__1_, connection_3__4__0_}), .i_en(i_en), .i_cmd({
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__2__1_, 
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__2__0_}) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_5 middle_stage_3__middle_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__7_, 
        connection_valid_2__6_}), .i_data_bus({connection_2__7__31_, 
        connection_2__7__30_, connection_2__7__29_, connection_2__7__28_, 
        connection_2__7__27_, connection_2__7__26_, connection_2__7__25_, 
        connection_2__7__24_, connection_2__7__23_, connection_2__7__22_, 
        connection_2__7__21_, connection_2__7__20_, connection_2__7__19_, 
        connection_2__7__18_, connection_2__7__17_, connection_2__7__16_, 
        connection_2__7__15_, connection_2__7__14_, connection_2__7__13_, 
        connection_2__7__12_, connection_2__7__11_, connection_2__7__10_, 
        connection_2__7__9_, connection_2__7__8_, connection_2__7__7_, 
        connection_2__7__6_, connection_2__7__5_, connection_2__7__4_, 
        connection_2__7__3_, connection_2__7__2_, connection_2__7__1_, 
        connection_2__7__0_, connection_2__6__31_, connection_2__6__30_, 
        connection_2__6__29_, connection_2__6__28_, connection_2__6__27_, 
        connection_2__6__26_, connection_2__6__25_, connection_2__6__24_, 
        connection_2__6__23_, connection_2__6__22_, connection_2__6__21_, 
        connection_2__6__20_, connection_2__6__19_, connection_2__6__18_, 
        connection_2__6__17_, connection_2__6__16_, connection_2__6__15_, 
        connection_2__6__14_, connection_2__6__13_, connection_2__6__12_, 
        connection_2__6__11_, connection_2__6__10_, connection_2__6__9_, 
        connection_2__6__8_, connection_2__6__7_, connection_2__6__6_, 
        connection_2__6__5_, connection_2__6__4_, connection_2__6__3_, 
        connection_2__6__2_, connection_2__6__1_, connection_2__6__0_}), 
        .o_valid({connection_valid_3__7_, connection_valid_3__6_}), 
        .o_data_bus({connection_3__7__31_, connection_3__7__30_, 
        connection_3__7__29_, connection_3__7__28_, connection_3__7__27_, 
        connection_3__7__26_, connection_3__7__25_, connection_3__7__24_, 
        connection_3__7__23_, connection_3__7__22_, connection_3__7__21_, 
        connection_3__7__20_, connection_3__7__19_, connection_3__7__18_, 
        connection_3__7__17_, connection_3__7__16_, connection_3__7__15_, 
        connection_3__7__14_, connection_3__7__13_, connection_3__7__12_, 
        connection_3__7__11_, connection_3__7__10_, connection_3__7__9_, 
        connection_3__7__8_, connection_3__7__7_, connection_3__7__6_, 
        connection_3__7__5_, connection_3__7__4_, connection_3__7__3_, 
        connection_3__7__2_, connection_3__7__1_, connection_3__7__0_, 
        connection_3__6__31_, connection_3__6__30_, connection_3__6__29_, 
        connection_3__6__28_, connection_3__6__27_, connection_3__6__26_, 
        connection_3__6__25_, connection_3__6__24_, connection_3__6__23_, 
        connection_3__6__22_, connection_3__6__21_, connection_3__6__20_, 
        connection_3__6__19_, connection_3__6__18_, connection_3__6__17_, 
        connection_3__6__16_, connection_3__6__15_, connection_3__6__14_, 
        connection_3__6__13_, connection_3__6__12_, connection_3__6__11_, 
        connection_3__6__10_, connection_3__6__9_, connection_3__6__8_, 
        connection_3__6__7_, connection_3__6__6_, connection_3__6__5_, 
        connection_3__6__4_, connection_3__6__3_, connection_3__6__2_, 
        connection_3__6__1_, connection_3__6__0_}), .i_en(i_en), .i_cmd({
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__3__1_, 
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__3__0_}) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_4 middle_stage_4__middle_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__9_, 
        connection_valid_2__8_}), .i_data_bus({connection_2__9__31_, 
        connection_2__9__30_, connection_2__9__29_, connection_2__9__28_, 
        connection_2__9__27_, connection_2__9__26_, connection_2__9__25_, 
        connection_2__9__24_, connection_2__9__23_, connection_2__9__22_, 
        connection_2__9__21_, connection_2__9__20_, connection_2__9__19_, 
        connection_2__9__18_, connection_2__9__17_, connection_2__9__16_, 
        connection_2__9__15_, connection_2__9__14_, connection_2__9__13_, 
        connection_2__9__12_, connection_2__9__11_, connection_2__9__10_, 
        connection_2__9__9_, connection_2__9__8_, connection_2__9__7_, 
        connection_2__9__6_, connection_2__9__5_, connection_2__9__4_, 
        connection_2__9__3_, connection_2__9__2_, connection_2__9__1_, 
        connection_2__9__0_, connection_2__8__31_, connection_2__8__30_, 
        connection_2__8__29_, connection_2__8__28_, connection_2__8__27_, 
        connection_2__8__26_, connection_2__8__25_, connection_2__8__24_, 
        connection_2__8__23_, connection_2__8__22_, connection_2__8__21_, 
        connection_2__8__20_, connection_2__8__19_, connection_2__8__18_, 
        connection_2__8__17_, connection_2__8__16_, connection_2__8__15_, 
        connection_2__8__14_, connection_2__8__13_, connection_2__8__12_, 
        connection_2__8__11_, connection_2__8__10_, connection_2__8__9_, 
        connection_2__8__8_, connection_2__8__7_, connection_2__8__6_, 
        connection_2__8__5_, connection_2__8__4_, connection_2__8__3_, 
        connection_2__8__2_, connection_2__8__1_, connection_2__8__0_}), 
        .o_valid({connection_valid_3__9_, connection_valid_3__8_}), 
        .o_data_bus({connection_3__9__31_, connection_3__9__30_, 
        connection_3__9__29_, connection_3__9__28_, connection_3__9__27_, 
        connection_3__9__26_, connection_3__9__25_, connection_3__9__24_, 
        connection_3__9__23_, connection_3__9__22_, connection_3__9__21_, 
        connection_3__9__20_, connection_3__9__19_, connection_3__9__18_, 
        connection_3__9__17_, connection_3__9__16_, connection_3__9__15_, 
        connection_3__9__14_, connection_3__9__13_, connection_3__9__12_, 
        connection_3__9__11_, connection_3__9__10_, connection_3__9__9_, 
        connection_3__9__8_, connection_3__9__7_, connection_3__9__6_, 
        connection_3__9__5_, connection_3__9__4_, connection_3__9__3_, 
        connection_3__9__2_, connection_3__9__1_, connection_3__9__0_, 
        connection_3__8__31_, connection_3__8__30_, connection_3__8__29_, 
        connection_3__8__28_, connection_3__8__27_, connection_3__8__26_, 
        connection_3__8__25_, connection_3__8__24_, connection_3__8__23_, 
        connection_3__8__22_, connection_3__8__21_, connection_3__8__20_, 
        connection_3__8__19_, connection_3__8__18_, connection_3__8__17_, 
        connection_3__8__16_, connection_3__8__15_, connection_3__8__14_, 
        connection_3__8__13_, connection_3__8__12_, connection_3__8__11_, 
        connection_3__8__10_, connection_3__8__9_, connection_3__8__8_, 
        connection_3__8__7_, connection_3__8__6_, connection_3__8__5_, 
        connection_3__8__4_, connection_3__8__3_, connection_3__8__2_, 
        connection_3__8__1_, connection_3__8__0_}), .i_en(i_en), .i_cmd({
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__4__1_, 
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__4__0_}) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_3 middle_stage_5__middle_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__11_, 
        connection_valid_2__10_}), .i_data_bus({connection_2__11__31_, 
        connection_2__11__30_, connection_2__11__29_, connection_2__11__28_, 
        connection_2__11__27_, connection_2__11__26_, connection_2__11__25_, 
        connection_2__11__24_, connection_2__11__23_, connection_2__11__22_, 
        connection_2__11__21_, connection_2__11__20_, connection_2__11__19_, 
        connection_2__11__18_, connection_2__11__17_, connection_2__11__16_, 
        connection_2__11__15_, connection_2__11__14_, connection_2__11__13_, 
        connection_2__11__12_, connection_2__11__11_, connection_2__11__10_, 
        connection_2__11__9_, connection_2__11__8_, connection_2__11__7_, 
        connection_2__11__6_, connection_2__11__5_, connection_2__11__4_, 
        connection_2__11__3_, connection_2__11__2_, connection_2__11__1_, 
        connection_2__11__0_, connection_2__10__31_, connection_2__10__30_, 
        connection_2__10__29_, connection_2__10__28_, connection_2__10__27_, 
        connection_2__10__26_, connection_2__10__25_, connection_2__10__24_, 
        connection_2__10__23_, connection_2__10__22_, connection_2__10__21_, 
        connection_2__10__20_, connection_2__10__19_, connection_2__10__18_, 
        connection_2__10__17_, connection_2__10__16_, connection_2__10__15_, 
        connection_2__10__14_, connection_2__10__13_, connection_2__10__12_, 
        connection_2__10__11_, connection_2__10__10_, connection_2__10__9_, 
        connection_2__10__8_, connection_2__10__7_, connection_2__10__6_, 
        connection_2__10__5_, connection_2__10__4_, connection_2__10__3_, 
        connection_2__10__2_, connection_2__10__1_, connection_2__10__0_}), 
        .o_valid({connection_valid_3__11_, connection_valid_3__10_}), 
        .o_data_bus({connection_3__11__31_, connection_3__11__30_, 
        connection_3__11__29_, connection_3__11__28_, connection_3__11__27_, 
        connection_3__11__26_, connection_3__11__25_, connection_3__11__24_, 
        connection_3__11__23_, connection_3__11__22_, connection_3__11__21_, 
        connection_3__11__20_, connection_3__11__19_, connection_3__11__18_, 
        connection_3__11__17_, connection_3__11__16_, connection_3__11__15_, 
        connection_3__11__14_, connection_3__11__13_, connection_3__11__12_, 
        connection_3__11__11_, connection_3__11__10_, connection_3__11__9_, 
        connection_3__11__8_, connection_3__11__7_, connection_3__11__6_, 
        connection_3__11__5_, connection_3__11__4_, connection_3__11__3_, 
        connection_3__11__2_, connection_3__11__1_, connection_3__11__0_, 
        connection_3__10__31_, connection_3__10__30_, connection_3__10__29_, 
        connection_3__10__28_, connection_3__10__27_, connection_3__10__26_, 
        connection_3__10__25_, connection_3__10__24_, connection_3__10__23_, 
        connection_3__10__22_, connection_3__10__21_, connection_3__10__20_, 
        connection_3__10__19_, connection_3__10__18_, connection_3__10__17_, 
        connection_3__10__16_, connection_3__10__15_, connection_3__10__14_, 
        connection_3__10__13_, connection_3__10__12_, connection_3__10__11_, 
        connection_3__10__10_, connection_3__10__9_, connection_3__10__8_, 
        connection_3__10__7_, connection_3__10__6_, connection_3__10__5_, 
        connection_3__10__4_, connection_3__10__3_, connection_3__10__2_, 
        connection_3__10__1_, connection_3__10__0_}), .i_en(n533), .i_cmd({
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__5__1_, 
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__5__0_}) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_2 middle_stage_6__middle_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__13_, 
        connection_valid_2__12_}), .i_data_bus({connection_2__13__31_, 
        connection_2__13__30_, connection_2__13__29_, connection_2__13__28_, 
        connection_2__13__27_, connection_2__13__26_, connection_2__13__25_, 
        connection_2__13__24_, connection_2__13__23_, connection_2__13__22_, 
        connection_2__13__21_, connection_2__13__20_, connection_2__13__19_, 
        connection_2__13__18_, connection_2__13__17_, connection_2__13__16_, 
        connection_2__13__15_, connection_2__13__14_, connection_2__13__13_, 
        connection_2__13__12_, connection_2__13__11_, connection_2__13__10_, 
        connection_2__13__9_, connection_2__13__8_, connection_2__13__7_, 
        connection_2__13__6_, connection_2__13__5_, connection_2__13__4_, 
        connection_2__13__3_, connection_2__13__2_, connection_2__13__1_, 
        connection_2__13__0_, connection_2__12__31_, connection_2__12__30_, 
        connection_2__12__29_, connection_2__12__28_, connection_2__12__27_, 
        connection_2__12__26_, connection_2__12__25_, connection_2__12__24_, 
        connection_2__12__23_, connection_2__12__22_, connection_2__12__21_, 
        connection_2__12__20_, connection_2__12__19_, connection_2__12__18_, 
        connection_2__12__17_, connection_2__12__16_, connection_2__12__15_, 
        connection_2__12__14_, connection_2__12__13_, connection_2__12__12_, 
        connection_2__12__11_, connection_2__12__10_, connection_2__12__9_, 
        connection_2__12__8_, connection_2__12__7_, connection_2__12__6_, 
        connection_2__12__5_, connection_2__12__4_, connection_2__12__3_, 
        connection_2__12__2_, connection_2__12__1_, connection_2__12__0_}), 
        .o_valid({connection_valid_3__13_, connection_valid_3__12_}), 
        .o_data_bus({connection_3__13__31_, connection_3__13__30_, 
        connection_3__13__29_, connection_3__13__28_, connection_3__13__27_, 
        connection_3__13__26_, connection_3__13__25_, connection_3__13__24_, 
        connection_3__13__23_, connection_3__13__22_, connection_3__13__21_, 
        connection_3__13__20_, connection_3__13__19_, connection_3__13__18_, 
        connection_3__13__17_, connection_3__13__16_, connection_3__13__15_, 
        connection_3__13__14_, connection_3__13__13_, connection_3__13__12_, 
        connection_3__13__11_, connection_3__13__10_, connection_3__13__9_, 
        connection_3__13__8_, connection_3__13__7_, connection_3__13__6_, 
        connection_3__13__5_, connection_3__13__4_, connection_3__13__3_, 
        connection_3__13__2_, connection_3__13__1_, connection_3__13__0_, 
        connection_3__12__31_, connection_3__12__30_, connection_3__12__29_, 
        connection_3__12__28_, connection_3__12__27_, connection_3__12__26_, 
        connection_3__12__25_, connection_3__12__24_, connection_3__12__23_, 
        connection_3__12__22_, connection_3__12__21_, connection_3__12__20_, 
        connection_3__12__19_, connection_3__12__18_, connection_3__12__17_, 
        connection_3__12__16_, connection_3__12__15_, connection_3__12__14_, 
        connection_3__12__13_, connection_3__12__12_, connection_3__12__11_, 
        connection_3__12__10_, connection_3__12__9_, connection_3__12__8_, 
        connection_3__12__7_, connection_3__12__6_, connection_3__12__5_, 
        connection_3__12__4_, connection_3__12__3_, connection_3__12__2_, 
        connection_3__12__1_, connection_3__12__0_}), .i_en(i_en), .i_cmd({
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__6__1_, 
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__6__0_}) );
  distribute_2x2_simple_seq_DATA_WIDTH32_COMMAND_WIDTH2_1 middle_stage_7__middle_stage ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_2__15_, 
        connection_valid_2__14_}), .i_data_bus({connection_2__15__31_, 
        connection_2__15__30_, connection_2__15__29_, connection_2__15__28_, 
        connection_2__15__27_, connection_2__15__26_, connection_2__15__25_, 
        connection_2__15__24_, connection_2__15__23_, connection_2__15__22_, 
        connection_2__15__21_, connection_2__15__20_, connection_2__15__19_, 
        connection_2__15__18_, connection_2__15__17_, connection_2__15__16_, 
        connection_2__15__15_, connection_2__15__14_, connection_2__15__13_, 
        connection_2__15__12_, connection_2__15__11_, connection_2__15__10_, 
        connection_2__15__9_, connection_2__15__8_, connection_2__15__7_, 
        connection_2__15__6_, connection_2__15__5_, connection_2__15__4_, 
        connection_2__15__3_, connection_2__15__2_, connection_2__15__1_, 
        connection_2__15__0_, connection_2__14__31_, connection_2__14__30_, 
        connection_2__14__29_, connection_2__14__28_, connection_2__14__27_, 
        connection_2__14__26_, connection_2__14__25_, connection_2__14__24_, 
        connection_2__14__23_, connection_2__14__22_, connection_2__14__21_, 
        connection_2__14__20_, connection_2__14__19_, connection_2__14__18_, 
        connection_2__14__17_, connection_2__14__16_, connection_2__14__15_, 
        connection_2__14__14_, connection_2__14__13_, connection_2__14__12_, 
        connection_2__14__11_, connection_2__14__10_, connection_2__14__9_, 
        connection_2__14__8_, connection_2__14__7_, connection_2__14__6_, 
        connection_2__14__5_, connection_2__14__4_, connection_2__14__3_, 
        connection_2__14__2_, connection_2__14__1_, connection_2__14__0_}), 
        .o_valid({connection_valid_3__15_, connection_valid_3__14_}), 
        .o_data_bus({connection_3__15__31_, connection_3__15__30_, 
        connection_3__15__29_, connection_3__15__28_, connection_3__15__27_, 
        connection_3__15__26_, connection_3__15__25_, connection_3__15__24_, 
        connection_3__15__23_, connection_3__15__22_, connection_3__15__21_, 
        connection_3__15__20_, connection_3__15__19_, connection_3__15__18_, 
        connection_3__15__17_, connection_3__15__16_, connection_3__15__15_, 
        connection_3__15__14_, connection_3__15__13_, connection_3__15__12_, 
        connection_3__15__11_, connection_3__15__10_, connection_3__15__9_, 
        connection_3__15__8_, connection_3__15__7_, connection_3__15__6_, 
        connection_3__15__5_, connection_3__15__4_, connection_3__15__3_, 
        connection_3__15__2_, connection_3__15__1_, connection_3__15__0_, 
        connection_3__14__31_, connection_3__14__30_, connection_3__14__29_, 
        connection_3__14__28_, connection_3__14__27_, connection_3__14__26_, 
        connection_3__14__25_, connection_3__14__24_, connection_3__14__23_, 
        connection_3__14__22_, connection_3__14__21_, connection_3__14__20_, 
        connection_3__14__19_, connection_3__14__18_, connection_3__14__17_, 
        connection_3__14__16_, connection_3__14__15_, connection_3__14__14_, 
        connection_3__14__13_, connection_3__14__12_, connection_3__14__11_, 
        connection_3__14__10_, connection_3__14__9_, connection_3__14__8_, 
        connection_3__14__7_, connection_3__14__6_, connection_3__14__5_, 
        connection_3__14__4_, connection_3__14__3_, connection_3__14__2_, 
        connection_3__14__1_, connection_3__14__0_}), .i_en(n533), .i_cmd({
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__7__1_, 
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__7__0_}) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_24 second_half_stages_4__sw_group_0__upper_group_0__upper_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_3__1_, 
        connection_valid_3__0_}), .i_data_bus({connection_3__1__31_, 
        connection_3__1__30_, connection_3__1__29_, connection_3__1__28_, 
        connection_3__1__27_, connection_3__1__26_, connection_3__1__25_, 
        connection_3__1__24_, connection_3__1__23_, connection_3__1__22_, 
        connection_3__1__21_, connection_3__1__20_, connection_3__1__19_, 
        connection_3__1__18_, connection_3__1__17_, connection_3__1__16_, 
        connection_3__1__15_, connection_3__1__14_, connection_3__1__13_, 
        connection_3__1__12_, connection_3__1__11_, connection_3__1__10_, 
        connection_3__1__9_, connection_3__1__8_, connection_3__1__7_, 
        connection_3__1__6_, connection_3__1__5_, connection_3__1__4_, 
        connection_3__1__3_, connection_3__1__2_, connection_3__1__1_, 
        connection_3__1__0_, connection_3__0__31_, connection_3__0__30_, 
        connection_3__0__29_, connection_3__0__28_, connection_3__0__27_, 
        connection_3__0__26_, connection_3__0__25_, connection_3__0__24_, 
        connection_3__0__23_, connection_3__0__22_, connection_3__0__21_, 
        connection_3__0__20_, connection_3__0__19_, connection_3__0__18_, 
        connection_3__0__17_, connection_3__0__16_, connection_3__0__15_, 
        connection_3__0__14_, connection_3__0__13_, connection_3__0__12_, 
        connection_3__0__11_, connection_3__0__10_, connection_3__0__9_, 
        connection_3__0__8_, connection_3__0__7_, connection_3__0__6_, 
        connection_3__0__5_, connection_3__0__4_, connection_3__0__3_, 
        connection_3__0__2_, connection_3__0__1_, connection_3__0__0_}), 
        .o_valid({connection_valid_4__1_, connection_valid_4__0_}), 
        .o_data_bus({connection_4__1__31_, connection_4__1__30_, 
        connection_4__1__29_, connection_4__1__28_, connection_4__1__27_, 
        connection_4__1__26_, connection_4__1__25_, connection_4__1__24_, 
        connection_4__1__23_, connection_4__1__22_, connection_4__1__21_, 
        connection_4__1__20_, connection_4__1__19_, connection_4__1__18_, 
        connection_4__1__17_, connection_4__1__16_, connection_4__1__15_, 
        connection_4__1__14_, connection_4__1__13_, connection_4__1__12_, 
        connection_4__1__11_, connection_4__1__10_, connection_4__1__9_, 
        connection_4__1__8_, connection_4__1__7_, connection_4__1__6_, 
        connection_4__1__5_, connection_4__1__4_, connection_4__1__3_, 
        connection_4__1__2_, connection_4__1__1_, connection_4__1__0_, 
        connection_4__0__31_, connection_4__0__30_, connection_4__0__29_, 
        connection_4__0__28_, connection_4__0__27_, connection_4__0__26_, 
        connection_4__0__25_, connection_4__0__24_, connection_4__0__23_, 
        connection_4__0__22_, connection_4__0__21_, connection_4__0__20_, 
        connection_4__0__19_, connection_4__0__18_, connection_4__0__17_, 
        connection_4__0__16_, connection_4__0__15_, connection_4__0__14_, 
        connection_4__0__13_, connection_4__0__12_, connection_4__0__11_, 
        connection_4__0__10_, connection_4__0__9_, connection_4__0__8_, 
        connection_4__0__7_, connection_4__0__6_, connection_4__0__5_, 
        connection_4__0__4_, connection_4__0__3_, connection_4__0__2_, 
        connection_4__0__1_, connection_4__0__0_}), .i_fwd_valid(
        fwd_connection_valid_sec_half[23]), .i_fwd_data_bus(
        fwd_connection_sec_half[767:736]), .o_fwd_valid(
        fwd_connection_valid_sec_half[22]), .o_fwd_data_bus(
        fwd_connection_sec_half[735:704]), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[119:115]) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_23 second_half_stages_4__sw_group_0__bottom_group_0__bottom_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_3__3_, 
        connection_valid_3__2_}), .i_data_bus({connection_3__3__31_, 
        connection_3__3__30_, connection_3__3__29_, connection_3__3__28_, 
        connection_3__3__27_, connection_3__3__26_, connection_3__3__25_, 
        connection_3__3__24_, connection_3__3__23_, connection_3__3__22_, 
        connection_3__3__21_, connection_3__3__20_, connection_3__3__19_, 
        connection_3__3__18_, connection_3__3__17_, connection_3__3__16_, 
        connection_3__3__15_, connection_3__3__14_, connection_3__3__13_, 
        connection_3__3__12_, connection_3__3__11_, connection_3__3__10_, 
        connection_3__3__9_, connection_3__3__8_, connection_3__3__7_, 
        connection_3__3__6_, connection_3__3__5_, connection_3__3__4_, 
        connection_3__3__3_, connection_3__3__2_, connection_3__3__1_, 
        connection_3__3__0_, connection_3__2__31_, connection_3__2__30_, 
        connection_3__2__29_, connection_3__2__28_, connection_3__2__27_, 
        connection_3__2__26_, connection_3__2__25_, connection_3__2__24_, 
        connection_3__2__23_, connection_3__2__22_, connection_3__2__21_, 
        connection_3__2__20_, connection_3__2__19_, connection_3__2__18_, 
        connection_3__2__17_, connection_3__2__16_, connection_3__2__15_, 
        connection_3__2__14_, connection_3__2__13_, connection_3__2__12_, 
        connection_3__2__11_, connection_3__2__10_, connection_3__2__9_, 
        connection_3__2__8_, connection_3__2__7_, connection_3__2__6_, 
        connection_3__2__5_, connection_3__2__4_, connection_3__2__3_, 
        connection_3__2__2_, connection_3__2__1_, connection_3__2__0_}), 
        .o_valid({connection_valid_4__3_, connection_valid_4__2_}), 
        .o_data_bus({connection_4__3__31_, connection_4__3__30_, 
        connection_4__3__29_, connection_4__3__28_, connection_4__3__27_, 
        connection_4__3__26_, connection_4__3__25_, connection_4__3__24_, 
        connection_4__3__23_, connection_4__3__22_, connection_4__3__21_, 
        connection_4__3__20_, connection_4__3__19_, connection_4__3__18_, 
        connection_4__3__17_, connection_4__3__16_, connection_4__3__15_, 
        connection_4__3__14_, connection_4__3__13_, connection_4__3__12_, 
        connection_4__3__11_, connection_4__3__10_, connection_4__3__9_, 
        connection_4__3__8_, connection_4__3__7_, connection_4__3__6_, 
        connection_4__3__5_, connection_4__3__4_, connection_4__3__3_, 
        connection_4__3__2_, connection_4__3__1_, connection_4__3__0_, 
        connection_4__2__31_, connection_4__2__30_, connection_4__2__29_, 
        connection_4__2__28_, connection_4__2__27_, connection_4__2__26_, 
        connection_4__2__25_, connection_4__2__24_, connection_4__2__23_, 
        connection_4__2__22_, connection_4__2__21_, connection_4__2__20_, 
        connection_4__2__19_, connection_4__2__18_, connection_4__2__17_, 
        connection_4__2__16_, connection_4__2__15_, connection_4__2__14_, 
        connection_4__2__13_, connection_4__2__12_, connection_4__2__11_, 
        connection_4__2__10_, connection_4__2__9_, connection_4__2__8_, 
        connection_4__2__7_, connection_4__2__6_, connection_4__2__5_, 
        connection_4__2__4_, connection_4__2__3_, connection_4__2__2_, 
        connection_4__2__1_, connection_4__2__0_}), .i_fwd_valid(
        fwd_connection_valid_sec_half[22]), .i_fwd_data_bus(
        fwd_connection_sec_half[735:704]), .o_fwd_valid(
        fwd_connection_valid_sec_half[23]), .o_fwd_data_bus(
        fwd_connection_sec_half[767:736]), .i_en(n533), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[114:110]) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_22 second_half_stages_4__sw_group_1__upper_group_0__upper_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_3__5_, 
        connection_valid_3__4_}), .i_data_bus({connection_3__5__31_, 
        connection_3__5__30_, connection_3__5__29_, connection_3__5__28_, 
        connection_3__5__27_, connection_3__5__26_, connection_3__5__25_, 
        connection_3__5__24_, connection_3__5__23_, connection_3__5__22_, 
        connection_3__5__21_, connection_3__5__20_, connection_3__5__19_, 
        connection_3__5__18_, connection_3__5__17_, connection_3__5__16_, 
        connection_3__5__15_, connection_3__5__14_, connection_3__5__13_, 
        connection_3__5__12_, connection_3__5__11_, connection_3__5__10_, 
        connection_3__5__9_, connection_3__5__8_, connection_3__5__7_, 
        connection_3__5__6_, connection_3__5__5_, connection_3__5__4_, 
        connection_3__5__3_, connection_3__5__2_, connection_3__5__1_, 
        connection_3__5__0_, connection_3__4__31_, connection_3__4__30_, 
        connection_3__4__29_, connection_3__4__28_, connection_3__4__27_, 
        connection_3__4__26_, connection_3__4__25_, connection_3__4__24_, 
        connection_3__4__23_, connection_3__4__22_, connection_3__4__21_, 
        connection_3__4__20_, connection_3__4__19_, connection_3__4__18_, 
        connection_3__4__17_, connection_3__4__16_, connection_3__4__15_, 
        connection_3__4__14_, connection_3__4__13_, connection_3__4__12_, 
        connection_3__4__11_, connection_3__4__10_, connection_3__4__9_, 
        connection_3__4__8_, connection_3__4__7_, connection_3__4__6_, 
        connection_3__4__5_, connection_3__4__4_, connection_3__4__3_, 
        connection_3__4__2_, connection_3__4__1_, connection_3__4__0_}), 
        .o_valid({connection_valid_4__5_, connection_valid_4__4_}), 
        .o_data_bus({connection_4__5__31_, connection_4__5__30_, 
        connection_4__5__29_, connection_4__5__28_, connection_4__5__27_, 
        connection_4__5__26_, connection_4__5__25_, connection_4__5__24_, 
        connection_4__5__23_, connection_4__5__22_, connection_4__5__21_, 
        connection_4__5__20_, connection_4__5__19_, connection_4__5__18_, 
        connection_4__5__17_, connection_4__5__16_, connection_4__5__15_, 
        connection_4__5__14_, connection_4__5__13_, connection_4__5__12_, 
        connection_4__5__11_, connection_4__5__10_, connection_4__5__9_, 
        connection_4__5__8_, connection_4__5__7_, connection_4__5__6_, 
        connection_4__5__5_, connection_4__5__4_, connection_4__5__3_, 
        connection_4__5__2_, connection_4__5__1_, connection_4__5__0_, 
        connection_4__4__31_, connection_4__4__30_, connection_4__4__29_, 
        connection_4__4__28_, connection_4__4__27_, connection_4__4__26_, 
        connection_4__4__25_, connection_4__4__24_, connection_4__4__23_, 
        connection_4__4__22_, connection_4__4__21_, connection_4__4__20_, 
        connection_4__4__19_, connection_4__4__18_, connection_4__4__17_, 
        connection_4__4__16_, connection_4__4__15_, connection_4__4__14_, 
        connection_4__4__13_, connection_4__4__12_, connection_4__4__11_, 
        connection_4__4__10_, connection_4__4__9_, connection_4__4__8_, 
        connection_4__4__7_, connection_4__4__6_, connection_4__4__5_, 
        connection_4__4__4_, connection_4__4__3_, connection_4__4__2_, 
        connection_4__4__1_, connection_4__4__0_}), .i_fwd_valid(
        fwd_connection_valid_sec_half[21]), .i_fwd_data_bus(
        fwd_connection_sec_half[703:672]), .o_fwd_valid(
        fwd_connection_valid_sec_half[20]), .o_fwd_data_bus(
        fwd_connection_sec_half[671:640]), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[109:105]) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_21 second_half_stages_4__sw_group_1__bottom_group_0__bottom_sw ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__7_, 
        connection_valid_3__6_}), .i_data_bus({connection_3__7__31_, 
        connection_3__7__30_, connection_3__7__29_, connection_3__7__28_, 
        connection_3__7__27_, connection_3__7__26_, connection_3__7__25_, 
        connection_3__7__24_, connection_3__7__23_, connection_3__7__22_, 
        connection_3__7__21_, connection_3__7__20_, connection_3__7__19_, 
        connection_3__7__18_, connection_3__7__17_, connection_3__7__16_, 
        connection_3__7__15_, connection_3__7__14_, connection_3__7__13_, 
        connection_3__7__12_, connection_3__7__11_, connection_3__7__10_, 
        connection_3__7__9_, connection_3__7__8_, connection_3__7__7_, 
        connection_3__7__6_, connection_3__7__5_, connection_3__7__4_, 
        connection_3__7__3_, connection_3__7__2_, connection_3__7__1_, 
        connection_3__7__0_, connection_3__6__31_, connection_3__6__30_, 
        connection_3__6__29_, connection_3__6__28_, connection_3__6__27_, 
        connection_3__6__26_, connection_3__6__25_, connection_3__6__24_, 
        connection_3__6__23_, connection_3__6__22_, connection_3__6__21_, 
        connection_3__6__20_, connection_3__6__19_, connection_3__6__18_, 
        connection_3__6__17_, connection_3__6__16_, connection_3__6__15_, 
        connection_3__6__14_, connection_3__6__13_, connection_3__6__12_, 
        connection_3__6__11_, connection_3__6__10_, connection_3__6__9_, 
        connection_3__6__8_, connection_3__6__7_, connection_3__6__6_, 
        connection_3__6__5_, connection_3__6__4_, connection_3__6__3_, 
        connection_3__6__2_, connection_3__6__1_, connection_3__6__0_}), 
        .o_valid({connection_valid_4__7_, connection_valid_4__6_}), 
        .o_data_bus({connection_4__7__31_, connection_4__7__30_, 
        connection_4__7__29_, connection_4__7__28_, connection_4__7__27_, 
        connection_4__7__26_, connection_4__7__25_, connection_4__7__24_, 
        connection_4__7__23_, connection_4__7__22_, connection_4__7__21_, 
        connection_4__7__20_, connection_4__7__19_, connection_4__7__18_, 
        connection_4__7__17_, connection_4__7__16_, connection_4__7__15_, 
        connection_4__7__14_, connection_4__7__13_, connection_4__7__12_, 
        connection_4__7__11_, connection_4__7__10_, connection_4__7__9_, 
        connection_4__7__8_, connection_4__7__7_, connection_4__7__6_, 
        connection_4__7__5_, connection_4__7__4_, connection_4__7__3_, 
        connection_4__7__2_, connection_4__7__1_, connection_4__7__0_, 
        connection_4__6__31_, connection_4__6__30_, connection_4__6__29_, 
        connection_4__6__28_, connection_4__6__27_, connection_4__6__26_, 
        connection_4__6__25_, connection_4__6__24_, connection_4__6__23_, 
        connection_4__6__22_, connection_4__6__21_, connection_4__6__20_, 
        connection_4__6__19_, connection_4__6__18_, connection_4__6__17_, 
        connection_4__6__16_, connection_4__6__15_, connection_4__6__14_, 
        connection_4__6__13_, connection_4__6__12_, connection_4__6__11_, 
        connection_4__6__10_, connection_4__6__9_, connection_4__6__8_, 
        connection_4__6__7_, connection_4__6__6_, connection_4__6__5_, 
        connection_4__6__4_, connection_4__6__3_, connection_4__6__2_, 
        connection_4__6__1_, connection_4__6__0_}), .i_fwd_valid(
        fwd_connection_valid_sec_half[20]), .i_fwd_data_bus(
        fwd_connection_sec_half[671:640]), .o_fwd_valid(
        fwd_connection_valid_sec_half[21]), .o_fwd_data_bus(
        fwd_connection_sec_half[703:672]), .i_en(n533), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[104:100]) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_20 second_half_stages_4__sw_group_2__upper_group_0__upper_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_3__9_, 
        connection_valid_3__8_}), .i_data_bus({connection_3__9__31_, 
        connection_3__9__30_, connection_3__9__29_, connection_3__9__28_, 
        connection_3__9__27_, connection_3__9__26_, connection_3__9__25_, 
        connection_3__9__24_, connection_3__9__23_, connection_3__9__22_, 
        connection_3__9__21_, connection_3__9__20_, connection_3__9__19_, 
        connection_3__9__18_, connection_3__9__17_, connection_3__9__16_, 
        connection_3__9__15_, connection_3__9__14_, connection_3__9__13_, 
        connection_3__9__12_, connection_3__9__11_, connection_3__9__10_, 
        connection_3__9__9_, connection_3__9__8_, connection_3__9__7_, 
        connection_3__9__6_, connection_3__9__5_, connection_3__9__4_, 
        connection_3__9__3_, connection_3__9__2_, connection_3__9__1_, 
        connection_3__9__0_, connection_3__8__31_, connection_3__8__30_, 
        connection_3__8__29_, connection_3__8__28_, connection_3__8__27_, 
        connection_3__8__26_, connection_3__8__25_, connection_3__8__24_, 
        connection_3__8__23_, connection_3__8__22_, connection_3__8__21_, 
        connection_3__8__20_, connection_3__8__19_, connection_3__8__18_, 
        connection_3__8__17_, connection_3__8__16_, connection_3__8__15_, 
        connection_3__8__14_, connection_3__8__13_, connection_3__8__12_, 
        connection_3__8__11_, connection_3__8__10_, connection_3__8__9_, 
        connection_3__8__8_, connection_3__8__7_, connection_3__8__6_, 
        connection_3__8__5_, connection_3__8__4_, connection_3__8__3_, 
        connection_3__8__2_, connection_3__8__1_, connection_3__8__0_}), 
        .o_valid({connection_valid_4__9_, connection_valid_4__8_}), 
        .o_data_bus({connection_4__9__31_, connection_4__9__30_, 
        connection_4__9__29_, connection_4__9__28_, connection_4__9__27_, 
        connection_4__9__26_, connection_4__9__25_, connection_4__9__24_, 
        connection_4__9__23_, connection_4__9__22_, connection_4__9__21_, 
        connection_4__9__20_, connection_4__9__19_, connection_4__9__18_, 
        connection_4__9__17_, connection_4__9__16_, connection_4__9__15_, 
        connection_4__9__14_, connection_4__9__13_, connection_4__9__12_, 
        connection_4__9__11_, connection_4__9__10_, connection_4__9__9_, 
        connection_4__9__8_, connection_4__9__7_, connection_4__9__6_, 
        connection_4__9__5_, connection_4__9__4_, connection_4__9__3_, 
        connection_4__9__2_, connection_4__9__1_, connection_4__9__0_, 
        connection_4__8__31_, connection_4__8__30_, connection_4__8__29_, 
        connection_4__8__28_, connection_4__8__27_, connection_4__8__26_, 
        connection_4__8__25_, connection_4__8__24_, connection_4__8__23_, 
        connection_4__8__22_, connection_4__8__21_, connection_4__8__20_, 
        connection_4__8__19_, connection_4__8__18_, connection_4__8__17_, 
        connection_4__8__16_, connection_4__8__15_, connection_4__8__14_, 
        connection_4__8__13_, connection_4__8__12_, connection_4__8__11_, 
        connection_4__8__10_, connection_4__8__9_, connection_4__8__8_, 
        connection_4__8__7_, connection_4__8__6_, connection_4__8__5_, 
        connection_4__8__4_, connection_4__8__3_, connection_4__8__2_, 
        connection_4__8__1_, connection_4__8__0_}), .i_fwd_valid(
        fwd_connection_valid_sec_half[19]), .i_fwd_data_bus(
        fwd_connection_sec_half[639:608]), .o_fwd_valid(
        fwd_connection_valid_sec_half[18]), .o_fwd_data_bus(
        fwd_connection_sec_half[607:576]), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[99:95]) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_19 second_half_stages_4__sw_group_2__bottom_group_0__bottom_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_3__11_, 
        connection_valid_3__10_}), .i_data_bus({connection_3__11__31_, 
        connection_3__11__30_, connection_3__11__29_, connection_3__11__28_, 
        connection_3__11__27_, connection_3__11__26_, connection_3__11__25_, 
        connection_3__11__24_, connection_3__11__23_, connection_3__11__22_, 
        connection_3__11__21_, connection_3__11__20_, connection_3__11__19_, 
        connection_3__11__18_, connection_3__11__17_, connection_3__11__16_, 
        connection_3__11__15_, connection_3__11__14_, connection_3__11__13_, 
        connection_3__11__12_, connection_3__11__11_, connection_3__11__10_, 
        connection_3__11__9_, connection_3__11__8_, connection_3__11__7_, 
        connection_3__11__6_, connection_3__11__5_, connection_3__11__4_, 
        connection_3__11__3_, connection_3__11__2_, connection_3__11__1_, 
        connection_3__11__0_, connection_3__10__31_, connection_3__10__30_, 
        connection_3__10__29_, connection_3__10__28_, connection_3__10__27_, 
        connection_3__10__26_, connection_3__10__25_, connection_3__10__24_, 
        connection_3__10__23_, connection_3__10__22_, connection_3__10__21_, 
        connection_3__10__20_, connection_3__10__19_, connection_3__10__18_, 
        connection_3__10__17_, connection_3__10__16_, connection_3__10__15_, 
        connection_3__10__14_, connection_3__10__13_, connection_3__10__12_, 
        connection_3__10__11_, connection_3__10__10_, connection_3__10__9_, 
        connection_3__10__8_, connection_3__10__7_, connection_3__10__6_, 
        connection_3__10__5_, connection_3__10__4_, connection_3__10__3_, 
        connection_3__10__2_, connection_3__10__1_, connection_3__10__0_}), 
        .o_valid({connection_valid_4__11_, connection_valid_4__10_}), 
        .o_data_bus({connection_4__11__31_, connection_4__11__30_, 
        connection_4__11__29_, connection_4__11__28_, connection_4__11__27_, 
        connection_4__11__26_, connection_4__11__25_, connection_4__11__24_, 
        connection_4__11__23_, connection_4__11__22_, connection_4__11__21_, 
        connection_4__11__20_, connection_4__11__19_, connection_4__11__18_, 
        connection_4__11__17_, connection_4__11__16_, connection_4__11__15_, 
        connection_4__11__14_, connection_4__11__13_, connection_4__11__12_, 
        connection_4__11__11_, connection_4__11__10_, connection_4__11__9_, 
        connection_4__11__8_, connection_4__11__7_, connection_4__11__6_, 
        connection_4__11__5_, connection_4__11__4_, connection_4__11__3_, 
        connection_4__11__2_, connection_4__11__1_, connection_4__11__0_, 
        connection_4__10__31_, connection_4__10__30_, connection_4__10__29_, 
        connection_4__10__28_, connection_4__10__27_, connection_4__10__26_, 
        connection_4__10__25_, connection_4__10__24_, connection_4__10__23_, 
        connection_4__10__22_, connection_4__10__21_, connection_4__10__20_, 
        connection_4__10__19_, connection_4__10__18_, connection_4__10__17_, 
        connection_4__10__16_, connection_4__10__15_, connection_4__10__14_, 
        connection_4__10__13_, connection_4__10__12_, connection_4__10__11_, 
        connection_4__10__10_, connection_4__10__9_, connection_4__10__8_, 
        connection_4__10__7_, connection_4__10__6_, connection_4__10__5_, 
        connection_4__10__4_, connection_4__10__3_, connection_4__10__2_, 
        connection_4__10__1_, connection_4__10__0_}), .i_fwd_valid(
        fwd_connection_valid_sec_half[18]), .i_fwd_data_bus(
        fwd_connection_sec_half[607:576]), .o_fwd_valid(
        fwd_connection_valid_sec_half[19]), .o_fwd_data_bus(
        fwd_connection_sec_half[639:608]), .i_en(n533), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[94:90]) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_18 second_half_stages_4__sw_group_3__upper_group_0__upper_sw ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_3__13_, 
        connection_valid_3__12_}), .i_data_bus({connection_3__13__31_, 
        connection_3__13__30_, connection_3__13__29_, connection_3__13__28_, 
        connection_3__13__27_, connection_3__13__26_, connection_3__13__25_, 
        connection_3__13__24_, connection_3__13__23_, connection_3__13__22_, 
        connection_3__13__21_, connection_3__13__20_, connection_3__13__19_, 
        connection_3__13__18_, connection_3__13__17_, connection_3__13__16_, 
        connection_3__13__15_, connection_3__13__14_, connection_3__13__13_, 
        connection_3__13__12_, connection_3__13__11_, connection_3__13__10_, 
        connection_3__13__9_, connection_3__13__8_, connection_3__13__7_, 
        connection_3__13__6_, connection_3__13__5_, connection_3__13__4_, 
        connection_3__13__3_, connection_3__13__2_, connection_3__13__1_, 
        connection_3__13__0_, connection_3__12__31_, connection_3__12__30_, 
        connection_3__12__29_, connection_3__12__28_, connection_3__12__27_, 
        connection_3__12__26_, connection_3__12__25_, connection_3__12__24_, 
        connection_3__12__23_, connection_3__12__22_, connection_3__12__21_, 
        connection_3__12__20_, connection_3__12__19_, connection_3__12__18_, 
        connection_3__12__17_, connection_3__12__16_, connection_3__12__15_, 
        connection_3__12__14_, connection_3__12__13_, connection_3__12__12_, 
        connection_3__12__11_, connection_3__12__10_, connection_3__12__9_, 
        connection_3__12__8_, connection_3__12__7_, connection_3__12__6_, 
        connection_3__12__5_, connection_3__12__4_, connection_3__12__3_, 
        connection_3__12__2_, connection_3__12__1_, connection_3__12__0_}), 
        .o_valid({connection_valid_4__13_, connection_valid_4__12_}), 
        .o_data_bus({connection_4__13__31_, connection_4__13__30_, 
        connection_4__13__29_, connection_4__13__28_, connection_4__13__27_, 
        connection_4__13__26_, connection_4__13__25_, connection_4__13__24_, 
        connection_4__13__23_, connection_4__13__22_, connection_4__13__21_, 
        connection_4__13__20_, connection_4__13__19_, connection_4__13__18_, 
        connection_4__13__17_, connection_4__13__16_, connection_4__13__15_, 
        connection_4__13__14_, connection_4__13__13_, connection_4__13__12_, 
        connection_4__13__11_, connection_4__13__10_, connection_4__13__9_, 
        connection_4__13__8_, connection_4__13__7_, connection_4__13__6_, 
        connection_4__13__5_, connection_4__13__4_, connection_4__13__3_, 
        connection_4__13__2_, connection_4__13__1_, connection_4__13__0_, 
        connection_4__12__31_, connection_4__12__30_, connection_4__12__29_, 
        connection_4__12__28_, connection_4__12__27_, connection_4__12__26_, 
        connection_4__12__25_, connection_4__12__24_, connection_4__12__23_, 
        connection_4__12__22_, connection_4__12__21_, connection_4__12__20_, 
        connection_4__12__19_, connection_4__12__18_, connection_4__12__17_, 
        connection_4__12__16_, connection_4__12__15_, connection_4__12__14_, 
        connection_4__12__13_, connection_4__12__12_, connection_4__12__11_, 
        connection_4__12__10_, connection_4__12__9_, connection_4__12__8_, 
        connection_4__12__7_, connection_4__12__6_, connection_4__12__5_, 
        connection_4__12__4_, connection_4__12__3_, connection_4__12__2_, 
        connection_4__12__1_, connection_4__12__0_}), .i_fwd_valid(
        fwd_connection_valid_sec_half[17]), .i_fwd_data_bus(
        fwd_connection_sec_half[575:544]), .o_fwd_valid(
        fwd_connection_valid_sec_half[16]), .o_fwd_data_bus(
        fwd_connection_sec_half[543:512]), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[89:85]) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_17 second_half_stages_4__sw_group_3__bottom_group_0__bottom_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_3__15_, 
        connection_valid_3__14_}), .i_data_bus({connection_3__15__31_, 
        connection_3__15__30_, connection_3__15__29_, connection_3__15__28_, 
        connection_3__15__27_, connection_3__15__26_, connection_3__15__25_, 
        connection_3__15__24_, connection_3__15__23_, connection_3__15__22_, 
        connection_3__15__21_, connection_3__15__20_, connection_3__15__19_, 
        connection_3__15__18_, connection_3__15__17_, connection_3__15__16_, 
        connection_3__15__15_, connection_3__15__14_, connection_3__15__13_, 
        connection_3__15__12_, connection_3__15__11_, connection_3__15__10_, 
        connection_3__15__9_, connection_3__15__8_, connection_3__15__7_, 
        connection_3__15__6_, connection_3__15__5_, connection_3__15__4_, 
        connection_3__15__3_, connection_3__15__2_, connection_3__15__1_, 
        connection_3__15__0_, connection_3__14__31_, connection_3__14__30_, 
        connection_3__14__29_, connection_3__14__28_, connection_3__14__27_, 
        connection_3__14__26_, connection_3__14__25_, connection_3__14__24_, 
        connection_3__14__23_, connection_3__14__22_, connection_3__14__21_, 
        connection_3__14__20_, connection_3__14__19_, connection_3__14__18_, 
        connection_3__14__17_, connection_3__14__16_, connection_3__14__15_, 
        connection_3__14__14_, connection_3__14__13_, connection_3__14__12_, 
        connection_3__14__11_, connection_3__14__10_, connection_3__14__9_, 
        connection_3__14__8_, connection_3__14__7_, connection_3__14__6_, 
        connection_3__14__5_, connection_3__14__4_, connection_3__14__3_, 
        connection_3__14__2_, connection_3__14__1_, connection_3__14__0_}), 
        .o_valid({connection_valid_4__15_, connection_valid_4__14_}), 
        .o_data_bus({connection_4__15__31_, connection_4__15__30_, 
        connection_4__15__29_, connection_4__15__28_, connection_4__15__27_, 
        connection_4__15__26_, connection_4__15__25_, connection_4__15__24_, 
        connection_4__15__23_, connection_4__15__22_, connection_4__15__21_, 
        connection_4__15__20_, connection_4__15__19_, connection_4__15__18_, 
        connection_4__15__17_, connection_4__15__16_, connection_4__15__15_, 
        connection_4__15__14_, connection_4__15__13_, connection_4__15__12_, 
        connection_4__15__11_, connection_4__15__10_, connection_4__15__9_, 
        connection_4__15__8_, connection_4__15__7_, connection_4__15__6_, 
        connection_4__15__5_, connection_4__15__4_, connection_4__15__3_, 
        connection_4__15__2_, connection_4__15__1_, connection_4__15__0_, 
        connection_4__14__31_, connection_4__14__30_, connection_4__14__29_, 
        connection_4__14__28_, connection_4__14__27_, connection_4__14__26_, 
        connection_4__14__25_, connection_4__14__24_, connection_4__14__23_, 
        connection_4__14__22_, connection_4__14__21_, connection_4__14__20_, 
        connection_4__14__19_, connection_4__14__18_, connection_4__14__17_, 
        connection_4__14__16_, connection_4__14__15_, connection_4__14__14_, 
        connection_4__14__13_, connection_4__14__12_, connection_4__14__11_, 
        connection_4__14__10_, connection_4__14__9_, connection_4__14__8_, 
        connection_4__14__7_, connection_4__14__6_, connection_4__14__5_, 
        connection_4__14__4_, connection_4__14__3_, connection_4__14__2_, 
        connection_4__14__1_, connection_4__14__0_}), .i_fwd_valid(
        fwd_connection_valid_sec_half[16]), .i_fwd_data_bus(
        fwd_connection_sec_half[543:512]), .o_fwd_valid(
        fwd_connection_valid_sec_half[17]), .o_fwd_data_bus(
        fwd_connection_sec_half[575:544]), .i_en(n533), .i_cmd(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[84:80]) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_16 second_half_stages_5__sw_group_0__upper_group_0__upper_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_4__1_, 
        connection_valid_4__0_}), .i_data_bus({connection_4__1__31_, 
        connection_4__1__30_, connection_4__1__29_, connection_4__1__28_, 
        connection_4__1__27_, connection_4__1__26_, connection_4__1__25_, 
        connection_4__1__24_, connection_4__1__23_, connection_4__1__22_, 
        connection_4__1__21_, connection_4__1__20_, connection_4__1__19_, 
        connection_4__1__18_, connection_4__1__17_, connection_4__1__16_, 
        connection_4__1__15_, connection_4__1__14_, connection_4__1__13_, 
        connection_4__1__12_, connection_4__1__11_, connection_4__1__10_, 
        connection_4__1__9_, connection_4__1__8_, connection_4__1__7_, 
        connection_4__1__6_, connection_4__1__5_, connection_4__1__4_, 
        connection_4__1__3_, connection_4__1__2_, connection_4__1__1_, 
        connection_4__1__0_, connection_4__0__31_, connection_4__0__30_, 
        connection_4__0__29_, connection_4__0__28_, connection_4__0__27_, 
        connection_4__0__26_, connection_4__0__25_, connection_4__0__24_, 
        connection_4__0__23_, connection_4__0__22_, connection_4__0__21_, 
        connection_4__0__20_, connection_4__0__19_, connection_4__0__18_, 
        connection_4__0__17_, connection_4__0__16_, connection_4__0__15_, 
        connection_4__0__14_, connection_4__0__13_, connection_4__0__12_, 
        connection_4__0__11_, connection_4__0__10_, connection_4__0__9_, 
        connection_4__0__8_, connection_4__0__7_, connection_4__0__6_, 
        connection_4__0__5_, connection_4__0__4_, connection_4__0__3_, 
        connection_4__0__2_, connection_4__0__1_, connection_4__0__0_}), 
        .o_valid({connection_valid_5__1_, connection_valid_5__0_}), 
        .o_data_bus({connection_5__1__31_, connection_5__1__30_, 
        connection_5__1__29_, connection_5__1__28_, connection_5__1__27_, 
        connection_5__1__26_, connection_5__1__25_, connection_5__1__24_, 
        connection_5__1__23_, connection_5__1__22_, connection_5__1__21_, 
        connection_5__1__20_, connection_5__1__19_, connection_5__1__18_, 
        connection_5__1__17_, connection_5__1__16_, connection_5__1__15_, 
        connection_5__1__14_, connection_5__1__13_, connection_5__1__12_, 
        connection_5__1__11_, connection_5__1__10_, connection_5__1__9_, 
        connection_5__1__8_, connection_5__1__7_, connection_5__1__6_, 
        connection_5__1__5_, connection_5__1__4_, connection_5__1__3_, 
        connection_5__1__2_, connection_5__1__1_, connection_5__1__0_, 
        connection_5__0__31_, connection_5__0__30_, connection_5__0__29_, 
        connection_5__0__28_, connection_5__0__27_, connection_5__0__26_, 
        connection_5__0__25_, connection_5__0__24_, connection_5__0__23_, 
        connection_5__0__22_, connection_5__0__21_, connection_5__0__20_, 
        connection_5__0__19_, connection_5__0__18_, connection_5__0__17_, 
        connection_5__0__16_, connection_5__0__15_, connection_5__0__14_, 
        connection_5__0__13_, connection_5__0__12_, connection_5__0__11_, 
        connection_5__0__10_, connection_5__0__9_, connection_5__0__8_, 
        connection_5__0__7_, connection_5__0__6_, connection_5__0__5_, 
        connection_5__0__4_, connection_5__0__3_, connection_5__0__2_, 
        connection_5__0__1_, connection_5__0__0_}), .i_fwd_valid(
        fwd_connection_valid_sec_half[15]), .i_fwd_data_bus(
        fwd_connection_sec_half[511:480]), .o_fwd_valid(
        fwd_connection_valid_sec_half[13]), .o_fwd_data_bus(
        fwd_connection_sec_half[447:416]), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[79:75]) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_15 second_half_stages_5__sw_group_0__upper_group_1__upper_sw ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__3_, 
        connection_valid_4__2_}), .i_data_bus({connection_4__3__31_, 
        connection_4__3__30_, connection_4__3__29_, connection_4__3__28_, 
        connection_4__3__27_, connection_4__3__26_, connection_4__3__25_, 
        connection_4__3__24_, connection_4__3__23_, connection_4__3__22_, 
        connection_4__3__21_, connection_4__3__20_, connection_4__3__19_, 
        connection_4__3__18_, connection_4__3__17_, connection_4__3__16_, 
        connection_4__3__15_, connection_4__3__14_, connection_4__3__13_, 
        connection_4__3__12_, connection_4__3__11_, connection_4__3__10_, 
        connection_4__3__9_, connection_4__3__8_, connection_4__3__7_, 
        connection_4__3__6_, connection_4__3__5_, connection_4__3__4_, 
        connection_4__3__3_, connection_4__3__2_, connection_4__3__1_, 
        connection_4__3__0_, connection_4__2__31_, connection_4__2__30_, 
        connection_4__2__29_, connection_4__2__28_, connection_4__2__27_, 
        connection_4__2__26_, connection_4__2__25_, connection_4__2__24_, 
        connection_4__2__23_, connection_4__2__22_, connection_4__2__21_, 
        connection_4__2__20_, connection_4__2__19_, connection_4__2__18_, 
        connection_4__2__17_, connection_4__2__16_, connection_4__2__15_, 
        connection_4__2__14_, connection_4__2__13_, connection_4__2__12_, 
        connection_4__2__11_, connection_4__2__10_, connection_4__2__9_, 
        connection_4__2__8_, connection_4__2__7_, connection_4__2__6_, 
        connection_4__2__5_, connection_4__2__4_, connection_4__2__3_, 
        connection_4__2__2_, connection_4__2__1_, connection_4__2__0_}), 
        .o_valid({connection_valid_5__3_, connection_valid_5__2_}), 
        .o_data_bus({connection_5__3__31_, connection_5__3__30_, 
        connection_5__3__29_, connection_5__3__28_, connection_5__3__27_, 
        connection_5__3__26_, connection_5__3__25_, connection_5__3__24_, 
        connection_5__3__23_, connection_5__3__22_, connection_5__3__21_, 
        connection_5__3__20_, connection_5__3__19_, connection_5__3__18_, 
        connection_5__3__17_, connection_5__3__16_, connection_5__3__15_, 
        connection_5__3__14_, connection_5__3__13_, connection_5__3__12_, 
        connection_5__3__11_, connection_5__3__10_, connection_5__3__9_, 
        connection_5__3__8_, connection_5__3__7_, connection_5__3__6_, 
        connection_5__3__5_, connection_5__3__4_, connection_5__3__3_, 
        connection_5__3__2_, connection_5__3__1_, connection_5__3__0_, 
        connection_5__2__31_, connection_5__2__30_, connection_5__2__29_, 
        connection_5__2__28_, connection_5__2__27_, connection_5__2__26_, 
        connection_5__2__25_, connection_5__2__24_, connection_5__2__23_, 
        connection_5__2__22_, connection_5__2__21_, connection_5__2__20_, 
        connection_5__2__19_, connection_5__2__18_, connection_5__2__17_, 
        connection_5__2__16_, connection_5__2__15_, connection_5__2__14_, 
        connection_5__2__13_, connection_5__2__12_, connection_5__2__11_, 
        connection_5__2__10_, connection_5__2__9_, connection_5__2__8_, 
        connection_5__2__7_, connection_5__2__6_, connection_5__2__5_, 
        connection_5__2__4_, connection_5__2__3_, connection_5__2__2_, 
        connection_5__2__1_, connection_5__2__0_}), .i_fwd_valid(
        fwd_connection_valid_sec_half[14]), .i_fwd_data_bus(
        fwd_connection_sec_half[479:448]), .o_fwd_valid(
        fwd_connection_valid_sec_half[12]), .o_fwd_data_bus(
        fwd_connection_sec_half[415:384]), .i_en(n533), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[74:70]) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_14 second_half_stages_5__sw_group_0__bottom_group_0__bottom_sw ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__5_, 
        connection_valid_4__4_}), .i_data_bus({connection_4__5__31_, 
        connection_4__5__30_, connection_4__5__29_, connection_4__5__28_, 
        connection_4__5__27_, connection_4__5__26_, connection_4__5__25_, 
        connection_4__5__24_, connection_4__5__23_, connection_4__5__22_, 
        connection_4__5__21_, connection_4__5__20_, connection_4__5__19_, 
        connection_4__5__18_, connection_4__5__17_, connection_4__5__16_, 
        connection_4__5__15_, connection_4__5__14_, connection_4__5__13_, 
        connection_4__5__12_, connection_4__5__11_, connection_4__5__10_, 
        connection_4__5__9_, connection_4__5__8_, connection_4__5__7_, 
        connection_4__5__6_, connection_4__5__5_, connection_4__5__4_, 
        connection_4__5__3_, connection_4__5__2_, connection_4__5__1_, 
        connection_4__5__0_, connection_4__4__31_, connection_4__4__30_, 
        connection_4__4__29_, connection_4__4__28_, connection_4__4__27_, 
        connection_4__4__26_, connection_4__4__25_, connection_4__4__24_, 
        connection_4__4__23_, connection_4__4__22_, connection_4__4__21_, 
        connection_4__4__20_, connection_4__4__19_, connection_4__4__18_, 
        connection_4__4__17_, connection_4__4__16_, connection_4__4__15_, 
        connection_4__4__14_, connection_4__4__13_, connection_4__4__12_, 
        connection_4__4__11_, connection_4__4__10_, connection_4__4__9_, 
        connection_4__4__8_, connection_4__4__7_, connection_4__4__6_, 
        connection_4__4__5_, connection_4__4__4_, connection_4__4__3_, 
        connection_4__4__2_, connection_4__4__1_, connection_4__4__0_}), 
        .o_valid({connection_valid_5__5_, connection_valid_5__4_}), 
        .o_data_bus({connection_5__5__31_, connection_5__5__30_, 
        connection_5__5__29_, connection_5__5__28_, connection_5__5__27_, 
        connection_5__5__26_, connection_5__5__25_, connection_5__5__24_, 
        connection_5__5__23_, connection_5__5__22_, connection_5__5__21_, 
        connection_5__5__20_, connection_5__5__19_, connection_5__5__18_, 
        connection_5__5__17_, connection_5__5__16_, connection_5__5__15_, 
        connection_5__5__14_, connection_5__5__13_, connection_5__5__12_, 
        connection_5__5__11_, connection_5__5__10_, connection_5__5__9_, 
        connection_5__5__8_, connection_5__5__7_, connection_5__5__6_, 
        connection_5__5__5_, connection_5__5__4_, connection_5__5__3_, 
        connection_5__5__2_, connection_5__5__1_, connection_5__5__0_, 
        connection_5__4__31_, connection_5__4__30_, connection_5__4__29_, 
        connection_5__4__28_, connection_5__4__27_, connection_5__4__26_, 
        connection_5__4__25_, connection_5__4__24_, connection_5__4__23_, 
        connection_5__4__22_, connection_5__4__21_, connection_5__4__20_, 
        connection_5__4__19_, connection_5__4__18_, connection_5__4__17_, 
        connection_5__4__16_, connection_5__4__15_, connection_5__4__14_, 
        connection_5__4__13_, connection_5__4__12_, connection_5__4__11_, 
        connection_5__4__10_, connection_5__4__9_, connection_5__4__8_, 
        connection_5__4__7_, connection_5__4__6_, connection_5__4__5_, 
        connection_5__4__4_, connection_5__4__3_, connection_5__4__2_, 
        connection_5__4__1_, connection_5__4__0_}), .i_fwd_valid(
        fwd_connection_valid_sec_half[13]), .i_fwd_data_bus(
        fwd_connection_sec_half[447:416]), .o_fwd_valid(
        fwd_connection_valid_sec_half[15]), .o_fwd_data_bus(
        fwd_connection_sec_half[511:480]), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[69:65]) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_13 second_half_stages_5__sw_group_0__bottom_group_1__bottom_sw ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__7_, 
        connection_valid_4__6_}), .i_data_bus({connection_4__7__31_, 
        connection_4__7__30_, connection_4__7__29_, connection_4__7__28_, 
        connection_4__7__27_, connection_4__7__26_, connection_4__7__25_, 
        connection_4__7__24_, connection_4__7__23_, connection_4__7__22_, 
        connection_4__7__21_, connection_4__7__20_, connection_4__7__19_, 
        connection_4__7__18_, connection_4__7__17_, connection_4__7__16_, 
        connection_4__7__15_, connection_4__7__14_, connection_4__7__13_, 
        connection_4__7__12_, connection_4__7__11_, connection_4__7__10_, 
        connection_4__7__9_, connection_4__7__8_, connection_4__7__7_, 
        connection_4__7__6_, connection_4__7__5_, connection_4__7__4_, 
        connection_4__7__3_, connection_4__7__2_, connection_4__7__1_, 
        connection_4__7__0_, connection_4__6__31_, connection_4__6__30_, 
        connection_4__6__29_, connection_4__6__28_, connection_4__6__27_, 
        connection_4__6__26_, connection_4__6__25_, connection_4__6__24_, 
        connection_4__6__23_, connection_4__6__22_, connection_4__6__21_, 
        connection_4__6__20_, connection_4__6__19_, connection_4__6__18_, 
        connection_4__6__17_, connection_4__6__16_, connection_4__6__15_, 
        connection_4__6__14_, connection_4__6__13_, connection_4__6__12_, 
        connection_4__6__11_, connection_4__6__10_, connection_4__6__9_, 
        connection_4__6__8_, connection_4__6__7_, connection_4__6__6_, 
        connection_4__6__5_, connection_4__6__4_, connection_4__6__3_, 
        connection_4__6__2_, connection_4__6__1_, connection_4__6__0_}), 
        .o_valid({connection_valid_5__7_, connection_valid_5__6_}), 
        .o_data_bus({connection_5__7__31_, connection_5__7__30_, 
        connection_5__7__29_, connection_5__7__28_, connection_5__7__27_, 
        connection_5__7__26_, connection_5__7__25_, connection_5__7__24_, 
        connection_5__7__23_, connection_5__7__22_, connection_5__7__21_, 
        connection_5__7__20_, connection_5__7__19_, connection_5__7__18_, 
        connection_5__7__17_, connection_5__7__16_, connection_5__7__15_, 
        connection_5__7__14_, connection_5__7__13_, connection_5__7__12_, 
        connection_5__7__11_, connection_5__7__10_, connection_5__7__9_, 
        connection_5__7__8_, connection_5__7__7_, connection_5__7__6_, 
        connection_5__7__5_, connection_5__7__4_, connection_5__7__3_, 
        connection_5__7__2_, connection_5__7__1_, connection_5__7__0_, 
        connection_5__6__31_, connection_5__6__30_, connection_5__6__29_, 
        connection_5__6__28_, connection_5__6__27_, connection_5__6__26_, 
        connection_5__6__25_, connection_5__6__24_, connection_5__6__23_, 
        connection_5__6__22_, connection_5__6__21_, connection_5__6__20_, 
        connection_5__6__19_, connection_5__6__18_, connection_5__6__17_, 
        connection_5__6__16_, connection_5__6__15_, connection_5__6__14_, 
        connection_5__6__13_, connection_5__6__12_, connection_5__6__11_, 
        connection_5__6__10_, connection_5__6__9_, connection_5__6__8_, 
        connection_5__6__7_, connection_5__6__6_, connection_5__6__5_, 
        connection_5__6__4_, connection_5__6__3_, connection_5__6__2_, 
        connection_5__6__1_, connection_5__6__0_}), .i_fwd_valid(
        fwd_connection_valid_sec_half[12]), .i_fwd_data_bus(
        fwd_connection_sec_half[415:384]), .o_fwd_valid(
        fwd_connection_valid_sec_half[14]), .o_fwd_data_bus(
        fwd_connection_sec_half[479:448]), .i_en(n533), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[64:60]) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_12 second_half_stages_5__sw_group_1__upper_group_0__upper_sw ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__9_, 
        connection_valid_4__8_}), .i_data_bus({connection_4__9__31_, 
        connection_4__9__30_, connection_4__9__29_, connection_4__9__28_, 
        connection_4__9__27_, connection_4__9__26_, connection_4__9__25_, 
        connection_4__9__24_, connection_4__9__23_, connection_4__9__22_, 
        connection_4__9__21_, connection_4__9__20_, connection_4__9__19_, 
        connection_4__9__18_, connection_4__9__17_, connection_4__9__16_, 
        connection_4__9__15_, connection_4__9__14_, connection_4__9__13_, 
        connection_4__9__12_, connection_4__9__11_, connection_4__9__10_, 
        connection_4__9__9_, connection_4__9__8_, connection_4__9__7_, 
        connection_4__9__6_, connection_4__9__5_, connection_4__9__4_, 
        connection_4__9__3_, connection_4__9__2_, connection_4__9__1_, 
        connection_4__9__0_, connection_4__8__31_, connection_4__8__30_, 
        connection_4__8__29_, connection_4__8__28_, connection_4__8__27_, 
        connection_4__8__26_, connection_4__8__25_, connection_4__8__24_, 
        connection_4__8__23_, connection_4__8__22_, connection_4__8__21_, 
        connection_4__8__20_, connection_4__8__19_, connection_4__8__18_, 
        connection_4__8__17_, connection_4__8__16_, connection_4__8__15_, 
        connection_4__8__14_, connection_4__8__13_, connection_4__8__12_, 
        connection_4__8__11_, connection_4__8__10_, connection_4__8__9_, 
        connection_4__8__8_, connection_4__8__7_, connection_4__8__6_, 
        connection_4__8__5_, connection_4__8__4_, connection_4__8__3_, 
        connection_4__8__2_, connection_4__8__1_, connection_4__8__0_}), 
        .o_valid({connection_valid_5__9_, connection_valid_5__8_}), 
        .o_data_bus({connection_5__9__31_, connection_5__9__30_, 
        connection_5__9__29_, connection_5__9__28_, connection_5__9__27_, 
        connection_5__9__26_, connection_5__9__25_, connection_5__9__24_, 
        connection_5__9__23_, connection_5__9__22_, connection_5__9__21_, 
        connection_5__9__20_, connection_5__9__19_, connection_5__9__18_, 
        connection_5__9__17_, connection_5__9__16_, connection_5__9__15_, 
        connection_5__9__14_, connection_5__9__13_, connection_5__9__12_, 
        connection_5__9__11_, connection_5__9__10_, connection_5__9__9_, 
        connection_5__9__8_, connection_5__9__7_, connection_5__9__6_, 
        connection_5__9__5_, connection_5__9__4_, connection_5__9__3_, 
        connection_5__9__2_, connection_5__9__1_, connection_5__9__0_, 
        connection_5__8__31_, connection_5__8__30_, connection_5__8__29_, 
        connection_5__8__28_, connection_5__8__27_, connection_5__8__26_, 
        connection_5__8__25_, connection_5__8__24_, connection_5__8__23_, 
        connection_5__8__22_, connection_5__8__21_, connection_5__8__20_, 
        connection_5__8__19_, connection_5__8__18_, connection_5__8__17_, 
        connection_5__8__16_, connection_5__8__15_, connection_5__8__14_, 
        connection_5__8__13_, connection_5__8__12_, connection_5__8__11_, 
        connection_5__8__10_, connection_5__8__9_, connection_5__8__8_, 
        connection_5__8__7_, connection_5__8__6_, connection_5__8__5_, 
        connection_5__8__4_, connection_5__8__3_, connection_5__8__2_, 
        connection_5__8__1_, connection_5__8__0_}), .i_fwd_valid(
        fwd_connection_valid_sec_half[11]), .i_fwd_data_bus(
        fwd_connection_sec_half[383:352]), .o_fwd_valid(
        fwd_connection_valid_sec_half[9]), .o_fwd_data_bus(
        fwd_connection_sec_half[319:288]), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[59:55]) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_11 second_half_stages_5__sw_group_1__upper_group_1__upper_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_4__11_, 
        connection_valid_4__10_}), .i_data_bus({connection_4__11__31_, 
        connection_4__11__30_, connection_4__11__29_, connection_4__11__28_, 
        connection_4__11__27_, connection_4__11__26_, connection_4__11__25_, 
        connection_4__11__24_, connection_4__11__23_, connection_4__11__22_, 
        connection_4__11__21_, connection_4__11__20_, connection_4__11__19_, 
        connection_4__11__18_, connection_4__11__17_, connection_4__11__16_, 
        connection_4__11__15_, connection_4__11__14_, connection_4__11__13_, 
        connection_4__11__12_, connection_4__11__11_, connection_4__11__10_, 
        connection_4__11__9_, connection_4__11__8_, connection_4__11__7_, 
        connection_4__11__6_, connection_4__11__5_, connection_4__11__4_, 
        connection_4__11__3_, connection_4__11__2_, connection_4__11__1_, 
        connection_4__11__0_, connection_4__10__31_, connection_4__10__30_, 
        connection_4__10__29_, connection_4__10__28_, connection_4__10__27_, 
        connection_4__10__26_, connection_4__10__25_, connection_4__10__24_, 
        connection_4__10__23_, connection_4__10__22_, connection_4__10__21_, 
        connection_4__10__20_, connection_4__10__19_, connection_4__10__18_, 
        connection_4__10__17_, connection_4__10__16_, connection_4__10__15_, 
        connection_4__10__14_, connection_4__10__13_, connection_4__10__12_, 
        connection_4__10__11_, connection_4__10__10_, connection_4__10__9_, 
        connection_4__10__8_, connection_4__10__7_, connection_4__10__6_, 
        connection_4__10__5_, connection_4__10__4_, connection_4__10__3_, 
        connection_4__10__2_, connection_4__10__1_, connection_4__10__0_}), 
        .o_valid({connection_valid_5__11_, connection_valid_5__10_}), 
        .o_data_bus({connection_5__11__31_, connection_5__11__30_, 
        connection_5__11__29_, connection_5__11__28_, connection_5__11__27_, 
        connection_5__11__26_, connection_5__11__25_, connection_5__11__24_, 
        connection_5__11__23_, connection_5__11__22_, connection_5__11__21_, 
        connection_5__11__20_, connection_5__11__19_, connection_5__11__18_, 
        connection_5__11__17_, connection_5__11__16_, connection_5__11__15_, 
        connection_5__11__14_, connection_5__11__13_, connection_5__11__12_, 
        connection_5__11__11_, connection_5__11__10_, connection_5__11__9_, 
        connection_5__11__8_, connection_5__11__7_, connection_5__11__6_, 
        connection_5__11__5_, connection_5__11__4_, connection_5__11__3_, 
        connection_5__11__2_, connection_5__11__1_, connection_5__11__0_, 
        connection_5__10__31_, connection_5__10__30_, connection_5__10__29_, 
        connection_5__10__28_, connection_5__10__27_, connection_5__10__26_, 
        connection_5__10__25_, connection_5__10__24_, connection_5__10__23_, 
        connection_5__10__22_, connection_5__10__21_, connection_5__10__20_, 
        connection_5__10__19_, connection_5__10__18_, connection_5__10__17_, 
        connection_5__10__16_, connection_5__10__15_, connection_5__10__14_, 
        connection_5__10__13_, connection_5__10__12_, connection_5__10__11_, 
        connection_5__10__10_, connection_5__10__9_, connection_5__10__8_, 
        connection_5__10__7_, connection_5__10__6_, connection_5__10__5_, 
        connection_5__10__4_, connection_5__10__3_, connection_5__10__2_, 
        connection_5__10__1_, connection_5__10__0_}), .i_fwd_valid(
        fwd_connection_valid_sec_half[10]), .i_fwd_data_bus(
        fwd_connection_sec_half[351:320]), .o_fwd_valid(
        fwd_connection_valid_sec_half[8]), .o_fwd_data_bus(
        fwd_connection_sec_half[287:256]), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[54:50]) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_10 second_half_stages_5__sw_group_1__bottom_group_0__bottom_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_4__13_, 
        connection_valid_4__12_}), .i_data_bus({connection_4__13__31_, 
        connection_4__13__30_, connection_4__13__29_, connection_4__13__28_, 
        connection_4__13__27_, connection_4__13__26_, connection_4__13__25_, 
        connection_4__13__24_, connection_4__13__23_, connection_4__13__22_, 
        connection_4__13__21_, connection_4__13__20_, connection_4__13__19_, 
        connection_4__13__18_, connection_4__13__17_, connection_4__13__16_, 
        connection_4__13__15_, connection_4__13__14_, connection_4__13__13_, 
        connection_4__13__12_, connection_4__13__11_, connection_4__13__10_, 
        connection_4__13__9_, connection_4__13__8_, connection_4__13__7_, 
        connection_4__13__6_, connection_4__13__5_, connection_4__13__4_, 
        connection_4__13__3_, connection_4__13__2_, connection_4__13__1_, 
        connection_4__13__0_, connection_4__12__31_, connection_4__12__30_, 
        connection_4__12__29_, connection_4__12__28_, connection_4__12__27_, 
        connection_4__12__26_, connection_4__12__25_, connection_4__12__24_, 
        connection_4__12__23_, connection_4__12__22_, connection_4__12__21_, 
        connection_4__12__20_, connection_4__12__19_, connection_4__12__18_, 
        connection_4__12__17_, connection_4__12__16_, connection_4__12__15_, 
        connection_4__12__14_, connection_4__12__13_, connection_4__12__12_, 
        connection_4__12__11_, connection_4__12__10_, connection_4__12__9_, 
        connection_4__12__8_, connection_4__12__7_, connection_4__12__6_, 
        connection_4__12__5_, connection_4__12__4_, connection_4__12__3_, 
        connection_4__12__2_, connection_4__12__1_, connection_4__12__0_}), 
        .o_valid({connection_valid_5__13_, connection_valid_5__12_}), 
        .o_data_bus({connection_5__13__31_, connection_5__13__30_, 
        connection_5__13__29_, connection_5__13__28_, connection_5__13__27_, 
        connection_5__13__26_, connection_5__13__25_, connection_5__13__24_, 
        connection_5__13__23_, connection_5__13__22_, connection_5__13__21_, 
        connection_5__13__20_, connection_5__13__19_, connection_5__13__18_, 
        connection_5__13__17_, connection_5__13__16_, connection_5__13__15_, 
        connection_5__13__14_, connection_5__13__13_, connection_5__13__12_, 
        connection_5__13__11_, connection_5__13__10_, connection_5__13__9_, 
        connection_5__13__8_, connection_5__13__7_, connection_5__13__6_, 
        connection_5__13__5_, connection_5__13__4_, connection_5__13__3_, 
        connection_5__13__2_, connection_5__13__1_, connection_5__13__0_, 
        connection_5__12__31_, connection_5__12__30_, connection_5__12__29_, 
        connection_5__12__28_, connection_5__12__27_, connection_5__12__26_, 
        connection_5__12__25_, connection_5__12__24_, connection_5__12__23_, 
        connection_5__12__22_, connection_5__12__21_, connection_5__12__20_, 
        connection_5__12__19_, connection_5__12__18_, connection_5__12__17_, 
        connection_5__12__16_, connection_5__12__15_, connection_5__12__14_, 
        connection_5__12__13_, connection_5__12__12_, connection_5__12__11_, 
        connection_5__12__10_, connection_5__12__9_, connection_5__12__8_, 
        connection_5__12__7_, connection_5__12__6_, connection_5__12__5_, 
        connection_5__12__4_, connection_5__12__3_, connection_5__12__2_, 
        connection_5__12__1_, connection_5__12__0_}), .i_fwd_valid(
        fwd_connection_valid_sec_half[9]), .i_fwd_data_bus(
        fwd_connection_sec_half[319:288]), .o_fwd_valid(
        fwd_connection_valid_sec_half[11]), .o_fwd_data_bus(
        fwd_connection_sec_half[383:352]), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[49:45]) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_9 second_half_stages_5__sw_group_1__bottom_group_1__bottom_sw ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_4__15_, 
        connection_valid_4__14_}), .i_data_bus({connection_4__15__31_, 
        connection_4__15__30_, connection_4__15__29_, connection_4__15__28_, 
        connection_4__15__27_, connection_4__15__26_, connection_4__15__25_, 
        connection_4__15__24_, connection_4__15__23_, connection_4__15__22_, 
        connection_4__15__21_, connection_4__15__20_, connection_4__15__19_, 
        connection_4__15__18_, connection_4__15__17_, connection_4__15__16_, 
        connection_4__15__15_, connection_4__15__14_, connection_4__15__13_, 
        connection_4__15__12_, connection_4__15__11_, connection_4__15__10_, 
        connection_4__15__9_, connection_4__15__8_, connection_4__15__7_, 
        connection_4__15__6_, connection_4__15__5_, connection_4__15__4_, 
        connection_4__15__3_, connection_4__15__2_, connection_4__15__1_, 
        connection_4__15__0_, connection_4__14__31_, connection_4__14__30_, 
        connection_4__14__29_, connection_4__14__28_, connection_4__14__27_, 
        connection_4__14__26_, connection_4__14__25_, connection_4__14__24_, 
        connection_4__14__23_, connection_4__14__22_, connection_4__14__21_, 
        connection_4__14__20_, connection_4__14__19_, connection_4__14__18_, 
        connection_4__14__17_, connection_4__14__16_, connection_4__14__15_, 
        connection_4__14__14_, connection_4__14__13_, connection_4__14__12_, 
        connection_4__14__11_, connection_4__14__10_, connection_4__14__9_, 
        connection_4__14__8_, connection_4__14__7_, connection_4__14__6_, 
        connection_4__14__5_, connection_4__14__4_, connection_4__14__3_, 
        connection_4__14__2_, connection_4__14__1_, connection_4__14__0_}), 
        .o_valid({connection_valid_5__15_, connection_valid_5__14_}), 
        .o_data_bus({connection_5__15__31_, connection_5__15__30_, 
        connection_5__15__29_, connection_5__15__28_, connection_5__15__27_, 
        connection_5__15__26_, connection_5__15__25_, connection_5__15__24_, 
        connection_5__15__23_, connection_5__15__22_, connection_5__15__21_, 
        connection_5__15__20_, connection_5__15__19_, connection_5__15__18_, 
        connection_5__15__17_, connection_5__15__16_, connection_5__15__15_, 
        connection_5__15__14_, connection_5__15__13_, connection_5__15__12_, 
        connection_5__15__11_, connection_5__15__10_, connection_5__15__9_, 
        connection_5__15__8_, connection_5__15__7_, connection_5__15__6_, 
        connection_5__15__5_, connection_5__15__4_, connection_5__15__3_, 
        connection_5__15__2_, connection_5__15__1_, connection_5__15__0_, 
        connection_5__14__31_, connection_5__14__30_, connection_5__14__29_, 
        connection_5__14__28_, connection_5__14__27_, connection_5__14__26_, 
        connection_5__14__25_, connection_5__14__24_, connection_5__14__23_, 
        connection_5__14__22_, connection_5__14__21_, connection_5__14__20_, 
        connection_5__14__19_, connection_5__14__18_, connection_5__14__17_, 
        connection_5__14__16_, connection_5__14__15_, connection_5__14__14_, 
        connection_5__14__13_, connection_5__14__12_, connection_5__14__11_, 
        connection_5__14__10_, connection_5__14__9_, connection_5__14__8_, 
        connection_5__14__7_, connection_5__14__6_, connection_5__14__5_, 
        connection_5__14__4_, connection_5__14__3_, connection_5__14__2_, 
        connection_5__14__1_, connection_5__14__0_}), .i_fwd_valid(
        fwd_connection_valid_sec_half[8]), .i_fwd_data_bus(
        fwd_connection_sec_half[287:256]), .o_fwd_valid(
        fwd_connection_valid_sec_half[10]), .o_fwd_data_bus(
        fwd_connection_sec_half[351:320]), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[44:40]) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_8 second_half_stages_6__sw_group_0__upper_group_0__upper_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_5__1_, 
        connection_valid_5__0_}), .i_data_bus({connection_5__1__31_, 
        connection_5__1__30_, connection_5__1__29_, connection_5__1__28_, 
        connection_5__1__27_, connection_5__1__26_, connection_5__1__25_, 
        connection_5__1__24_, connection_5__1__23_, connection_5__1__22_, 
        connection_5__1__21_, connection_5__1__20_, connection_5__1__19_, 
        connection_5__1__18_, connection_5__1__17_, connection_5__1__16_, 
        connection_5__1__15_, connection_5__1__14_, connection_5__1__13_, 
        connection_5__1__12_, connection_5__1__11_, connection_5__1__10_, 
        connection_5__1__9_, connection_5__1__8_, connection_5__1__7_, 
        connection_5__1__6_, connection_5__1__5_, connection_5__1__4_, 
        connection_5__1__3_, connection_5__1__2_, connection_5__1__1_, 
        connection_5__1__0_, connection_5__0__31_, connection_5__0__30_, 
        connection_5__0__29_, connection_5__0__28_, connection_5__0__27_, 
        connection_5__0__26_, connection_5__0__25_, connection_5__0__24_, 
        connection_5__0__23_, connection_5__0__22_, connection_5__0__21_, 
        connection_5__0__20_, connection_5__0__19_, connection_5__0__18_, 
        connection_5__0__17_, connection_5__0__16_, connection_5__0__15_, 
        connection_5__0__14_, connection_5__0__13_, connection_5__0__12_, 
        connection_5__0__11_, connection_5__0__10_, connection_5__0__9_, 
        connection_5__0__8_, connection_5__0__7_, connection_5__0__6_, 
        connection_5__0__5_, connection_5__0__4_, connection_5__0__3_, 
        connection_5__0__2_, connection_5__0__1_, connection_5__0__0_}), 
        .o_valid({n549, n550}), .o_data_bus({n999, n1000, n1001, n1002, n1003, 
        n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, 
        n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, 
        n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, 
        n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, 
        n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, 
        n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062}), 
        .i_fwd_valid(fwd_connection_valid_sec_half[7]), .i_fwd_data_bus(
        fwd_connection_sec_half[255:224]), .o_fwd_valid(
        fwd_connection_valid_sec_half[3]), .o_fwd_data_bus(
        fwd_connection_sec_half[127:96]), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[39:35]) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_7 second_half_stages_6__sw_group_0__upper_group_1__upper_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_5__3_, 
        connection_valid_5__2_}), .i_data_bus({connection_5__3__31_, 
        connection_5__3__30_, connection_5__3__29_, connection_5__3__28_, 
        connection_5__3__27_, connection_5__3__26_, connection_5__3__25_, 
        connection_5__3__24_, connection_5__3__23_, connection_5__3__22_, 
        connection_5__3__21_, connection_5__3__20_, connection_5__3__19_, 
        connection_5__3__18_, connection_5__3__17_, connection_5__3__16_, 
        connection_5__3__15_, connection_5__3__14_, connection_5__3__13_, 
        connection_5__3__12_, connection_5__3__11_, connection_5__3__10_, 
        connection_5__3__9_, connection_5__3__8_, connection_5__3__7_, 
        connection_5__3__6_, connection_5__3__5_, connection_5__3__4_, 
        connection_5__3__3_, connection_5__3__2_, connection_5__3__1_, 
        connection_5__3__0_, connection_5__2__31_, connection_5__2__30_, 
        connection_5__2__29_, connection_5__2__28_, connection_5__2__27_, 
        connection_5__2__26_, connection_5__2__25_, connection_5__2__24_, 
        connection_5__2__23_, connection_5__2__22_, connection_5__2__21_, 
        connection_5__2__20_, connection_5__2__19_, connection_5__2__18_, 
        connection_5__2__17_, connection_5__2__16_, connection_5__2__15_, 
        connection_5__2__14_, connection_5__2__13_, connection_5__2__12_, 
        connection_5__2__11_, connection_5__2__10_, connection_5__2__9_, 
        connection_5__2__8_, connection_5__2__7_, connection_5__2__6_, 
        connection_5__2__5_, connection_5__2__4_, connection_5__2__3_, 
        connection_5__2__2_, connection_5__2__1_, connection_5__2__0_}), 
        .o_valid({n547, n548}), .o_data_bus({n935, n936, n937, n938, n939, 
        n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, 
        n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, 
        n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, 
        n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, 
        n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998}), 
        .i_fwd_valid(fwd_connection_valid_sec_half[6]), .i_fwd_data_bus(
        fwd_connection_sec_half[223:192]), .o_fwd_valid(
        fwd_connection_valid_sec_half[2]), .o_fwd_data_bus(
        fwd_connection_sec_half[95:64]), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[34:30]) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_6 second_half_stages_6__sw_group_0__upper_group_2__upper_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_5__5_, 
        connection_valid_5__4_}), .i_data_bus({connection_5__5__31_, 
        connection_5__5__30_, connection_5__5__29_, connection_5__5__28_, 
        connection_5__5__27_, connection_5__5__26_, connection_5__5__25_, 
        connection_5__5__24_, connection_5__5__23_, connection_5__5__22_, 
        connection_5__5__21_, connection_5__5__20_, connection_5__5__19_, 
        connection_5__5__18_, connection_5__5__17_, connection_5__5__16_, 
        connection_5__5__15_, connection_5__5__14_, connection_5__5__13_, 
        connection_5__5__12_, connection_5__5__11_, connection_5__5__10_, 
        connection_5__5__9_, connection_5__5__8_, connection_5__5__7_, 
        connection_5__5__6_, connection_5__5__5_, connection_5__5__4_, 
        connection_5__5__3_, connection_5__5__2_, connection_5__5__1_, 
        connection_5__5__0_, connection_5__4__31_, connection_5__4__30_, 
        connection_5__4__29_, connection_5__4__28_, connection_5__4__27_, 
        connection_5__4__26_, connection_5__4__25_, connection_5__4__24_, 
        connection_5__4__23_, connection_5__4__22_, connection_5__4__21_, 
        connection_5__4__20_, connection_5__4__19_, connection_5__4__18_, 
        connection_5__4__17_, connection_5__4__16_, connection_5__4__15_, 
        connection_5__4__14_, connection_5__4__13_, connection_5__4__12_, 
        connection_5__4__11_, connection_5__4__10_, connection_5__4__9_, 
        connection_5__4__8_, connection_5__4__7_, connection_5__4__6_, 
        connection_5__4__5_, connection_5__4__4_, connection_5__4__3_, 
        connection_5__4__2_, connection_5__4__1_, connection_5__4__0_}), 
        .o_valid({n545, n546}), .o_data_bus({n871, n872, n873, n874, n875, 
        n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, 
        n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, 
        n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, 
        n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, 
        n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934}), 
        .i_fwd_valid(fwd_connection_valid_sec_half[5]), .i_fwd_data_bus(
        fwd_connection_sec_half[191:160]), .o_fwd_valid(
        fwd_connection_valid_sec_half[1]), .o_fwd_data_bus(
        fwd_connection_sec_half[63:32]), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[29:25]) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_5 second_half_stages_6__sw_group_0__upper_group_3__upper_sw ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__7_, 
        connection_valid_5__6_}), .i_data_bus({connection_5__7__31_, 
        connection_5__7__30_, connection_5__7__29_, connection_5__7__28_, 
        connection_5__7__27_, connection_5__7__26_, connection_5__7__25_, 
        connection_5__7__24_, connection_5__7__23_, connection_5__7__22_, 
        connection_5__7__21_, connection_5__7__20_, connection_5__7__19_, 
        connection_5__7__18_, connection_5__7__17_, connection_5__7__16_, 
        connection_5__7__15_, connection_5__7__14_, connection_5__7__13_, 
        connection_5__7__12_, connection_5__7__11_, connection_5__7__10_, 
        connection_5__7__9_, connection_5__7__8_, connection_5__7__7_, 
        connection_5__7__6_, connection_5__7__5_, connection_5__7__4_, 
        connection_5__7__3_, connection_5__7__2_, connection_5__7__1_, 
        connection_5__7__0_, connection_5__6__31_, connection_5__6__30_, 
        connection_5__6__29_, connection_5__6__28_, connection_5__6__27_, 
        connection_5__6__26_, connection_5__6__25_, connection_5__6__24_, 
        connection_5__6__23_, connection_5__6__22_, connection_5__6__21_, 
        connection_5__6__20_, connection_5__6__19_, connection_5__6__18_, 
        connection_5__6__17_, connection_5__6__16_, connection_5__6__15_, 
        connection_5__6__14_, connection_5__6__13_, connection_5__6__12_, 
        connection_5__6__11_, connection_5__6__10_, connection_5__6__9_, 
        connection_5__6__8_, connection_5__6__7_, connection_5__6__6_, 
        connection_5__6__5_, connection_5__6__4_, connection_5__6__3_, 
        connection_5__6__2_, connection_5__6__1_, connection_5__6__0_}), 
        .o_valid({n543, n544}), .o_data_bus({n807, n808, n809, n810, n811, 
        n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, 
        n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, 
        n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, 
        n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, 
        n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870}), 
        .i_fwd_valid(fwd_connection_valid_sec_half[4]), .i_fwd_data_bus(
        fwd_connection_sec_half[159:128]), .o_fwd_valid(
        fwd_connection_valid_sec_half[0]), .o_fwd_data_bus(
        fwd_connection_sec_half[31:0]), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[24:20]) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_4 second_half_stages_6__sw_group_0__bottom_group_0__bottom_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_5__9_, 
        connection_valid_5__8_}), .i_data_bus({connection_5__9__31_, 
        connection_5__9__30_, connection_5__9__29_, connection_5__9__28_, 
        connection_5__9__27_, connection_5__9__26_, connection_5__9__25_, 
        connection_5__9__24_, connection_5__9__23_, connection_5__9__22_, 
        connection_5__9__21_, connection_5__9__20_, connection_5__9__19_, 
        connection_5__9__18_, connection_5__9__17_, connection_5__9__16_, 
        connection_5__9__15_, connection_5__9__14_, connection_5__9__13_, 
        connection_5__9__12_, connection_5__9__11_, connection_5__9__10_, 
        connection_5__9__9_, connection_5__9__8_, connection_5__9__7_, 
        connection_5__9__6_, connection_5__9__5_, connection_5__9__4_, 
        connection_5__9__3_, connection_5__9__2_, connection_5__9__1_, 
        connection_5__9__0_, connection_5__8__31_, connection_5__8__30_, 
        connection_5__8__29_, connection_5__8__28_, connection_5__8__27_, 
        connection_5__8__26_, connection_5__8__25_, connection_5__8__24_, 
        connection_5__8__23_, connection_5__8__22_, connection_5__8__21_, 
        connection_5__8__20_, connection_5__8__19_, connection_5__8__18_, 
        connection_5__8__17_, connection_5__8__16_, connection_5__8__15_, 
        connection_5__8__14_, connection_5__8__13_, connection_5__8__12_, 
        connection_5__8__11_, connection_5__8__10_, connection_5__8__9_, 
        connection_5__8__8_, connection_5__8__7_, connection_5__8__6_, 
        connection_5__8__5_, connection_5__8__4_, connection_5__8__3_, 
        connection_5__8__2_, connection_5__8__1_, connection_5__8__0_}), 
        .o_valid({n541, n542}), .o_data_bus({n743, n744, n745, n746, n747, 
        n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, 
        n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, 
        n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, 
        n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, 
        n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806}), 
        .i_fwd_valid(fwd_connection_valid_sec_half[3]), .i_fwd_data_bus(
        fwd_connection_sec_half[127:96]), .o_fwd_valid(
        fwd_connection_valid_sec_half[7]), .o_fwd_data_bus(
        fwd_connection_sec_half[255:224]), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[19:15]) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_3 second_half_stages_6__sw_group_0__bottom_group_1__bottom_sw ( 
        .clk(clk), .rst(n532), .i_valid({connection_valid_5__11_, 
        connection_valid_5__10_}), .i_data_bus({connection_5__11__31_, 
        connection_5__11__30_, connection_5__11__29_, connection_5__11__28_, 
        connection_5__11__27_, connection_5__11__26_, connection_5__11__25_, 
        connection_5__11__24_, connection_5__11__23_, connection_5__11__22_, 
        connection_5__11__21_, connection_5__11__20_, connection_5__11__19_, 
        connection_5__11__18_, connection_5__11__17_, connection_5__11__16_, 
        connection_5__11__15_, connection_5__11__14_, connection_5__11__13_, 
        connection_5__11__12_, connection_5__11__11_, connection_5__11__10_, 
        connection_5__11__9_, connection_5__11__8_, connection_5__11__7_, 
        connection_5__11__6_, connection_5__11__5_, connection_5__11__4_, 
        connection_5__11__3_, connection_5__11__2_, connection_5__11__1_, 
        connection_5__11__0_, connection_5__10__31_, connection_5__10__30_, 
        connection_5__10__29_, connection_5__10__28_, connection_5__10__27_, 
        connection_5__10__26_, connection_5__10__25_, connection_5__10__24_, 
        connection_5__10__23_, connection_5__10__22_, connection_5__10__21_, 
        connection_5__10__20_, connection_5__10__19_, connection_5__10__18_, 
        connection_5__10__17_, connection_5__10__16_, connection_5__10__15_, 
        connection_5__10__14_, connection_5__10__13_, connection_5__10__12_, 
        connection_5__10__11_, connection_5__10__10_, connection_5__10__9_, 
        connection_5__10__8_, connection_5__10__7_, connection_5__10__6_, 
        connection_5__10__5_, connection_5__10__4_, connection_5__10__3_, 
        connection_5__10__2_, connection_5__10__1_, connection_5__10__0_}), 
        .o_valid({n539, n540}), .o_data_bus({n679, n680, n681, n682, n683, 
        n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, 
        n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, 
        n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, 
        n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, 
        n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742}), 
        .i_fwd_valid(fwd_connection_valid_sec_half[2]), .i_fwd_data_bus(
        fwd_connection_sec_half[95:64]), .o_fwd_valid(
        fwd_connection_valid_sec_half[6]), .o_fwd_data_bus(
        fwd_connection_sec_half[223:192]), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[14:10]) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_2 second_half_stages_6__sw_group_0__bottom_group_2__bottom_sw ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__13_, 
        connection_valid_5__12_}), .i_data_bus({connection_5__13__31_, 
        connection_5__13__30_, connection_5__13__29_, connection_5__13__28_, 
        connection_5__13__27_, connection_5__13__26_, connection_5__13__25_, 
        connection_5__13__24_, connection_5__13__23_, connection_5__13__22_, 
        connection_5__13__21_, connection_5__13__20_, connection_5__13__19_, 
        connection_5__13__18_, connection_5__13__17_, connection_5__13__16_, 
        connection_5__13__15_, connection_5__13__14_, connection_5__13__13_, 
        connection_5__13__12_, connection_5__13__11_, connection_5__13__10_, 
        connection_5__13__9_, connection_5__13__8_, connection_5__13__7_, 
        connection_5__13__6_, connection_5__13__5_, connection_5__13__4_, 
        connection_5__13__3_, connection_5__13__2_, connection_5__13__1_, 
        connection_5__13__0_, connection_5__12__31_, connection_5__12__30_, 
        connection_5__12__29_, connection_5__12__28_, connection_5__12__27_, 
        connection_5__12__26_, connection_5__12__25_, connection_5__12__24_, 
        connection_5__12__23_, connection_5__12__22_, connection_5__12__21_, 
        connection_5__12__20_, connection_5__12__19_, connection_5__12__18_, 
        connection_5__12__17_, connection_5__12__16_, connection_5__12__15_, 
        connection_5__12__14_, connection_5__12__13_, connection_5__12__12_, 
        connection_5__12__11_, connection_5__12__10_, connection_5__12__9_, 
        connection_5__12__8_, connection_5__12__7_, connection_5__12__6_, 
        connection_5__12__5_, connection_5__12__4_, connection_5__12__3_, 
        connection_5__12__2_, connection_5__12__1_, connection_5__12__0_}), 
        .o_valid({n537, n538}), .o_data_bus({n615, n616, n617, n618, n619, 
        n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, 
        n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, 
        n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, 
        n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, 
        n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678}), 
        .i_fwd_valid(fwd_connection_valid_sec_half[1]), .i_fwd_data_bus(
        fwd_connection_sec_half[63:32]), .o_fwd_valid(
        fwd_connection_valid_sec_half[5]), .o_fwd_data_bus(
        fwd_connection_sec_half[191:160]), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[9:5]) );
  distribute_3x3_simple_seq_DATA_WIDTH32_COMMAND_WIDTH5_1 second_half_stages_6__sw_group_0__bottom_group_3__bottom_sw ( 
        .clk(clk), .rst(rst), .i_valid({connection_valid_5__15_, 
        connection_valid_5__14_}), .i_data_bus({connection_5__15__31_, 
        connection_5__15__30_, connection_5__15__29_, connection_5__15__28_, 
        connection_5__15__27_, connection_5__15__26_, connection_5__15__25_, 
        connection_5__15__24_, connection_5__15__23_, connection_5__15__22_, 
        connection_5__15__21_, connection_5__15__20_, connection_5__15__19_, 
        connection_5__15__18_, connection_5__15__17_, connection_5__15__16_, 
        connection_5__15__15_, connection_5__15__14_, connection_5__15__13_, 
        connection_5__15__12_, connection_5__15__11_, connection_5__15__10_, 
        connection_5__15__9_, connection_5__15__8_, connection_5__15__7_, 
        connection_5__15__6_, connection_5__15__5_, connection_5__15__4_, 
        connection_5__15__3_, connection_5__15__2_, connection_5__15__1_, 
        connection_5__15__0_, connection_5__14__31_, connection_5__14__30_, 
        connection_5__14__29_, connection_5__14__28_, connection_5__14__27_, 
        connection_5__14__26_, connection_5__14__25_, connection_5__14__24_, 
        connection_5__14__23_, connection_5__14__22_, connection_5__14__21_, 
        connection_5__14__20_, connection_5__14__19_, connection_5__14__18_, 
        connection_5__14__17_, connection_5__14__16_, connection_5__14__15_, 
        connection_5__14__14_, connection_5__14__13_, connection_5__14__12_, 
        connection_5__14__11_, connection_5__14__10_, connection_5__14__9_, 
        connection_5__14__8_, connection_5__14__7_, connection_5__14__6_, 
        connection_5__14__5_, connection_5__14__4_, connection_5__14__3_, 
        connection_5__14__2_, connection_5__14__1_, connection_5__14__0_}), 
        .o_valid({n535, n536}), .o_data_bus({n551, n552, n553, n554, n555, 
        n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, 
        n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, 
        n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, 
        n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, 
        n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614}), 
        .i_fwd_valid(fwd_connection_valid_sec_half[0]), .i_fwd_data_bus(
        fwd_connection_sec_half[31:0]), .o_fwd_valid(
        fwd_connection_valid_sec_half[4]), .o_fwd_data_bus(
        fwd_connection_sec_half[159:128]), .i_en(i_en), .i_cmd(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[4:0]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__0__4_ ( 
        .D(i_cmd[44]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__0__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__0__3_ ( 
        .D(i_cmd[43]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__0__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__0__2_ ( 
        .D(i_cmd[42]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__0__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__0__1_ ( 
        .D(i_cmd[41]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__0__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__0__0_ ( 
        .D(i_cmd[40]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__0__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__1__4_ ( 
        .D(i_cmd[49]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__1__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__1__3_ ( 
        .D(i_cmd[48]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__1__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__1__2_ ( 
        .D(i_cmd[47]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__1__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__1__1_ ( 
        .D(i_cmd[46]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__1__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__1__0_ ( 
        .D(i_cmd[45]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__1__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__2__4_ ( 
        .D(i_cmd[54]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__2__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__2__3_ ( 
        .D(i_cmd[53]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__2__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__2__2_ ( 
        .D(i_cmd[52]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__2__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__2__1_ ( 
        .D(i_cmd[51]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__2__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__2__0_ ( 
        .D(i_cmd[50]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__2__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__3__4_ ( 
        .D(i_cmd[59]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__3__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__3__3_ ( 
        .D(i_cmd[58]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__3__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__3__2_ ( 
        .D(i_cmd[57]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__3__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__3__1_ ( 
        .D(i_cmd[56]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__3__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__3__0_ ( 
        .D(i_cmd[55]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__3__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__4__4_ ( 
        .D(i_cmd[64]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__4__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__4__3_ ( 
        .D(i_cmd[63]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__4__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__4__2_ ( 
        .D(i_cmd[62]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__4__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__4__1_ ( 
        .D(i_cmd[61]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__4__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__4__0_ ( 
        .D(i_cmd[60]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__4__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__5__4_ ( 
        .D(i_cmd[69]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__5__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__5__3_ ( 
        .D(i_cmd[68]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__5__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__5__2_ ( 
        .D(i_cmd[67]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__5__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__5__1_ ( 
        .D(i_cmd[66]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__5__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__5__0_ ( 
        .D(i_cmd[65]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__5__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__6__4_ ( 
        .D(i_cmd[74]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__6__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__6__3_ ( 
        .D(i_cmd[73]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__6__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__6__2_ ( 
        .D(i_cmd[72]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__6__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__6__1_ ( 
        .D(i_cmd[71]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__6__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__6__0_ ( 
        .D(i_cmd[70]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__6__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__7__4_ ( 
        .D(i_cmd[79]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__7__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__7__3_ ( 
        .D(i_cmd[78]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__7__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__7__2_ ( 
        .D(i_cmd[77]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__7__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__7__1_ ( 
        .D(i_cmd[76]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__7__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_0__7__0_ ( 
        .D(i_cmd[75]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_0__7__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__0__4_ ( 
        .D(i_cmd[84]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__0__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__0__3_ ( 
        .D(i_cmd[83]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__0__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__0__2_ ( 
        .D(i_cmd[82]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__0__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__0__1_ ( 
        .D(i_cmd[81]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__0__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__0__0_ ( 
        .D(i_cmd[80]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__0__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__1__4_ ( 
        .D(i_cmd[89]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__1__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__1__3_ ( 
        .D(i_cmd[88]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__1__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__1__2_ ( 
        .D(i_cmd[87]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__1__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__1__1_ ( 
        .D(i_cmd[86]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__1__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__1__0_ ( 
        .D(i_cmd[85]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__1__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__2__4_ ( 
        .D(i_cmd[94]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__2__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__2__3_ ( 
        .D(i_cmd[93]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__2__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__2__2_ ( 
        .D(i_cmd[92]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__2__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__2__1_ ( 
        .D(i_cmd[91]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__2__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__2__0_ ( 
        .D(i_cmd[90]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__2__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__3__4_ ( 
        .D(i_cmd[99]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__3__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__3__3_ ( 
        .D(i_cmd[98]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__3__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__3__2_ ( 
        .D(i_cmd[97]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__3__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__3__1_ ( 
        .D(i_cmd[96]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__3__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__3__0_ ( 
        .D(i_cmd[95]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__3__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__4__4_ ( 
        .D(i_cmd[104]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__4__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__4__3_ ( 
        .D(i_cmd[103]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__4__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__4__2_ ( 
        .D(i_cmd[102]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__4__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__4__1_ ( 
        .D(i_cmd[101]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__4__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__4__0_ ( 
        .D(i_cmd[100]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__4__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__5__4_ ( 
        .D(i_cmd[109]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__5__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__5__3_ ( 
        .D(i_cmd[108]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__5__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__5__2_ ( 
        .D(i_cmd[107]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__5__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__5__1_ ( 
        .D(i_cmd[106]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__5__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__5__0_ ( 
        .D(i_cmd[105]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__5__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__6__4_ ( 
        .D(i_cmd[114]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__6__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__6__3_ ( 
        .D(i_cmd[113]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__6__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__6__2_ ( 
        .D(i_cmd[112]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__6__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__6__1_ ( 
        .D(i_cmd[111]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__6__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__6__0_ ( 
        .D(i_cmd[110]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__6__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__7__4_ ( 
        .D(i_cmd[119]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__7__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__7__3_ ( 
        .D(i_cmd[118]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__7__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__7__2_ ( 
        .D(i_cmd[117]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__7__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__7__1_ ( 
        .D(i_cmd[116]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__7__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_1__7__0_ ( 
        .D(i_cmd[115]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__7__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__0__1_ ( 
        .D(i_cmd[121]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__0__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__0__0_ ( 
        .D(i_cmd[120]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__0__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__1__1_ ( 
        .D(i_cmd[126]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__1__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__1__0_ ( 
        .D(i_cmd[125]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__1__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__2__1_ ( 
        .D(i_cmd[131]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__2__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__2__0_ ( 
        .D(i_cmd[130]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__2__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__3__1_ ( 
        .D(i_cmd[136]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__3__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__3__0_ ( 
        .D(i_cmd[135]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__3__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__4__1_ ( 
        .D(i_cmd[141]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__4__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__4__0_ ( 
        .D(i_cmd[140]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__4__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__5__1_ ( 
        .D(i_cmd[146]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__5__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__5__0_ ( 
        .D(i_cmd[145]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__5__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__6__1_ ( 
        .D(i_cmd[151]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__6__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__6__0_ ( 
        .D(i_cmd[150]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__6__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__7__1_ ( 
        .D(i_cmd[156]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__7__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_2__7__0_ ( 
        .D(i_cmd[155]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__7__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__0__4_ ( 
        .D(i_cmd[164]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__0__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__0__3_ ( 
        .D(i_cmd[163]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__0__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__0__2_ ( 
        .D(i_cmd[162]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__0__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__0__1_ ( 
        .D(i_cmd[161]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__0__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__0__0_ ( 
        .D(i_cmd[160]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__0__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__1__4_ ( 
        .D(i_cmd[169]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__1__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__1__3_ ( 
        .D(i_cmd[168]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__1__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__1__2_ ( 
        .D(i_cmd[167]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__1__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__1__1_ ( 
        .D(i_cmd[166]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__1__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__1__0_ ( 
        .D(i_cmd[165]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__1__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__2__4_ ( 
        .D(i_cmd[174]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__2__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__2__3_ ( 
        .D(i_cmd[173]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__2__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__2__2_ ( 
        .D(i_cmd[172]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__2__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__2__1_ ( 
        .D(i_cmd[171]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__2__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__2__0_ ( 
        .D(i_cmd[170]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__2__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__3__4_ ( 
        .D(i_cmd[179]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__3__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__3__3_ ( 
        .D(i_cmd[178]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__3__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__3__2_ ( 
        .D(i_cmd[177]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__3__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__3__1_ ( 
        .D(i_cmd[176]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__3__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__3__0_ ( 
        .D(i_cmd[175]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__3__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__4__4_ ( 
        .D(i_cmd[184]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__4__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__4__3_ ( 
        .D(i_cmd[183]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__4__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__4__2_ ( 
        .D(i_cmd[182]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__4__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__4__1_ ( 
        .D(i_cmd[181]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__4__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__4__0_ ( 
        .D(i_cmd[180]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__4__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__5__4_ ( 
        .D(i_cmd[189]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__5__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__5__3_ ( 
        .D(i_cmd[188]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__5__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__5__2_ ( 
        .D(i_cmd[187]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__5__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__5__1_ ( 
        .D(i_cmd[186]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__5__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__5__0_ ( 
        .D(i_cmd[185]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__5__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__6__4_ ( 
        .D(i_cmd[194]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__6__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__6__3_ ( 
        .D(i_cmd[193]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__6__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__6__2_ ( 
        .D(i_cmd[192]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__6__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__6__1_ ( 
        .D(i_cmd[191]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__6__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__6__0_ ( 
        .D(i_cmd[190]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__6__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__7__4_ ( 
        .D(i_cmd[199]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__7__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__7__3_ ( 
        .D(i_cmd[198]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__7__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__7__2_ ( 
        .D(i_cmd[197]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__7__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__7__1_ ( 
        .D(i_cmd[196]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__7__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_3__7__0_ ( 
        .D(i_cmd[195]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__7__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__0__4_ ( 
        .D(i_cmd[204]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__0__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__0__3_ ( 
        .D(i_cmd[203]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__0__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__0__2_ ( 
        .D(i_cmd[202]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__0__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__0__1_ ( 
        .D(i_cmd[201]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__0__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__0__0_ ( 
        .D(i_cmd[200]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__0__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__1__4_ ( 
        .D(i_cmd[209]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__1__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__1__3_ ( 
        .D(i_cmd[208]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__1__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__1__2_ ( 
        .D(i_cmd[207]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__1__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__1__1_ ( 
        .D(i_cmd[206]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__1__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__1__0_ ( 
        .D(i_cmd[205]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__1__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__2__4_ ( 
        .D(i_cmd[214]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__2__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__2__3_ ( 
        .D(i_cmd[213]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__2__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__2__2_ ( 
        .D(i_cmd[212]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__2__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__2__1_ ( 
        .D(i_cmd[211]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__2__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__2__0_ ( 
        .D(i_cmd[210]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__2__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__3__4_ ( 
        .D(i_cmd[219]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__3__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__3__3_ ( 
        .D(i_cmd[218]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__3__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__3__2_ ( 
        .D(i_cmd[217]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__3__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__3__1_ ( 
        .D(i_cmd[216]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__3__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__3__0_ ( 
        .D(i_cmd[215]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__3__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__4__4_ ( 
        .D(i_cmd[224]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__4__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__4__3_ ( 
        .D(i_cmd[223]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__4__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__4__2_ ( 
        .D(i_cmd[222]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__4__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__4__1_ ( 
        .D(i_cmd[221]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__4__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__4__0_ ( 
        .D(i_cmd[220]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__4__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__5__4_ ( 
        .D(i_cmd[229]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__5__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__5__3_ ( 
        .D(i_cmd[228]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__5__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__5__2_ ( 
        .D(i_cmd[227]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__5__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__5__1_ ( 
        .D(i_cmd[226]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__5__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__5__0_ ( 
        .D(i_cmd[225]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__5__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__6__4_ ( 
        .D(i_cmd[234]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__6__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__6__3_ ( 
        .D(i_cmd[233]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__6__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__6__2_ ( 
        .D(i_cmd[232]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__6__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__6__1_ ( 
        .D(i_cmd[231]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__6__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__6__0_ ( 
        .D(i_cmd[230]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__6__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__7__4_ ( 
        .D(i_cmd[239]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__7__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__7__3_ ( 
        .D(i_cmd[238]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__7__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__7__2_ ( 
        .D(i_cmd[237]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__7__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__7__1_ ( 
        .D(i_cmd[236]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__7__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_4__7__0_ ( 
        .D(i_cmd[235]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__7__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__0__4_ ( 
        .D(i_cmd[244]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__0__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__0__3_ ( 
        .D(i_cmd[243]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__0__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__0__2_ ( 
        .D(i_cmd[242]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__0__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__0__1_ ( 
        .D(i_cmd[241]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__0__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__0__0_ ( 
        .D(i_cmd[240]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__0__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__1__4_ ( 
        .D(i_cmd[249]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__1__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__1__3_ ( 
        .D(i_cmd[248]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__1__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__1__2_ ( 
        .D(i_cmd[247]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__1__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__1__1_ ( 
        .D(i_cmd[246]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__1__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__1__0_ ( 
        .D(i_cmd[245]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__1__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__2__4_ ( 
        .D(i_cmd[254]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__2__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__2__3_ ( 
        .D(i_cmd[253]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__2__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__2__2_ ( 
        .D(i_cmd[252]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__2__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__2__1_ ( 
        .D(i_cmd[251]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__2__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__2__0_ ( 
        .D(i_cmd[250]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__2__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__3__4_ ( 
        .D(i_cmd[259]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__3__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__3__3_ ( 
        .D(i_cmd[258]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__3__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__3__2_ ( 
        .D(i_cmd[257]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__3__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__3__1_ ( 
        .D(i_cmd[256]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__3__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__3__0_ ( 
        .D(i_cmd[255]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__3__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__4__4_ ( 
        .D(i_cmd[264]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__4__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__4__3_ ( 
        .D(i_cmd[263]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__4__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__4__2_ ( 
        .D(i_cmd[262]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__4__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__4__1_ ( 
        .D(i_cmd[261]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__4__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__4__0_ ( 
        .D(i_cmd[260]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__4__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__5__4_ ( 
        .D(i_cmd[269]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__5__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__5__3_ ( 
        .D(i_cmd[268]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__5__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__5__2_ ( 
        .D(i_cmd[267]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__5__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__5__1_ ( 
        .D(i_cmd[266]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__5__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__5__0_ ( 
        .D(i_cmd[265]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__5__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__6__4_ ( 
        .D(i_cmd[274]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__6__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__6__3_ ( 
        .D(i_cmd[273]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__6__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__6__2_ ( 
        .D(i_cmd[272]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__6__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__6__1_ ( 
        .D(i_cmd[271]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__6__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__6__0_ ( 
        .D(i_cmd[270]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__6__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__7__4_ ( 
        .D(i_cmd[279]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__7__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__7__3_ ( 
        .D(i_cmd[278]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__7__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__7__2_ ( 
        .D(i_cmd[277]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__7__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__7__1_ ( 
        .D(i_cmd[276]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__7__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_0__pipeline_i_cmd_reg_reg_5__7__0_ ( 
        .D(i_cmd[275]), .CP(clk), .Q(
        cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__7__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__0__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__0__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__0__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__0__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__0__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__0__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__0__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__0__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__0__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__0__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__0__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__0__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__0__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__0__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__0__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__1__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__1__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__1__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__1__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__1__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__1__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__1__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__1__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__1__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__1__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__1__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__1__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__1__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__1__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__1__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__2__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__2__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__2__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__2__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__2__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__2__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__2__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__2__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__2__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__2__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__2__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__2__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__2__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__2__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__2__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__3__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__3__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__3__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__3__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__3__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__3__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__3__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__3__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__3__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__3__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__3__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__3__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__3__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__3__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__3__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__4__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__4__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__4__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__4__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__4__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__4__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__4__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__4__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__4__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__4__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__4__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__4__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__4__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__4__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__4__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__5__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__5__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__5__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__5__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__5__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__5__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__5__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__5__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__5__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__5__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__5__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__5__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__5__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__5__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__5__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__6__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__6__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__6__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__6__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__6__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__6__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__6__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__6__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__6__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__6__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__6__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__6__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__6__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__6__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__6__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__7__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__7__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__7__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__7__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__7__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__7__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__7__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__7__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__7__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__7__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__7__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__7__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_0__7__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_1__7__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_0__7__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__0__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__0__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__0__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__0__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__0__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__0__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__1__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__1__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__1__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__1__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__1__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__1__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__2__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__2__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__2__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__2__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__2__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__2__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__3__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__3__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__3__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__3__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__3__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__3__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__4__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__4__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__4__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__4__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__4__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__4__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__5__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__5__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__5__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__5__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__5__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__5__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__6__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__6__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__6__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__6__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__6__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__6__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__7__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__7__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__7__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_1__7__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_2__7__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__7__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__0__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__0__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__0__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__0__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__0__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__0__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__0__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__0__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__0__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__0__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__0__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__0__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__0__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__0__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__0__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__1__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__1__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__1__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__1__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__1__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__1__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__1__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__1__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__1__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__1__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__1__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__1__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__1__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__1__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__1__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__2__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__2__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__2__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__2__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__2__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__2__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__2__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__2__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__2__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__2__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__2__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__2__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__2__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__2__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__2__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__3__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__3__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__3__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__3__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__3__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__3__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__3__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__3__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__3__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__3__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__3__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__3__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__3__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__3__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__3__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__4__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__4__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__4__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__4__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__4__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__4__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__4__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__4__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__4__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__4__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__4__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__4__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__4__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__4__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__4__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__5__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__5__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__5__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__5__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__5__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__5__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__5__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__5__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__5__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__5__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__5__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__5__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__5__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__5__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__5__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__6__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__6__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__6__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__6__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__6__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__6__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__6__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__6__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__6__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__6__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__6__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__6__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__6__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__6__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__6__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__7__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__7__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__7__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__7__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__7__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__7__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__7__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__7__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__7__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__7__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__7__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__7__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_2__7__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_3__7__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__7__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__0__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__0__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__0__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__0__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__0__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__0__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__0__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__0__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__0__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__0__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__0__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__0__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__0__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__0__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__0__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__1__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__1__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__1__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__1__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__1__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__1__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__1__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__1__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__1__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__1__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__1__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__1__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__1__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__1__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__1__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__2__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__2__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__2__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__2__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__2__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__2__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__2__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__2__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__2__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__2__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__2__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__2__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__2__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__2__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__2__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__3__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__3__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__3__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__3__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__3__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__3__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__3__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__3__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__3__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__3__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__3__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__3__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__3__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__3__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__3__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__4__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__4__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__4__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__4__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__4__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__4__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__4__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__4__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__4__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__4__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__4__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__4__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__4__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__4__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__4__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__5__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__5__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__5__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__5__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__5__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__5__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__5__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__5__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__5__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__5__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__5__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__5__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__5__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__5__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__5__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__6__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__6__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__6__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__6__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__6__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__6__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__6__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__6__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__6__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__6__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__6__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__6__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__6__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__6__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__6__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__7__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__7__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__7__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__7__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__7__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__7__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__7__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__7__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__7__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__7__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__7__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__7__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_3__7__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_4__7__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__7__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__0__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__0__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__0__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__0__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__0__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__0__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__0__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__0__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__0__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__0__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__0__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__0__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__0__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__0__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__0__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__1__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__1__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__1__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__1__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__1__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__1__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__1__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__1__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__1__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__1__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__1__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__1__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__1__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__1__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__1__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__2__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__2__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__2__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__2__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__2__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__2__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__2__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__2__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__2__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__2__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__2__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__2__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__2__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__2__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__2__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__3__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__3__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__3__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__3__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__3__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__3__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__3__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__3__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__3__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__3__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__3__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__3__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__3__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__3__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__3__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__4__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__4__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__4__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__4__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__4__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__4__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__4__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__4__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__4__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__4__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__4__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__4__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__4__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__4__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__4__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__5__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__5__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__5__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__5__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__5__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__5__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__5__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__5__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__5__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__5__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__5__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__5__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__5__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__5__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__5__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__6__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__6__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__6__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__6__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__6__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__6__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__6__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__6__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__6__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__6__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__6__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__6__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__6__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__6__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__6__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__7__4_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__7__4_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__7__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__7__3_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__7__3_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__7__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__7__2_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__7__2_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__7__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__7__1_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__7__1_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__7__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_1__pipeline_i_cmd_reg_reg_4__7__0_ ( 
        .D(cmd_pipeline_stage_0__pipeline_i_cmd_reg_5__7__0_), .CP(clk), .Q(
        cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__7__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__0__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__0__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__0__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__0__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__0__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__0__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__1__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__1__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__1__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__1__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__1__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__1__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__2__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__2__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__2__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__2__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__2__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__2__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__3__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__3__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__3__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__3__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__3__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__3__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__4__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__4__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__4__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__4__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__4__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__4__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__5__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__5__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__5__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__5__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__5__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__5__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__6__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__6__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__6__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__6__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__6__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__6__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__7__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__7__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__7__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_0__7__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_1__7__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_0__7__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__0__4_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__0__4_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__0__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__0__3_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__0__3_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__0__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__0__2_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__0__2_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__0__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__0__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__0__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__0__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__0__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__0__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__0__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__1__4_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__1__4_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__1__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__1__3_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__1__3_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__1__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__1__2_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__1__2_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__1__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__1__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__1__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__1__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__1__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__1__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__1__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__2__4_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__2__4_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__2__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__2__3_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__2__3_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__2__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__2__2_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__2__2_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__2__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__2__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__2__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__2__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__2__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__2__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__2__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__3__4_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__3__4_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__3__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__3__3_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__3__3_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__3__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__3__2_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__3__2_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__3__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__3__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__3__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__3__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__3__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__3__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__3__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__4__4_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__4__4_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__4__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__4__3_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__4__3_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__4__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__4__2_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__4__2_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__4__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__4__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__4__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__4__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__4__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__4__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__4__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__5__4_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__5__4_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__5__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__5__3_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__5__3_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__5__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__5__2_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__5__2_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__5__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__5__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__5__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__5__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__5__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__5__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__5__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__6__4_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__6__4_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__6__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__6__3_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__6__3_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__6__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__6__2_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__6__2_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__6__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__6__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__6__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__6__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__6__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__6__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__6__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__7__4_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__7__4_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__7__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__7__3_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__7__3_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__7__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__7__2_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__7__2_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__7__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__7__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__7__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__7__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_1__7__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_2__7__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__7__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__0__4_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__0__4_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__0__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__0__3_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__0__3_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__0__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__0__2_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__0__2_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__0__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__0__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__0__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__0__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__0__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__0__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__0__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__1__4_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__1__4_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__1__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__1__3_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__1__3_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__1__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__1__2_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__1__2_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__1__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__1__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__1__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__1__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__1__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__1__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__1__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__2__4_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__2__4_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__2__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__2__3_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__2__3_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__2__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__2__2_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__2__2_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__2__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__2__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__2__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__2__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__2__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__2__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__2__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__3__4_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__3__4_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__3__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__3__3_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__3__3_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__3__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__3__2_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__3__2_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__3__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__3__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__3__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__3__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__3__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__3__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__3__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__4__4_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__4__4_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__4__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__4__3_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__4__3_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__4__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__4__2_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__4__2_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__4__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__4__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__4__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__4__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__4__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__4__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__4__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__5__4_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__5__4_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__5__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__5__3_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__5__3_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__5__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__5__2_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__5__2_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__5__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__5__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__5__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__5__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__5__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__5__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__5__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__6__4_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__6__4_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__6__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__6__3_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__6__3_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__6__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__6__2_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__6__2_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__6__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__6__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__6__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__6__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__6__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__6__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__6__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__7__4_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__7__4_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__7__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__7__3_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__7__3_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__7__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__7__2_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__7__2_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__7__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__7__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__7__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__7__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_2__7__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_3__7__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__7__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__0__4_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__0__4_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__0__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__0__3_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__0__3_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__0__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__0__2_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__0__2_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__0__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__0__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__0__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__0__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__0__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__0__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__0__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__1__4_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__1__4_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__1__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__1__3_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__1__3_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__1__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__1__2_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__1__2_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__1__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__1__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__1__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__1__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__1__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__1__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__1__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__2__4_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__2__4_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__2__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__2__3_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__2__3_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__2__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__2__2_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__2__2_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__2__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__2__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__2__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__2__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__2__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__2__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__2__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__3__4_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__3__4_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__3__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__3__3_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__3__3_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__3__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__3__2_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__3__2_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__3__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__3__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__3__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__3__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__3__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__3__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__3__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__4__4_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__4__4_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__4__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__4__3_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__4__3_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__4__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__4__2_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__4__2_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__4__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__4__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__4__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__4__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__4__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__4__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__4__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__5__4_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__5__4_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__5__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__5__3_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__5__3_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__5__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__5__2_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__5__2_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__5__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__5__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__5__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__5__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__5__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__5__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__5__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__6__4_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__6__4_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__6__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__6__3_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__6__3_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__6__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__6__2_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__6__2_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__6__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__6__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__6__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__6__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__6__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__6__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__6__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__7__4_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__7__4_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__7__4_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__7__3_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__7__3_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__7__3_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__7__2_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__7__2_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__7__2_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__7__1_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__7__1_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__7__1_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_2__pipeline_i_cmd_reg_reg_3__7__0_ ( 
        .D(cmd_pipeline_stage_1__pipeline_i_cmd_reg_4__7__0_), .CP(clk), .Q(
        cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__7__0_) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__0__4_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__0__4_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[119]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__0__3_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__0__3_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[118]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__0__2_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__0__2_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[117]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__0__1_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__0__1_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[116]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__0__0_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__0__0_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[115]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__1__4_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__1__4_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[114]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__1__3_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__1__3_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[113]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__1__2_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__1__2_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[112]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__1__1_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__1__1_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[111]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__1__0_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__1__0_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[110]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__2__4_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__2__4_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[109]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__2__3_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__2__3_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[108]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__2__2_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__2__2_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[107]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__2__0_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__2__0_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[105]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__3__2_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__3__2_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[102]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__4__4_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__4__4_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[99]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__4__3_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__4__3_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[98]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__4__2_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__4__2_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[97]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__4__1_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__4__1_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[96]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__4__0_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__4__0_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[95]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__5__4_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__5__4_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[94]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__5__3_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__5__3_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[93]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__5__2_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__5__2_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[92]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__5__1_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__5__1_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[91]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__5__0_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__5__0_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[90]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__6__4_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__6__4_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[89]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__6__3_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__6__3_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[88]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__6__2_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__6__2_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[87]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__6__0_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__6__0_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[85]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__7__4_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__7__4_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[84]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__7__3_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__7__3_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[83]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__7__2_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__7__2_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[82]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__0__4_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__0__4_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[79]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__0__3_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__0__3_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[78]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__0__2_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__0__2_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[77]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__0__1_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__0__1_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[76]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__0__0_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__0__0_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[75]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__1__4_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__1__4_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[74]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__1__3_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__1__3_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[73]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__1__2_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__1__2_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[72]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__1__1_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__1__1_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[71]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__1__0_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__1__0_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[70]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__2__4_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__2__4_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[69]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__2__3_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__2__3_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[68]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__2__2_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__2__2_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[67]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__2__1_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__2__1_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[66]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__2__0_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__2__0_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[65]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__3__4_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__3__4_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[64]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__3__3_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__3__3_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[63]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__3__2_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__3__2_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[62]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__3__1_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__3__1_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[61]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__3__0_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__3__0_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[60]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__4__4_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__4__4_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[59]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__4__3_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__4__3_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[58]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__4__2_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__4__2_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[57]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__4__1_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__4__1_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[56]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__4__0_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__4__0_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[55]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__5__4_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__5__4_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[54]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__5__3_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__5__3_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[53]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__5__2_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__5__2_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[52]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__5__1_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__5__1_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[51]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__5__0_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__5__0_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[50]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__6__4_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__6__4_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[49]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__6__3_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__6__3_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[48]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__6__2_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__6__2_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[47]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__6__1_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__6__1_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[46]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__6__0_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__6__0_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[45]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__7__4_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__7__4_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[44]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__7__3_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__7__3_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[43]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__7__2_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__7__2_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[42]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__7__1_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__7__1_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[41]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_1__7__0_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_2__7__0_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[40]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__0__4_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__0__4_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[39]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__0__3_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__0__3_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[38]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__0__2_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__0__2_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[37]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__0__1_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__0__1_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[36]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__0__0_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__0__0_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[35]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__1__4_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__1__4_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[34]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__1__3_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__1__3_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[33]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__1__2_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__1__2_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[32]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__1__1_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__1__1_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[31]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__1__0_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__1__0_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[30]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__2__4_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__2__4_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[29]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__2__3_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__2__3_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[28]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__2__2_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__2__2_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[27]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__2__1_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__2__1_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[26]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__2__0_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__2__0_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[25]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__3__4_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__3__4_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[24]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__3__3_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__3__3_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[23]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__3__2_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__3__2_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[22]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__3__1_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__3__1_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[21]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__3__0_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__3__0_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[20]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__4__4_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__4__4_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[19]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__4__3_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__4__3_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[18]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__4__2_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__4__2_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[17]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__4__1_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__4__1_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[16]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__4__0_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__4__0_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[15]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__5__4_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__5__4_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[14]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__5__3_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__5__3_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[13]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__5__2_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__5__2_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[12]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__5__1_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__5__1_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[11]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__5__0_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__5__0_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[10]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__6__4_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__6__4_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[9]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__6__3_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__6__3_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[8]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__6__2_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__6__2_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__6__1_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__6__1_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__6__0_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__6__0_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__7__4_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__7__4_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__7__3_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__7__3_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__7__2_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__7__2_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__7__1_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__7__1_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_2__7__0_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_3__7__0_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__0__4_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[79]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[79]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__0__3_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[78]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[78]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__0__1_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[76]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[76]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__0__0_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[75]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[75]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__1__4_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[74]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[74]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__1__3_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[73]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[73]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__1__2_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[72]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[72]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__1__1_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[71]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[71]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__1__0_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[70]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[70]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__2__4_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[69]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[69]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__2__3_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[68]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[68]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__2__2_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[67]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[67]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__2__1_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[66]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[66]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__2__0_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[65]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[65]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__3__4_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[64]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[64]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__3__3_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[63]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[63]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__3__2_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[62]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[62]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__3__1_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[61]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[61]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__3__0_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[60]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[60]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__4__4_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[59]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[59]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__4__2_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[57]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[57]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__4__1_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[56]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[56]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__4__0_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[55]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[55]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__5__4_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[54]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[54]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__5__3_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[53]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[53]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__5__2_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[52]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[52]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__5__1_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[51]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[51]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__5__0_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[50]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[50]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__6__4_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[49]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[49]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__6__3_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[48]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[48]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__6__2_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[47]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[47]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__6__1_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[46]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[46]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__6__0_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[45]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[45]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__7__4_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[44]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[44]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__7__3_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[43]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[43]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__7__2_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[42]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[42]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__7__1_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[41]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[41]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__7__0_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[40]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[40]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__0__4_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[39]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[39]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__0__3_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[38]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[38]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__0__2_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[37]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[37]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__0__1_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[36]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[36]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__0__0_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[35]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[35]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__1__4_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[34]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[34]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__1__3_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[33]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[33]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__1__2_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[32]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[32]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__1__1_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[31]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[31]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__1__0_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[30]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[30]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__2__4_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[29]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[29]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__2__3_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[28]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[28]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__2__2_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[27]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[27]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__2__1_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[26]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[26]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__2__0_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[25]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[25]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__3__4_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[24]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[24]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__3__3_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[23]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[23]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__3__2_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[22]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[22]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__3__1_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[21]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[21]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__3__0_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[20]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[20]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__4__4_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[19]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[19]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__4__3_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[18]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[18]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__4__2_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[17]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[17]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__4__1_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[16]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[16]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__4__0_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[15]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[15]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__5__4_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[14]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[14]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__5__3_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[13]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[13]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__5__2_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[12]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[12]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__5__1_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[11]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[11]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__5__0_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[10]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[10]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__6__4_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[9]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[9]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__6__3_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[8]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[8]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__6__2_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[7]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__6__1_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[6]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__6__0_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[5]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__7__4_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[4]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__7__3_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[3]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__7__2_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[2]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__7__1_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[1]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_1__7__0_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[0]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__0__4_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[39]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[39]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__0__3_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[38]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[38]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__0__2_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[37]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[37]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__0__1_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[36]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[36]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__0__0_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[35]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[35]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__1__4_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[34]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[34]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__1__3_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[33]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[33]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__1__2_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[32]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[32]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__1__1_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[31]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[31]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__1__0_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[30]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[30]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__2__4_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[29]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[29]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__2__3_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[28]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[28]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__2__2_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[27]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[27]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__2__1_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[26]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[26]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__2__0_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[25]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[25]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__3__4_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[24]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[24]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__3__3_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[23]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[23]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__3__2_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[22]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[22]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__3__1_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[21]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[21]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__3__0_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[20]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[20]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__4__4_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[19]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[19]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__4__3_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[18]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[18]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__4__2_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[17]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[17]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__4__1_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[16]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[16]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__4__0_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[15]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[15]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__5__4_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[14]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[14]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__5__3_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[13]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[13]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__5__2_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[12]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[12]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__5__1_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[11]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[11]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__5__0_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[10]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[10]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__6__3_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[8]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[8]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__6__2_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[7]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__6__1_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[6]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__6__0_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[5]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__7__4_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[4]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__7__3_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[3]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__7__2_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[2]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__7__1_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[1]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__7__0_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[0]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__6__1_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__6__1_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[86]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__3__1_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__3__1_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[101]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__3__0_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__3__0_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[100]) );
  DFQD2BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__2__1_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__2__1_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[106]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__0__2_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[77]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[77]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_4__pipeline_i_cmd_reg_reg_0__4__3_ ( 
        .D(cmd_pipeline_stage_3__pipeline_i_cmd_reg[58]), .CP(clk), .Q(
        cmd_pipeline_stage_4__pipeline_i_cmd_reg[58]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_5__pipeline_i_cmd_reg_reg_0__6__4_ ( 
        .D(cmd_pipeline_stage_4__pipeline_i_cmd_reg[9]), .CP(clk), .Q(
        cmd_pipeline_stage_5__pipeline_i_cmd_reg[9]) );
  DFQD2BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__7__0_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__7__0_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[80]) );
  DFQD2BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__7__1_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__7__1_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[81]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__3__3_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__3__3_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[103]) );
  DFQD1BWP30P140LVT cmd_pipeline_stage_3__pipeline_i_cmd_reg_reg_0__3__4_ ( 
        .D(cmd_pipeline_stage_2__pipeline_i_cmd_reg_1__3__4_), .CP(clk), .Q(
        cmd_pipeline_stage_3__pipeline_i_cmd_reg[104]) );
  INVD3BWP30P140LVT U5 ( .I(n534), .ZN(n533) );
  INVD1BWP30P140LVT U6 ( .I(i_en), .ZN(n534) );
  INVD1BWP30P140LVT U7 ( .I(rst), .ZN(n531) );
  INVD6BWP30P140LVT U8 ( .I(n531), .ZN(n532) );
  BUFFD6BWP30P140LVT U9 ( .I(n785), .Z(o_data_bus[277]) );
  BUFFD6BWP30P140LVT U10 ( .I(n786), .Z(o_data_bus[276]) );
  BUFFD6BWP30P140LVT U11 ( .I(n784), .Z(o_data_bus[278]) );
  BUFFD6BWP30P140LVT U12 ( .I(n783), .Z(o_data_bus[279]) );
  BUFFD6BWP30P140LVT U13 ( .I(n782), .Z(o_data_bus[280]) );
  BUFFD6BWP30P140LVT U14 ( .I(n781), .Z(o_data_bus[281]) );
  BUFFD6BWP30P140LVT U15 ( .I(n780), .Z(o_data_bus[282]) );
  BUFFD6BWP30P140LVT U16 ( .I(n822), .Z(o_data_bus[240]) );
  BUFFD6BWP30P140LVT U17 ( .I(n778), .Z(o_data_bus[284]) );
  BUFFD6BWP30P140LVT U18 ( .I(n777), .Z(o_data_bus[285]) );
  BUFFD6BWP30P140LVT U19 ( .I(n776), .Z(o_data_bus[286]) );
  BUFFD6BWP30P140LVT U20 ( .I(n775), .Z(o_data_bus[287]) );
  BUFFD6BWP30P140LVT U21 ( .I(n779), .Z(o_data_bus[283]) );
  BUFFD6BWP30P140LVT U22 ( .I(n773), .Z(o_data_bus[289]) );
  BUFFD6BWP30P140LVT U23 ( .I(n772), .Z(o_data_bus[290]) );
  BUFFD6BWP30P140LVT U24 ( .I(n771), .Z(o_data_bus[291]) );
  BUFFD6BWP30P140LVT U25 ( .I(n770), .Z(o_data_bus[292]) );
  BUFFD6BWP30P140LVT U26 ( .I(n774), .Z(o_data_bus[288]) );
  BUFFD6BWP30P140LVT U27 ( .I(n768), .Z(o_data_bus[294]) );
  BUFFD6BWP30P140LVT U28 ( .I(n787), .Z(o_data_bus[275]) );
  BUFFD6BWP30P140LVT U29 ( .I(n788), .Z(o_data_bus[274]) );
  BUFFD6BWP30P140LVT U30 ( .I(n789), .Z(o_data_bus[273]) );
  BUFFD6BWP30P140LVT U31 ( .I(n790), .Z(o_data_bus[272]) );
  BUFFD6BWP30P140LVT U32 ( .I(n791), .Z(o_data_bus[271]) );
  BUFFD6BWP30P140LVT U33 ( .I(n792), .Z(o_data_bus[270]) );
  BUFFD6BWP30P140LVT U34 ( .I(n793), .Z(o_data_bus[269]) );
  BUFFD6BWP30P140LVT U35 ( .I(n794), .Z(o_data_bus[268]) );
  BUFFD6BWP30P140LVT U36 ( .I(n795), .Z(o_data_bus[267]) );
  BUFFD6BWP30P140LVT U37 ( .I(n796), .Z(o_data_bus[266]) );
  BUFFD6BWP30P140LVT U38 ( .I(n797), .Z(o_data_bus[265]) );
  BUFFD6BWP30P140LVT U39 ( .I(n767), .Z(o_data_bus[295]) );
  BUFFD6BWP30P140LVT U40 ( .I(n766), .Z(o_data_bus[296]) );
  BUFFD6BWP30P140LVT U41 ( .I(n798), .Z(o_data_bus[264]) );
  BUFFD6BWP30P140LVT U42 ( .I(n799), .Z(o_data_bus[263]) );
  BUFFD6BWP30P140LVT U43 ( .I(n765), .Z(o_data_bus[297]) );
  BUFFD6BWP30P140LVT U44 ( .I(n800), .Z(o_data_bus[262]) );
  BUFFD6BWP30P140LVT U45 ( .I(n801), .Z(o_data_bus[261]) );
  BUFFD6BWP30P140LVT U46 ( .I(n802), .Z(o_data_bus[260]) );
  BUFFD6BWP30P140LVT U47 ( .I(n803), .Z(o_data_bus[259]) );
  BUFFD6BWP30P140LVT U48 ( .I(n804), .Z(o_data_bus[258]) );
  BUFFD6BWP30P140LVT U49 ( .I(n805), .Z(o_data_bus[257]) );
  BUFFD6BWP30P140LVT U50 ( .I(n806), .Z(o_data_bus[256]) );
  BUFFD6BWP30P140LVT U51 ( .I(n764), .Z(o_data_bus[298]) );
  BUFFD6BWP30P140LVT U52 ( .I(n807), .Z(o_data_bus[255]) );
  BUFFD6BWP30P140LVT U53 ( .I(n763), .Z(o_data_bus[299]) );
  BUFFD6BWP30P140LVT U54 ( .I(n808), .Z(o_data_bus[254]) );
  BUFFD6BWP30P140LVT U55 ( .I(n809), .Z(o_data_bus[253]) );
  BUFFD6BWP30P140LVT U56 ( .I(n769), .Z(o_data_bus[293]) );
  BUFFD6BWP30P140LVT U57 ( .I(n810), .Z(o_data_bus[252]) );
  BUFFD6BWP30P140LVT U58 ( .I(n811), .Z(o_data_bus[251]) );
  BUFFD6BWP30P140LVT U59 ( .I(n812), .Z(o_data_bus[250]) );
  BUFFD6BWP30P140LVT U60 ( .I(n813), .Z(o_data_bus[249]) );
  BUFFD6BWP30P140LVT U61 ( .I(n814), .Z(o_data_bus[248]) );
  BUFFD6BWP30P140LVT U62 ( .I(n815), .Z(o_data_bus[247]) );
  BUFFD6BWP30P140LVT U63 ( .I(n816), .Z(o_data_bus[246]) );
  BUFFD6BWP30P140LVT U64 ( .I(n817), .Z(o_data_bus[245]) );
  BUFFD6BWP30P140LVT U65 ( .I(n818), .Z(o_data_bus[244]) );
  BUFFD6BWP30P140LVT U66 ( .I(n819), .Z(o_data_bus[243]) );
  BUFFD6BWP30P140LVT U67 ( .I(n820), .Z(o_data_bus[242]) );
  BUFFD6BWP30P140LVT U68 ( .I(n821), .Z(o_data_bus[241]) );
  BUFFD6BWP30P140LVT U69 ( .I(n1013), .Z(o_data_bus[49]) );
  BUFFD6BWP30P140LVT U70 ( .I(n762), .Z(o_data_bus[300]) );
  BUFFD6BWP30P140LVT U71 ( .I(n823), .Z(o_data_bus[239]) );
  BUFFD6BWP30P140LVT U72 ( .I(n824), .Z(o_data_bus[238]) );
  BUFFD6BWP30P140LVT U73 ( .I(n825), .Z(o_data_bus[237]) );
  BUFFD6BWP30P140LVT U74 ( .I(n826), .Z(o_data_bus[236]) );
  BUFFD6BWP30P140LVT U75 ( .I(n827), .Z(o_data_bus[235]) );
  BUFFD6BWP30P140LVT U76 ( .I(n828), .Z(o_data_bus[234]) );
  BUFFD6BWP30P140LVT U77 ( .I(n829), .Z(o_data_bus[233]) );
  BUFFD6BWP30P140LVT U78 ( .I(n830), .Z(o_data_bus[232]) );
  BUFFD6BWP30P140LVT U79 ( .I(n831), .Z(o_data_bus[231]) );
  BUFFD6BWP30P140LVT U80 ( .I(n832), .Z(o_data_bus[230]) );
  BUFFD6BWP30P140LVT U81 ( .I(n833), .Z(o_data_bus[229]) );
  BUFFD6BWP30P140LVT U82 ( .I(n834), .Z(o_data_bus[228]) );
  BUFFD6BWP30P140LVT U83 ( .I(n835), .Z(o_data_bus[227]) );
  BUFFD6BWP30P140LVT U84 ( .I(n836), .Z(o_data_bus[226]) );
  BUFFD6BWP30P140LVT U85 ( .I(n837), .Z(o_data_bus[225]) );
  BUFFD6BWP30P140LVT U86 ( .I(n838), .Z(o_data_bus[224]) );
  BUFFD6BWP30P140LVT U87 ( .I(n839), .Z(o_data_bus[223]) );
  BUFFD6BWP30P140LVT U88 ( .I(n840), .Z(o_data_bus[222]) );
  BUFFD6BWP30P140LVT U89 ( .I(n841), .Z(o_data_bus[221]) );
  BUFFD6BWP30P140LVT U90 ( .I(n842), .Z(o_data_bus[220]) );
  BUFFD6BWP30P140LVT U91 ( .I(n843), .Z(o_data_bus[219]) );
  BUFFD6BWP30P140LVT U92 ( .I(n844), .Z(o_data_bus[218]) );
  BUFFD6BWP30P140LVT U93 ( .I(n845), .Z(o_data_bus[217]) );
  BUFFD6BWP30P140LVT U94 ( .I(n846), .Z(o_data_bus[216]) );
  BUFFD6BWP30P140LVT U95 ( .I(n847), .Z(o_data_bus[215]) );
  BUFFD6BWP30P140LVT U96 ( .I(n848), .Z(o_data_bus[214]) );
  BUFFD6BWP30P140LVT U97 ( .I(n849), .Z(o_data_bus[213]) );
  BUFFD6BWP30P140LVT U98 ( .I(n850), .Z(o_data_bus[212]) );
  BUFFD6BWP30P140LVT U99 ( .I(n851), .Z(o_data_bus[211]) );
  BUFFD6BWP30P140LVT U100 ( .I(n852), .Z(o_data_bus[210]) );
  BUFFD6BWP30P140LVT U101 ( .I(n853), .Z(o_data_bus[209]) );
  BUFFD6BWP30P140LVT U102 ( .I(n854), .Z(o_data_bus[208]) );
  BUFFD6BWP30P140LVT U103 ( .I(n855), .Z(o_data_bus[207]) );
  BUFFD6BWP30P140LVT U104 ( .I(n856), .Z(o_data_bus[206]) );
  BUFFD6BWP30P140LVT U105 ( .I(n857), .Z(o_data_bus[205]) );
  BUFFD6BWP30P140LVT U106 ( .I(n858), .Z(o_data_bus[204]) );
  BUFFD6BWP30P140LVT U107 ( .I(n859), .Z(o_data_bus[203]) );
  BUFFD6BWP30P140LVT U108 ( .I(n860), .Z(o_data_bus[202]) );
  BUFFD6BWP30P140LVT U109 ( .I(n861), .Z(o_data_bus[201]) );
  BUFFD6BWP30P140LVT U110 ( .I(n862), .Z(o_data_bus[200]) );
  BUFFD6BWP30P140LVT U111 ( .I(n863), .Z(o_data_bus[199]) );
  BUFFD6BWP30P140LVT U112 ( .I(n864), .Z(o_data_bus[198]) );
  BUFFD6BWP30P140LVT U113 ( .I(n865), .Z(o_data_bus[197]) );
  BUFFD6BWP30P140LVT U114 ( .I(n866), .Z(o_data_bus[196]) );
  BUFFD6BWP30P140LVT U115 ( .I(n867), .Z(o_data_bus[195]) );
  BUFFD6BWP30P140LVT U116 ( .I(n868), .Z(o_data_bus[194]) );
  BUFFD6BWP30P140LVT U117 ( .I(n869), .Z(o_data_bus[193]) );
  BUFFD6BWP30P140LVT U118 ( .I(n870), .Z(o_data_bus[192]) );
  BUFFD6BWP30P140LVT U119 ( .I(n871), .Z(o_data_bus[191]) );
  BUFFD6BWP30P140LVT U120 ( .I(n872), .Z(o_data_bus[190]) );
  BUFFD6BWP30P140LVT U121 ( .I(n873), .Z(o_data_bus[189]) );
  BUFFD6BWP30P140LVT U122 ( .I(n874), .Z(o_data_bus[188]) );
  BUFFD6BWP30P140LVT U123 ( .I(n875), .Z(o_data_bus[187]) );
  BUFFD6BWP30P140LVT U124 ( .I(n876), .Z(o_data_bus[186]) );
  BUFFD6BWP30P140LVT U125 ( .I(n877), .Z(o_data_bus[185]) );
  BUFFD6BWP30P140LVT U126 ( .I(n878), .Z(o_data_bus[184]) );
  BUFFD6BWP30P140LVT U127 ( .I(n879), .Z(o_data_bus[183]) );
  BUFFD6BWP30P140LVT U128 ( .I(n880), .Z(o_data_bus[182]) );
  BUFFD6BWP30P140LVT U129 ( .I(n881), .Z(o_data_bus[181]) );
  BUFFD6BWP30P140LVT U130 ( .I(n882), .Z(o_data_bus[180]) );
  BUFFD6BWP30P140LVT U131 ( .I(n883), .Z(o_data_bus[179]) );
  BUFFD6BWP30P140LVT U132 ( .I(n884), .Z(o_data_bus[178]) );
  BUFFD6BWP30P140LVT U133 ( .I(n885), .Z(o_data_bus[177]) );
  BUFFD6BWP30P140LVT U134 ( .I(n761), .Z(o_data_bus[301]) );
  BUFFD6BWP30P140LVT U135 ( .I(n715), .Z(o_data_bus[347]) );
  BUFFD6BWP30P140LVT U136 ( .I(n714), .Z(o_data_bus[348]) );
  BUFFD6BWP30P140LVT U137 ( .I(n713), .Z(o_data_bus[349]) );
  BUFFD6BWP30P140LVT U138 ( .I(n712), .Z(o_data_bus[350]) );
  BUFFD6BWP30P140LVT U139 ( .I(n711), .Z(o_data_bus[351]) );
  BUFFD6BWP30P140LVT U140 ( .I(n710), .Z(o_data_bus[352]) );
  BUFFD6BWP30P140LVT U141 ( .I(n709), .Z(o_data_bus[353]) );
  BUFFD6BWP30P140LVT U142 ( .I(n708), .Z(o_data_bus[354]) );
  BUFFD6BWP30P140LVT U143 ( .I(n707), .Z(o_data_bus[355]) );
  BUFFD6BWP30P140LVT U144 ( .I(n706), .Z(o_data_bus[356]) );
  BUFFD6BWP30P140LVT U145 ( .I(n705), .Z(o_data_bus[357]) );
  BUFFD6BWP30P140LVT U146 ( .I(n704), .Z(o_data_bus[358]) );
  BUFFD6BWP30P140LVT U147 ( .I(n703), .Z(o_data_bus[359]) );
  BUFFD6BWP30P140LVT U148 ( .I(n702), .Z(o_data_bus[360]) );
  BUFFD6BWP30P140LVT U149 ( .I(n701), .Z(o_data_bus[361]) );
  BUFFD6BWP30P140LVT U150 ( .I(n700), .Z(o_data_bus[362]) );
  BUFFD6BWP30P140LVT U151 ( .I(n699), .Z(o_data_bus[363]) );
  BUFFD6BWP30P140LVT U152 ( .I(n698), .Z(o_data_bus[364]) );
  BUFFD6BWP30P140LVT U153 ( .I(n697), .Z(o_data_bus[365]) );
  BUFFD6BWP30P140LVT U154 ( .I(n696), .Z(o_data_bus[366]) );
  BUFFD6BWP30P140LVT U155 ( .I(n695), .Z(o_data_bus[367]) );
  BUFFD6BWP30P140LVT U156 ( .I(n694), .Z(o_data_bus[368]) );
  BUFFD6BWP30P140LVT U157 ( .I(n693), .Z(o_data_bus[369]) );
  BUFFD6BWP30P140LVT U158 ( .I(n692), .Z(o_data_bus[370]) );
  BUFFD6BWP30P140LVT U159 ( .I(n691), .Z(o_data_bus[371]) );
  BUFFD6BWP30P140LVT U160 ( .I(n690), .Z(o_data_bus[372]) );
  BUFFD6BWP30P140LVT U161 ( .I(n689), .Z(o_data_bus[373]) );
  BUFFD6BWP30P140LVT U162 ( .I(n688), .Z(o_data_bus[374]) );
  BUFFD6BWP30P140LVT U163 ( .I(n687), .Z(o_data_bus[375]) );
  BUFFD6BWP30P140LVT U164 ( .I(n686), .Z(o_data_bus[376]) );
  BUFFD6BWP30P140LVT U165 ( .I(n718), .Z(o_data_bus[344]) );
  BUFFD6BWP30P140LVT U166 ( .I(n685), .Z(o_data_bus[377]) );
  BUFFD6BWP30P140LVT U167 ( .I(n719), .Z(o_data_bus[343]) );
  BUFFD6BWP30P140LVT U168 ( .I(n720), .Z(o_data_bus[342]) );
  BUFFD6BWP30P140LVT U169 ( .I(n684), .Z(o_data_bus[378]) );
  BUFFD6BWP30P140LVT U170 ( .I(n683), .Z(o_data_bus[379]) );
  BUFFD6BWP30P140LVT U171 ( .I(n721), .Z(o_data_bus[341]) );
  BUFFD6BWP30P140LVT U172 ( .I(n722), .Z(o_data_bus[340]) );
  BUFFD6BWP30P140LVT U173 ( .I(n682), .Z(o_data_bus[380]) );
  BUFFD6BWP30P140LVT U174 ( .I(n681), .Z(o_data_bus[381]) );
  BUFFD6BWP30P140LVT U175 ( .I(n680), .Z(o_data_bus[382]) );
  BUFFD6BWP30P140LVT U176 ( .I(n723), .Z(o_data_bus[339]) );
  BUFFD6BWP30P140LVT U177 ( .I(n724), .Z(o_data_bus[338]) );
  BUFFD6BWP30P140LVT U178 ( .I(n679), .Z(o_data_bus[383]) );
  BUFFD6BWP30P140LVT U179 ( .I(n678), .Z(o_data_bus[384]) );
  BUFFD6BWP30P140LVT U180 ( .I(n725), .Z(o_data_bus[337]) );
  BUFFD6BWP30P140LVT U181 ( .I(n726), .Z(o_data_bus[336]) );
  BUFFD6BWP30P140LVT U182 ( .I(n677), .Z(o_data_bus[385]) );
  BUFFD6BWP30P140LVT U183 ( .I(n676), .Z(o_data_bus[386]) );
  BUFFD6BWP30P140LVT U184 ( .I(n727), .Z(o_data_bus[335]) );
  BUFFD6BWP30P140LVT U185 ( .I(n728), .Z(o_data_bus[334]) );
  BUFFD6BWP30P140LVT U186 ( .I(n675), .Z(o_data_bus[387]) );
  BUFFD6BWP30P140LVT U187 ( .I(n674), .Z(o_data_bus[388]) );
  BUFFD6BWP30P140LVT U188 ( .I(n729), .Z(o_data_bus[333]) );
  BUFFD6BWP30P140LVT U189 ( .I(n730), .Z(o_data_bus[332]) );
  BUFFD6BWP30P140LVT U190 ( .I(n673), .Z(o_data_bus[389]) );
  BUFFD6BWP30P140LVT U191 ( .I(n672), .Z(o_data_bus[390]) );
  BUFFD6BWP30P140LVT U192 ( .I(n731), .Z(o_data_bus[331]) );
  BUFFD6BWP30P140LVT U193 ( .I(n732), .Z(o_data_bus[330]) );
  BUFFD6BWP30P140LVT U194 ( .I(n671), .Z(o_data_bus[391]) );
  BUFFD6BWP30P140LVT U195 ( .I(n670), .Z(o_data_bus[392]) );
  BUFFD6BWP30P140LVT U196 ( .I(n733), .Z(o_data_bus[329]) );
  BUFFD6BWP30P140LVT U197 ( .I(n734), .Z(o_data_bus[328]) );
  BUFFD6BWP30P140LVT U198 ( .I(n669), .Z(o_data_bus[393]) );
  BUFFD6BWP30P140LVT U199 ( .I(n668), .Z(o_data_bus[394]) );
  BUFFD6BWP30P140LVT U200 ( .I(n735), .Z(o_data_bus[327]) );
  BUFFD6BWP30P140LVT U201 ( .I(n736), .Z(o_data_bus[326]) );
  BUFFD6BWP30P140LVT U202 ( .I(n667), .Z(o_data_bus[395]) );
  BUFFD6BWP30P140LVT U203 ( .I(n666), .Z(o_data_bus[396]) );
  BUFFD6BWP30P140LVT U204 ( .I(n737), .Z(o_data_bus[325]) );
  BUFFD6BWP30P140LVT U205 ( .I(n738), .Z(o_data_bus[324]) );
  BUFFD6BWP30P140LVT U206 ( .I(n665), .Z(o_data_bus[397]) );
  BUFFD6BWP30P140LVT U207 ( .I(n664), .Z(o_data_bus[398]) );
  BUFFD6BWP30P140LVT U208 ( .I(n663), .Z(o_data_bus[399]) );
  BUFFD6BWP30P140LVT U209 ( .I(n662), .Z(o_data_bus[400]) );
  BUFFD6BWP30P140LVT U210 ( .I(n661), .Z(o_data_bus[401]) );
  BUFFD6BWP30P140LVT U211 ( .I(n660), .Z(o_data_bus[402]) );
  BUFFD6BWP30P140LVT U212 ( .I(n886), .Z(o_data_bus[176]) );
  BUFFD6BWP30P140LVT U213 ( .I(n658), .Z(o_data_bus[404]) );
  BUFFD6BWP30P140LVT U214 ( .I(n657), .Z(o_data_bus[405]) );
  BUFFD6BWP30P140LVT U215 ( .I(n716), .Z(o_data_bus[346]) );
  BUFFD6BWP30P140LVT U216 ( .I(n656), .Z(o_data_bus[406]) );
  BUFFD6BWP30P140LVT U217 ( .I(n655), .Z(o_data_bus[407]) );
  BUFFD6BWP30P140LVT U218 ( .I(n654), .Z(o_data_bus[408]) );
  BUFFD6BWP30P140LVT U219 ( .I(n739), .Z(o_data_bus[323]) );
  BUFFD6BWP30P140LVT U220 ( .I(n653), .Z(o_data_bus[409]) );
  BUFFD6BWP30P140LVT U221 ( .I(n652), .Z(o_data_bus[410]) );
  BUFFD6BWP30P140LVT U222 ( .I(n651), .Z(o_data_bus[411]) );
  BUFFD6BWP30P140LVT U223 ( .I(n650), .Z(o_data_bus[412]) );
  BUFFD6BWP30P140LVT U224 ( .I(n649), .Z(o_data_bus[413]) );
  BUFFD6BWP30P140LVT U225 ( .I(n648), .Z(o_data_bus[414]) );
  BUFFD6BWP30P140LVT U226 ( .I(n647), .Z(o_data_bus[415]) );
  BUFFD6BWP30P140LVT U227 ( .I(n646), .Z(o_data_bus[416]) );
  BUFFD6BWP30P140LVT U228 ( .I(n645), .Z(o_data_bus[417]) );
  BUFFD6BWP30P140LVT U229 ( .I(n644), .Z(o_data_bus[418]) );
  BUFFD6BWP30P140LVT U230 ( .I(n643), .Z(o_data_bus[419]) );
  BUFFD6BWP30P140LVT U231 ( .I(n642), .Z(o_data_bus[420]) );
  BUFFD6BWP30P140LVT U232 ( .I(n641), .Z(o_data_bus[421]) );
  BUFFD6BWP30P140LVT U233 ( .I(n640), .Z(o_data_bus[422]) );
  BUFFD6BWP30P140LVT U234 ( .I(n639), .Z(o_data_bus[423]) );
  BUFFD6BWP30P140LVT U235 ( .I(n638), .Z(o_data_bus[424]) );
  BUFFD6BWP30P140LVT U236 ( .I(n637), .Z(o_data_bus[425]) );
  BUFFD6BWP30P140LVT U237 ( .I(n636), .Z(o_data_bus[426]) );
  BUFFD6BWP30P140LVT U238 ( .I(n635), .Z(o_data_bus[427]) );
  BUFFD6BWP30P140LVT U239 ( .I(n634), .Z(o_data_bus[428]) );
  BUFFD6BWP30P140LVT U240 ( .I(n633), .Z(o_data_bus[429]) );
  BUFFD6BWP30P140LVT U241 ( .I(n632), .Z(o_data_bus[430]) );
  BUFFD6BWP30P140LVT U242 ( .I(n631), .Z(o_data_bus[431]) );
  BUFFD6BWP30P140LVT U243 ( .I(n630), .Z(o_data_bus[432]) );
  BUFFD6BWP30P140LVT U244 ( .I(n629), .Z(o_data_bus[433]) );
  BUFFD6BWP30P140LVT U245 ( .I(n628), .Z(o_data_bus[434]) );
  BUFFD6BWP30P140LVT U246 ( .I(n627), .Z(o_data_bus[435]) );
  BUFFD6BWP30P140LVT U247 ( .I(n626), .Z(o_data_bus[436]) );
  BUFFD6BWP30P140LVT U248 ( .I(n625), .Z(o_data_bus[437]) );
  BUFFD6BWP30P140LVT U249 ( .I(n624), .Z(o_data_bus[438]) );
  BUFFD6BWP30P140LVT U250 ( .I(n623), .Z(o_data_bus[439]) );
  BUFFD6BWP30P140LVT U251 ( .I(n622), .Z(o_data_bus[440]) );
  BUFFD6BWP30P140LVT U252 ( .I(n740), .Z(o_data_bus[322]) );
  BUFFD6BWP30P140LVT U253 ( .I(n621), .Z(o_data_bus[441]) );
  BUFFD6BWP30P140LVT U254 ( .I(n620), .Z(o_data_bus[442]) );
  BUFFD6BWP30P140LVT U255 ( .I(n619), .Z(o_data_bus[443]) );
  BUFFD6BWP30P140LVT U256 ( .I(n618), .Z(o_data_bus[444]) );
  BUFFD6BWP30P140LVT U257 ( .I(n617), .Z(o_data_bus[445]) );
  BUFFD6BWP30P140LVT U258 ( .I(n616), .Z(o_data_bus[446]) );
  BUFFD6BWP30P140LVT U259 ( .I(n615), .Z(o_data_bus[447]) );
  BUFFD6BWP30P140LVT U260 ( .I(n614), .Z(o_data_bus[448]) );
  BUFFD6BWP30P140LVT U261 ( .I(n613), .Z(o_data_bus[449]) );
  BUFFD6BWP30P140LVT U262 ( .I(n612), .Z(o_data_bus[450]) );
  BUFFD6BWP30P140LVT U263 ( .I(n611), .Z(o_data_bus[451]) );
  BUFFD6BWP30P140LVT U264 ( .I(n610), .Z(o_data_bus[452]) );
  BUFFD6BWP30P140LVT U265 ( .I(n609), .Z(o_data_bus[453]) );
  BUFFD6BWP30P140LVT U266 ( .I(n608), .Z(o_data_bus[454]) );
  BUFFD6BWP30P140LVT U267 ( .I(n607), .Z(o_data_bus[455]) );
  BUFFD6BWP30P140LVT U268 ( .I(n606), .Z(o_data_bus[456]) );
  BUFFD6BWP30P140LVT U269 ( .I(n605), .Z(o_data_bus[457]) );
  BUFFD6BWP30P140LVT U270 ( .I(n604), .Z(o_data_bus[458]) );
  BUFFD6BWP30P140LVT U271 ( .I(n603), .Z(o_data_bus[459]) );
  BUFFD6BWP30P140LVT U272 ( .I(n602), .Z(o_data_bus[460]) );
  BUFFD6BWP30P140LVT U273 ( .I(n601), .Z(o_data_bus[461]) );
  BUFFD6BWP30P140LVT U274 ( .I(n600), .Z(o_data_bus[462]) );
  BUFFD6BWP30P140LVT U275 ( .I(n741), .Z(o_data_bus[321]) );
  BUFFD6BWP30P140LVT U276 ( .I(n742), .Z(o_data_bus[320]) );
  BUFFD6BWP30P140LVT U277 ( .I(n743), .Z(o_data_bus[319]) );
  BUFFD6BWP30P140LVT U278 ( .I(n744), .Z(o_data_bus[318]) );
  BUFFD6BWP30P140LVT U279 ( .I(n745), .Z(o_data_bus[317]) );
  BUFFD6BWP30P140LVT U280 ( .I(n746), .Z(o_data_bus[316]) );
  BUFFD6BWP30P140LVT U281 ( .I(n747), .Z(o_data_bus[315]) );
  BUFFD6BWP30P140LVT U282 ( .I(n748), .Z(o_data_bus[314]) );
  BUFFD6BWP30P140LVT U283 ( .I(n749), .Z(o_data_bus[313]) );
  BUFFD6BWP30P140LVT U284 ( .I(n750), .Z(o_data_bus[312]) );
  BUFFD6BWP30P140LVT U285 ( .I(n751), .Z(o_data_bus[311]) );
  BUFFD6BWP30P140LVT U286 ( .I(n752), .Z(o_data_bus[310]) );
  BUFFD6BWP30P140LVT U287 ( .I(n753), .Z(o_data_bus[309]) );
  BUFFD6BWP30P140LVT U288 ( .I(n754), .Z(o_data_bus[308]) );
  BUFFD6BWP30P140LVT U289 ( .I(n755), .Z(o_data_bus[307]) );
  BUFFD6BWP30P140LVT U290 ( .I(n756), .Z(o_data_bus[306]) );
  BUFFD6BWP30P140LVT U291 ( .I(n757), .Z(o_data_bus[305]) );
  BUFFD6BWP30P140LVT U292 ( .I(n758), .Z(o_data_bus[304]) );
  BUFFD6BWP30P140LVT U293 ( .I(n759), .Z(o_data_bus[303]) );
  BUFFD6BWP30P140LVT U294 ( .I(n760), .Z(o_data_bus[302]) );
  BUFFD6BWP30P140LVT U295 ( .I(n659), .Z(o_data_bus[403]) );
  BUFFD6BWP30P140LVT U296 ( .I(n887), .Z(o_data_bus[175]) );
  BUFFD6BWP30P140LVT U297 ( .I(n961), .Z(o_data_bus[101]) );
  BUFFD6BWP30P140LVT U298 ( .I(n962), .Z(o_data_bus[100]) );
  BUFFD6BWP30P140LVT U299 ( .I(n963), .Z(o_data_bus[99]) );
  BUFFD6BWP30P140LVT U300 ( .I(n964), .Z(o_data_bus[98]) );
  BUFFD6BWP30P140LVT U301 ( .I(n965), .Z(o_data_bus[97]) );
  BUFFD6BWP30P140LVT U302 ( .I(n966), .Z(o_data_bus[96]) );
  BUFFD6BWP30P140LVT U303 ( .I(n967), .Z(o_data_bus[95]) );
  BUFFD6BWP30P140LVT U304 ( .I(n968), .Z(o_data_bus[94]) );
  BUFFD6BWP30P140LVT U305 ( .I(n969), .Z(o_data_bus[93]) );
  BUFFD6BWP30P140LVT U306 ( .I(n970), .Z(o_data_bus[92]) );
  BUFFD6BWP30P140LVT U307 ( .I(n971), .Z(o_data_bus[91]) );
  BUFFD6BWP30P140LVT U308 ( .I(n972), .Z(o_data_bus[90]) );
  BUFFD6BWP30P140LVT U309 ( .I(n973), .Z(o_data_bus[89]) );
  BUFFD6BWP30P140LVT U310 ( .I(n974), .Z(o_data_bus[88]) );
  BUFFD6BWP30P140LVT U311 ( .I(n975), .Z(o_data_bus[87]) );
  BUFFD6BWP30P140LVT U312 ( .I(n976), .Z(o_data_bus[86]) );
  BUFFD6BWP30P140LVT U313 ( .I(n977), .Z(o_data_bus[85]) );
  BUFFD6BWP30P140LVT U314 ( .I(n978), .Z(o_data_bus[84]) );
  BUFFD6BWP30P140LVT U315 ( .I(n979), .Z(o_data_bus[83]) );
  BUFFD6BWP30P140LVT U316 ( .I(n980), .Z(o_data_bus[82]) );
  BUFFD6BWP30P140LVT U317 ( .I(n981), .Z(o_data_bus[81]) );
  BUFFD6BWP30P140LVT U318 ( .I(n982), .Z(o_data_bus[80]) );
  BUFFD6BWP30P140LVT U319 ( .I(n983), .Z(o_data_bus[79]) );
  BUFFD6BWP30P140LVT U320 ( .I(n536), .Z(o_valid[14]) );
  BUFFD6BWP30P140LVT U321 ( .I(n569), .Z(o_data_bus[493]) );
  BUFFD6BWP30P140LVT U322 ( .I(n568), .Z(o_data_bus[494]) );
  BUFFD6BWP30P140LVT U323 ( .I(n567), .Z(o_data_bus[495]) );
  BUFFD6BWP30P140LVT U324 ( .I(n566), .Z(o_data_bus[496]) );
  BUFFD6BWP30P140LVT U325 ( .I(n565), .Z(o_data_bus[497]) );
  BUFFD6BWP30P140LVT U326 ( .I(n564), .Z(o_data_bus[498]) );
  BUFFD6BWP30P140LVT U327 ( .I(n984), .Z(o_data_bus[78]) );
  BUFFD6BWP30P140LVT U328 ( .I(n985), .Z(o_data_bus[77]) );
  BUFFD6BWP30P140LVT U329 ( .I(n986), .Z(o_data_bus[76]) );
  BUFFD6BWP30P140LVT U330 ( .I(n563), .Z(o_data_bus[499]) );
  BUFFD6BWP30P140LVT U331 ( .I(n562), .Z(o_data_bus[500]) );
  BUFFD6BWP30P140LVT U332 ( .I(n561), .Z(o_data_bus[501]) );
  BUFFD6BWP30P140LVT U333 ( .I(n560), .Z(o_data_bus[502]) );
  BUFFD6BWP30P140LVT U334 ( .I(n559), .Z(o_data_bus[503]) );
  BUFFD6BWP30P140LVT U335 ( .I(n558), .Z(o_data_bus[504]) );
  BUFFD6BWP30P140LVT U336 ( .I(n557), .Z(o_data_bus[505]) );
  BUFFD6BWP30P140LVT U337 ( .I(n556), .Z(o_data_bus[506]) );
  BUFFD6BWP30P140LVT U338 ( .I(n555), .Z(o_data_bus[507]) );
  BUFFD6BWP30P140LVT U339 ( .I(n554), .Z(o_data_bus[508]) );
  BUFFD6BWP30P140LVT U340 ( .I(n553), .Z(o_data_bus[509]) );
  BUFFD6BWP30P140LVT U341 ( .I(n552), .Z(o_data_bus[510]) );
  BUFFD6BWP30P140LVT U342 ( .I(n551), .Z(o_data_bus[511]) );
  BUFFD6BWP30P140LVT U343 ( .I(n550), .Z(o_valid[0]) );
  BUFFD6BWP30P140LVT U344 ( .I(n549), .Z(o_valid[1]) );
  BUFFD6BWP30P140LVT U345 ( .I(n548), .Z(o_valid[2]) );
  BUFFD6BWP30P140LVT U346 ( .I(n547), .Z(o_valid[3]) );
  BUFFD6BWP30P140LVT U347 ( .I(n987), .Z(o_data_bus[75]) );
  BUFFD6BWP30P140LVT U348 ( .I(n988), .Z(o_data_bus[74]) );
  BUFFD6BWP30P140LVT U349 ( .I(n989), .Z(o_data_bus[73]) );
  BUFFD6BWP30P140LVT U350 ( .I(n990), .Z(o_data_bus[72]) );
  BUFFD6BWP30P140LVT U351 ( .I(n991), .Z(o_data_bus[71]) );
  BUFFD6BWP30P140LVT U352 ( .I(n992), .Z(o_data_bus[70]) );
  BUFFD6BWP30P140LVT U353 ( .I(n993), .Z(o_data_bus[69]) );
  BUFFD6BWP30P140LVT U354 ( .I(n994), .Z(o_data_bus[68]) );
  BUFFD6BWP30P140LVT U355 ( .I(n995), .Z(o_data_bus[67]) );
  BUFFD6BWP30P140LVT U356 ( .I(n996), .Z(o_data_bus[66]) );
  BUFFD6BWP30P140LVT U357 ( .I(n997), .Z(o_data_bus[65]) );
  BUFFD6BWP30P140LVT U358 ( .I(n546), .Z(o_valid[4]) );
  BUFFD6BWP30P140LVT U359 ( .I(n545), .Z(o_valid[5]) );
  BUFFD6BWP30P140LVT U360 ( .I(n544), .Z(o_valid[6]) );
  BUFFD6BWP30P140LVT U361 ( .I(n543), .Z(o_valid[7]) );
  BUFFD6BWP30P140LVT U362 ( .I(n542), .Z(o_valid[8]) );
  BUFFD6BWP30P140LVT U363 ( .I(n541), .Z(o_valid[9]) );
  BUFFD6BWP30P140LVT U364 ( .I(n960), .Z(o_data_bus[102]) );
  BUFFD6BWP30P140LVT U365 ( .I(n998), .Z(o_data_bus[64]) );
  BUFFD6BWP30P140LVT U366 ( .I(n999), .Z(o_data_bus[63]) );
  BUFFD6BWP30P140LVT U367 ( .I(n1000), .Z(o_data_bus[62]) );
  BUFFD6BWP30P140LVT U368 ( .I(n1001), .Z(o_data_bus[61]) );
  BUFFD6BWP30P140LVT U369 ( .I(n1002), .Z(o_data_bus[60]) );
  BUFFD6BWP30P140LVT U370 ( .I(n1003), .Z(o_data_bus[59]) );
  BUFFD6BWP30P140LVT U371 ( .I(n1004), .Z(o_data_bus[58]) );
  BUFFD6BWP30P140LVT U372 ( .I(n1005), .Z(o_data_bus[57]) );
  BUFFD6BWP30P140LVT U373 ( .I(n1006), .Z(o_data_bus[56]) );
  BUFFD6BWP30P140LVT U374 ( .I(n1007), .Z(o_data_bus[55]) );
  BUFFD6BWP30P140LVT U375 ( .I(n1008), .Z(o_data_bus[54]) );
  BUFFD6BWP30P140LVT U376 ( .I(n1009), .Z(o_data_bus[53]) );
  BUFFD6BWP30P140LVT U377 ( .I(n1010), .Z(o_data_bus[52]) );
  BUFFD6BWP30P140LVT U378 ( .I(n1011), .Z(o_data_bus[51]) );
  BUFFD6BWP30P140LVT U379 ( .I(n1012), .Z(o_data_bus[50]) );
  BUFFD6BWP30P140LVT U380 ( .I(n540), .Z(o_valid[10]) );
  BUFFD6BWP30P140LVT U381 ( .I(n539), .Z(o_valid[11]) );
  BUFFD6BWP30P140LVT U382 ( .I(n1062), .Z(o_data_bus[0]) );
  BUFFD6BWP30P140LVT U383 ( .I(n1061), .Z(o_data_bus[1]) );
  BUFFD6BWP30P140LVT U384 ( .I(n1060), .Z(o_data_bus[2]) );
  BUFFD6BWP30P140LVT U385 ( .I(n1059), .Z(o_data_bus[3]) );
  BUFFD6BWP30P140LVT U386 ( .I(n1058), .Z(o_data_bus[4]) );
  BUFFD6BWP30P140LVT U387 ( .I(n1057), .Z(o_data_bus[5]) );
  BUFFD6BWP30P140LVT U388 ( .I(n1056), .Z(o_data_bus[6]) );
  BUFFD6BWP30P140LVT U389 ( .I(n1055), .Z(o_data_bus[7]) );
  BUFFD6BWP30P140LVT U390 ( .I(n1054), .Z(o_data_bus[8]) );
  BUFFD6BWP30P140LVT U391 ( .I(n1053), .Z(o_data_bus[9]) );
  BUFFD6BWP30P140LVT U392 ( .I(n1052), .Z(o_data_bus[10]) );
  BUFFD6BWP30P140LVT U393 ( .I(n1051), .Z(o_data_bus[11]) );
  BUFFD6BWP30P140LVT U394 ( .I(n1050), .Z(o_data_bus[12]) );
  BUFFD6BWP30P140LVT U395 ( .I(n1049), .Z(o_data_bus[13]) );
  BUFFD6BWP30P140LVT U396 ( .I(n1048), .Z(o_data_bus[14]) );
  BUFFD6BWP30P140LVT U397 ( .I(n538), .Z(o_valid[12]) );
  BUFFD6BWP30P140LVT U398 ( .I(n1047), .Z(o_data_bus[15]) );
  BUFFD6BWP30P140LVT U399 ( .I(n1046), .Z(o_data_bus[16]) );
  BUFFD6BWP30P140LVT U400 ( .I(n1045), .Z(o_data_bus[17]) );
  BUFFD6BWP30P140LVT U401 ( .I(n1044), .Z(o_data_bus[18]) );
  BUFFD6BWP30P140LVT U402 ( .I(n1043), .Z(o_data_bus[19]) );
  BUFFD6BWP30P140LVT U403 ( .I(n1042), .Z(o_data_bus[20]) );
  BUFFD6BWP30P140LVT U404 ( .I(n1041), .Z(o_data_bus[21]) );
  BUFFD6BWP30P140LVT U405 ( .I(n1040), .Z(o_data_bus[22]) );
  BUFFD6BWP30P140LVT U406 ( .I(n1039), .Z(o_data_bus[23]) );
  BUFFD6BWP30P140LVT U407 ( .I(n1038), .Z(o_data_bus[24]) );
  BUFFD6BWP30P140LVT U408 ( .I(n1037), .Z(o_data_bus[25]) );
  BUFFD6BWP30P140LVT U409 ( .I(n1036), .Z(o_data_bus[26]) );
  BUFFD6BWP30P140LVT U410 ( .I(n1035), .Z(o_data_bus[27]) );
  BUFFD6BWP30P140LVT U411 ( .I(n1034), .Z(o_data_bus[28]) );
  BUFFD6BWP30P140LVT U412 ( .I(n1033), .Z(o_data_bus[29]) );
  BUFFD6BWP30P140LVT U413 ( .I(n1032), .Z(o_data_bus[30]) );
  BUFFD6BWP30P140LVT U414 ( .I(n1031), .Z(o_data_bus[31]) );
  BUFFD6BWP30P140LVT U415 ( .I(n1030), .Z(o_data_bus[32]) );
  BUFFD6BWP30P140LVT U416 ( .I(n1029), .Z(o_data_bus[33]) );
  BUFFD6BWP30P140LVT U417 ( .I(n1028), .Z(o_data_bus[34]) );
  BUFFD6BWP30P140LVT U418 ( .I(n1027), .Z(o_data_bus[35]) );
  BUFFD6BWP30P140LVT U419 ( .I(n1026), .Z(o_data_bus[36]) );
  BUFFD6BWP30P140LVT U420 ( .I(n1025), .Z(o_data_bus[37]) );
  BUFFD6BWP30P140LVT U421 ( .I(n1024), .Z(o_data_bus[38]) );
  BUFFD6BWP30P140LVT U422 ( .I(n1023), .Z(o_data_bus[39]) );
  BUFFD6BWP30P140LVT U423 ( .I(n1022), .Z(o_data_bus[40]) );
  BUFFD6BWP30P140LVT U424 ( .I(n1021), .Z(o_data_bus[41]) );
  BUFFD6BWP30P140LVT U425 ( .I(n1020), .Z(o_data_bus[42]) );
  BUFFD6BWP30P140LVT U426 ( .I(n1019), .Z(o_data_bus[43]) );
  BUFFD6BWP30P140LVT U427 ( .I(n1018), .Z(o_data_bus[44]) );
  BUFFD6BWP30P140LVT U428 ( .I(n1017), .Z(o_data_bus[45]) );
  BUFFD6BWP30P140LVT U429 ( .I(n1016), .Z(o_data_bus[46]) );
  BUFFD6BWP30P140LVT U430 ( .I(n537), .Z(o_valid[13]) );
  BUFFD6BWP30P140LVT U431 ( .I(n1015), .Z(o_data_bus[47]) );
  BUFFD6BWP30P140LVT U432 ( .I(n1014), .Z(o_data_bus[48]) );
  BUFFD6BWP30P140LVT U433 ( .I(n888), .Z(o_data_bus[174]) );
  BUFFD6BWP30P140LVT U434 ( .I(n889), .Z(o_data_bus[173]) );
  BUFFD6BWP30P140LVT U435 ( .I(n890), .Z(o_data_bus[172]) );
  BUFFD6BWP30P140LVT U436 ( .I(n891), .Z(o_data_bus[171]) );
  BUFFD6BWP30P140LVT U437 ( .I(n892), .Z(o_data_bus[170]) );
  BUFFD6BWP30P140LVT U438 ( .I(n893), .Z(o_data_bus[169]) );
  BUFFD6BWP30P140LVT U439 ( .I(n894), .Z(o_data_bus[168]) );
  BUFFD6BWP30P140LVT U440 ( .I(n895), .Z(o_data_bus[167]) );
  BUFFD6BWP30P140LVT U441 ( .I(n896), .Z(o_data_bus[166]) );
  BUFFD6BWP30P140LVT U442 ( .I(n897), .Z(o_data_bus[165]) );
  BUFFD6BWP30P140LVT U443 ( .I(n898), .Z(o_data_bus[164]) );
  BUFFD6BWP30P140LVT U444 ( .I(n899), .Z(o_data_bus[163]) );
  BUFFD6BWP30P140LVT U445 ( .I(n900), .Z(o_data_bus[162]) );
  BUFFD6BWP30P140LVT U446 ( .I(n901), .Z(o_data_bus[161]) );
  BUFFD6BWP30P140LVT U447 ( .I(n902), .Z(o_data_bus[160]) );
  BUFFD6BWP30P140LVT U448 ( .I(n717), .Z(o_data_bus[345]) );
  BUFFD6BWP30P140LVT U449 ( .I(n904), .Z(o_data_bus[158]) );
  BUFFD6BWP30P140LVT U450 ( .I(n905), .Z(o_data_bus[157]) );
  BUFFD6BWP30P140LVT U451 ( .I(n906), .Z(o_data_bus[156]) );
  BUFFD6BWP30P140LVT U452 ( .I(n907), .Z(o_data_bus[155]) );
  BUFFD6BWP30P140LVT U453 ( .I(n908), .Z(o_data_bus[154]) );
  BUFFD6BWP30P140LVT U454 ( .I(n909), .Z(o_data_bus[153]) );
  BUFFD6BWP30P140LVT U455 ( .I(n910), .Z(o_data_bus[152]) );
  BUFFD6BWP30P140LVT U456 ( .I(n911), .Z(o_data_bus[151]) );
  BUFFD6BWP30P140LVT U457 ( .I(n912), .Z(o_data_bus[150]) );
  BUFFD6BWP30P140LVT U458 ( .I(n913), .Z(o_data_bus[149]) );
  BUFFD6BWP30P140LVT U459 ( .I(n914), .Z(o_data_bus[148]) );
  BUFFD6BWP30P140LVT U460 ( .I(n915), .Z(o_data_bus[147]) );
  BUFFD6BWP30P140LVT U461 ( .I(n916), .Z(o_data_bus[146]) );
  BUFFD6BWP30P140LVT U462 ( .I(n917), .Z(o_data_bus[145]) );
  BUFFD6BWP30P140LVT U463 ( .I(n918), .Z(o_data_bus[144]) );
  BUFFD6BWP30P140LVT U464 ( .I(n919), .Z(o_data_bus[143]) );
  BUFFD6BWP30P140LVT U465 ( .I(n920), .Z(o_data_bus[142]) );
  BUFFD6BWP30P140LVT U466 ( .I(n921), .Z(o_data_bus[141]) );
  BUFFD6BWP30P140LVT U467 ( .I(n922), .Z(o_data_bus[140]) );
  BUFFD6BWP30P140LVT U468 ( .I(n923), .Z(o_data_bus[139]) );
  BUFFD6BWP30P140LVT U469 ( .I(n924), .Z(o_data_bus[138]) );
  BUFFD6BWP30P140LVT U470 ( .I(n925), .Z(o_data_bus[137]) );
  BUFFD6BWP30P140LVT U471 ( .I(n926), .Z(o_data_bus[136]) );
  BUFFD6BWP30P140LVT U472 ( .I(n927), .Z(o_data_bus[135]) );
  BUFFD6BWP30P140LVT U473 ( .I(n928), .Z(o_data_bus[134]) );
  BUFFD6BWP30P140LVT U474 ( .I(n599), .Z(o_data_bus[463]) );
  BUFFD6BWP30P140LVT U475 ( .I(n598), .Z(o_data_bus[464]) );
  BUFFD6BWP30P140LVT U476 ( .I(n597), .Z(o_data_bus[465]) );
  BUFFD6BWP30P140LVT U477 ( .I(n929), .Z(o_data_bus[133]) );
  BUFFD6BWP30P140LVT U478 ( .I(n930), .Z(o_data_bus[132]) );
  BUFFD6BWP30P140LVT U479 ( .I(n596), .Z(o_data_bus[466]) );
  BUFFD6BWP30P140LVT U480 ( .I(n595), .Z(o_data_bus[467]) );
  BUFFD6BWP30P140LVT U481 ( .I(n931), .Z(o_data_bus[131]) );
  BUFFD6BWP30P140LVT U482 ( .I(n932), .Z(o_data_bus[130]) );
  BUFFD6BWP30P140LVT U483 ( .I(n594), .Z(o_data_bus[468]) );
  BUFFD6BWP30P140LVT U484 ( .I(n593), .Z(o_data_bus[469]) );
  BUFFD6BWP30P140LVT U485 ( .I(n933), .Z(o_data_bus[129]) );
  BUFFD6BWP30P140LVT U486 ( .I(n934), .Z(o_data_bus[128]) );
  BUFFD6BWP30P140LVT U487 ( .I(n592), .Z(o_data_bus[470]) );
  BUFFD6BWP30P140LVT U488 ( .I(n591), .Z(o_data_bus[471]) );
  BUFFD6BWP30P140LVT U489 ( .I(n935), .Z(o_data_bus[127]) );
  BUFFD6BWP30P140LVT U490 ( .I(n936), .Z(o_data_bus[126]) );
  BUFFD6BWP30P140LVT U491 ( .I(n590), .Z(o_data_bus[472]) );
  BUFFD6BWP30P140LVT U492 ( .I(n589), .Z(o_data_bus[473]) );
  BUFFD6BWP30P140LVT U493 ( .I(n937), .Z(o_data_bus[125]) );
  BUFFD6BWP30P140LVT U494 ( .I(n938), .Z(o_data_bus[124]) );
  BUFFD6BWP30P140LVT U495 ( .I(n588), .Z(o_data_bus[474]) );
  BUFFD6BWP30P140LVT U496 ( .I(n587), .Z(o_data_bus[475]) );
  BUFFD6BWP30P140LVT U497 ( .I(n939), .Z(o_data_bus[123]) );
  BUFFD6BWP30P140LVT U498 ( .I(n586), .Z(o_data_bus[476]) );
  BUFFD6BWP30P140LVT U499 ( .I(n585), .Z(o_data_bus[477]) );
  BUFFD6BWP30P140LVT U500 ( .I(n584), .Z(o_data_bus[478]) );
  BUFFD6BWP30P140LVT U501 ( .I(n940), .Z(o_data_bus[122]) );
  BUFFD6BWP30P140LVT U502 ( .I(n941), .Z(o_data_bus[121]) );
  BUFFD6BWP30P140LVT U503 ( .I(n583), .Z(o_data_bus[479]) );
  BUFFD6BWP30P140LVT U504 ( .I(n582), .Z(o_data_bus[480]) );
  BUFFD6BWP30P140LVT U505 ( .I(n942), .Z(o_data_bus[120]) );
  BUFFD6BWP30P140LVT U506 ( .I(n943), .Z(o_data_bus[119]) );
  BUFFD6BWP30P140LVT U507 ( .I(n581), .Z(o_data_bus[481]) );
  BUFFD6BWP30P140LVT U508 ( .I(n580), .Z(o_data_bus[482]) );
  BUFFD6BWP30P140LVT U509 ( .I(n579), .Z(o_data_bus[483]) );
  BUFFD6BWP30P140LVT U510 ( .I(n944), .Z(o_data_bus[118]) );
  BUFFD6BWP30P140LVT U511 ( .I(n945), .Z(o_data_bus[117]) );
  BUFFD6BWP30P140LVT U512 ( .I(n578), .Z(o_data_bus[484]) );
  BUFFD6BWP30P140LVT U513 ( .I(n903), .Z(o_data_bus[159]) );
  BUFFD6BWP30P140LVT U514 ( .I(n577), .Z(o_data_bus[485]) );
  BUFFD6BWP30P140LVT U515 ( .I(n946), .Z(o_data_bus[116]) );
  BUFFD6BWP30P140LVT U516 ( .I(n947), .Z(o_data_bus[115]) );
  BUFFD6BWP30P140LVT U517 ( .I(n948), .Z(o_data_bus[114]) );
  BUFFD6BWP30P140LVT U518 ( .I(n576), .Z(o_data_bus[486]) );
  BUFFD6BWP30P140LVT U519 ( .I(n949), .Z(o_data_bus[113]) );
  BUFFD6BWP30P140LVT U520 ( .I(n950), .Z(o_data_bus[112]) );
  BUFFD6BWP30P140LVT U521 ( .I(n575), .Z(o_data_bus[487]) );
  BUFFD6BWP30P140LVT U522 ( .I(n574), .Z(o_data_bus[488]) );
  BUFFD6BWP30P140LVT U523 ( .I(n951), .Z(o_data_bus[111]) );
  BUFFD6BWP30P140LVT U524 ( .I(n955), .Z(o_data_bus[107]) );
  BUFFD6BWP30P140LVT U525 ( .I(n956), .Z(o_data_bus[106]) );
  BUFFD6BWP30P140LVT U526 ( .I(n953), .Z(o_data_bus[109]) );
  BUFFD6BWP30P140LVT U527 ( .I(n952), .Z(o_data_bus[110]) );
  BUFFD6BWP30P140LVT U528 ( .I(n571), .Z(o_data_bus[491]) );
  BUFFD6BWP30P140LVT U529 ( .I(n535), .Z(o_valid[15]) );
  BUFFD6BWP30P140LVT U530 ( .I(n572), .Z(o_data_bus[490]) );
  BUFFD6BWP30P140LVT U531 ( .I(n958), .Z(o_data_bus[104]) );
  BUFFD6BWP30P140LVT U532 ( .I(n959), .Z(o_data_bus[103]) );
  BUFFD6BWP30P140LVT U533 ( .I(n573), .Z(o_data_bus[489]) );
  BUFFD6BWP30P140LVT U534 ( .I(n957), .Z(o_data_bus[105]) );
  BUFFD6BWP30P140LVT U535 ( .I(n570), .Z(o_data_bus[492]) );
  BUFFD6BWP30P140LVT U536 ( .I(n954), .Z(o_data_bus[108]) );
endmodule

