
module crossbar_one_hot_seq ( clk, rst, i_valid, i_data_bus, o_valid, 
        o_data_bus, i_en, i_cmd );
  input [31:0] i_valid;
  input [1023:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input [255:0] i_cmd;
  input clk, rst, i_en;
  wire   N542, N543, N544, N545, N546, N547, N548, N549, N550, N551, N552,
         N553, N554, N555, N556, N557, N558, N559, N560, N561, N562, N563,
         N564, N565, N566, N567, N568, N569, N570, N571, N572, N573, N574,
         N762, N763, N764, N765, N766, N767, N768, N769, N770, N771, N772,
         N773, N774, N775, N776, N777, N778, N779, N780, N781, N782, N783,
         N784, N785, N786, N787, N788, N789, N790, N791, N792, N793, N794,
         N982, N983, N984, N985, N986, N987, N988, N989, N990, N991, N992,
         N993, N994, N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003,
         N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013,
         N1014, N1202, N1203, N1204, N1205, N1206, N1207, N1208, N1209, N1210,
         N1211, N1212, N1213, N1214, N1215, N1216, N1217, N1218, N1219, N1220,
         N1221, N1222, N1223, N1224, N1225, N1226, N1227, N1228, N1229, N1230,
         N1231, N1232, N1233, N1234, N1422, N1423, N1424, N1425, N1426, N1427,
         N1428, N1429, N1430, N1431, N1432, N1433, N1434, N1435, N1436, N1437,
         N1438, N1439, N1440, N1441, N1442, N1443, N1444, N1445, N1446, N1447,
         N1448, N1449, N1450, N1451, N1452, N1453, N1454, N1642, N1643, N1644,
         N1645, N1646, N1647, N1648, N1649, N1650, N1651, N1652, N1653, N1654,
         N1655, N1656, N1657, N1658, N1659, N1660, N1661, N1662, N1663, N1664,
         N1665, N1666, N1667, N1668, N1669, N1670, N1671, N1672, N1673, N1674,
         N1862, N1863, N1864, N1865, N1866, N1867, N1868, N1869, N1870, N1871,
         N1872, N1873, N1874, N1875, N1876, N1877, N1878, N1879, N1880, N1881,
         N1882, N1883, N1884, N1885, N1886, N1887, N1888, N1889, N1890, N1891,
         N1892, N1893, N1894, N2082, N2083, N2084, N2085, N2086, N2087, N2088,
         N2089, N2090, N2091, N2092, N2093, N2094, N2095, N2096, N2097, N2098,
         N2099, N2100, N2101, N2102, N2103, N2104, N2105, N2106, N2107, N2108,
         N2109, N2110, N2111, N2112, N2113, N2114, N2228, N2229, N2230, N2231,
         N2232, N2233, N2234, N2235, N2236, N2237, N2238, N2239, N2240, N2241,
         N2242, N2243, N2244, N2245, N2246, N2247, N2248, N2249, N2250, N2251,
         N2252, N2253, N2254, N2255, N2256, N2257, N2258, N2259, N2260, N2444,
         N2445, N2446, N2447, N2448, N2449, N2450, N2451, N2452, N2453, N2454,
         N2455, N2456, N2457, N2458, N2459, N2460, N2461, N2462, N2463, N2464,
         N2465, N2466, N2467, N2468, N2469, N2470, N2471, N2472, N2473, N2474,
         N2475, N2476, N2660, N2661, N2662, N2663, N2664, N2665, N2666, N2667,
         N2668, N2669, N2670, N2671, N2672, N2673, N2674, N2675, N2676, N2677,
         N2678, N2679, N2680, N2681, N2682, N2683, N2684, N2685, N2686, N2687,
         N2688, N2689, N2690, N2691, N2692, N2876, N2877, N2878, N2879, N2880,
         N2881, N2882, N2883, N2884, N2885, N2886, N2887, N2888, N2889, N2890,
         N2891, N2892, N2893, N2894, N2895, N2896, N2897, N2898, N2899, N2900,
         N2901, N2902, N2903, N2904, N2905, N2906, N2907, N2908, N3092, N3093,
         N3094, N3095, N3096, N3097, N3098, N3099, N3100, N3101, N3102, N3103,
         N3104, N3105, N3106, N3107, N3108, N3109, N3110, N3111, N3112, N3113,
         N3114, N3115, N3116, N3117, N3118, N3119, N3120, N3121, N3122, N3123,
         N3124, N3308, N3309, N3310, N3311, N3312, N3313, N3314, N3315, N3316,
         N3317, N3318, N3319, N3320, N3321, N3322, N3323, N3324, N3325, N3326,
         N3327, N3328, N3329, N3330, N3331, N3332, N3333, N3334, N3335, N3336,
         N3337, N3338, N3339, N3340, N3524, N3525, N3526, N3527, N3528, N3529,
         N3530, N3531, N3532, N3533, N3534, N3535, N3536, N3537, N3538, N3539,
         N3540, N3541, N3542, N3543, N3544, N3545, N3546, N3547, N3548, N3549,
         N3550, N3551, N3552, N3553, N3554, N3555, N3556, N3740, N3741, N3742,
         N3743, N3744, N3745, N3746, N3747, N3748, N3749, N3750, N3751, N3752,
         N3753, N3754, N3755, N3756, N3757, N3758, N3759, N3760, N3761, N3762,
         N3763, N3764, N3765, N3766, N3767, N3768, N3769, N3770, N3771, N3772,
         N3956, N3957, N3958, N3959, N3960, N3961, N3962, N3963, N3964, N3965,
         N3966, N3967, N3968, N3969, N3970, N3971, N3972, N3973, N3974, N3975,
         N3976, N3977, N3978, N3979, N3980, N3981, N3982, N3983, N3984, N3985,
         N3986, N3987, N3988, N4102, N4103, N4104, N4105, N4106, N4107, N4108,
         N4109, N4110, N4111, N4112, N4113, N4114, N4115, N4116, N4117, N4118,
         N4119, N4120, N4121, N4122, N4123, N4124, N4125, N4126, N4127, N4128,
         N4129, N4130, N4131, N4132, N4133, N4134, N4318, N4319, N4320, N4321,
         N4322, N4323, N4324, N4325, N4326, N4327, N4328, N4329, N4330, N4331,
         N4332, N4333, N4334, N4335, N4336, N4337, N4338, N4339, N4340, N4341,
         N4342, N4343, N4344, N4345, N4346, N4347, N4348, N4349, N4350, N4534,
         N4535, N4536, N4537, N4538, N4539, N4540, N4541, N4542, N4543, N4544,
         N4545, N4546, N4547, N4548, N4549, N4550, N4551, N4552, N4553, N4554,
         N4555, N4556, N4557, N4558, N4559, N4560, N4561, N4562, N4563, N4564,
         N4565, N4566, N4750, N4751, N4752, N4753, N4754, N4755, N4756, N4757,
         N4758, N4759, N4760, N4761, N4762, N4763, N4764, N4765, N4766, N4767,
         N4768, N4769, N4770, N4771, N4772, N4773, N4774, N4775, N4776, N4777,
         N4778, N4779, N4780, N4781, N4782, N4966, N4967, N4968, N4969, N4970,
         N4971, N4972, N4973, N4974, N4975, N4976, N4977, N4978, N4979, N4980,
         N4981, N4982, N4983, N4984, N4985, N4986, N4987, N4988, N4989, N4990,
         N4991, N4992, N4993, N4994, N4995, N4996, N4997, N4998, N5182, N5183,
         N5184, N5185, N5186, N5187, N5188, N5189, N5190, N5191, N5192, N5193,
         N5194, N5195, N5196, N5197, N5198, N5199, N5200, N5201, N5202, N5203,
         N5204, N5205, N5206, N5207, N5208, N5209, N5210, N5211, N5212, N5213,
         N5214, N5398, N5399, N5400, N5401, N5402, N5403, N5404, N5405, N5406,
         N5407, N5408, N5409, N5410, N5411, N5412, N5413, N5414, N5415, N5416,
         N5417, N5418, N5419, N5420, N5421, N5422, N5423, N5424, N5425, N5426,
         N5427, N5428, N5429, N5430, N5614, N5615, N5616, N5617, N5618, N5619,
         N5620, N5621, N5622, N5623, N5624, N5625, N5626, N5627, N5628, N5629,
         N5630, N5631, N5632, N5633, N5634, N5635, N5636, N5637, N5638, N5639,
         N5640, N5641, N5642, N5643, N5644, N5645, N5646, N5830, N5831, N5832,
         N5833, N5834, N5835, N5836, N5837, N5838, N5839, N5840, N5841, N5842,
         N5843, N5844, N5845, N5846, N5847, N5848, N5849, N5850, N5851, N5852,
         N5853, N5854, N5855, N5856, N5857, N5858, N5859, N5860, N5861, N5862,
         N5976, N5977, N5978, N5979, N5980, N5981, N5982, N5983, N5984, N5985,
         N5986, N5987, N5988, N5989, N5990, N5991, N5992, N5993, N5994, N5995,
         N5996, N5997, N5998, N5999, N6000, N6001, N6002, N6003, N6004, N6005,
         N6006, N6007, N6008, N6192, N6193, N6194, N6195, N6196, N6197, N6198,
         N6199, N6200, N6201, N6202, N6203, N6204, N6205, N6206, N6207, N6208,
         N6209, N6210, N6211, N6212, N6213, N6214, N6215, N6216, N6217, N6218,
         N6219, N6220, N6221, N6222, N6223, N6224, N6408, N6409, N6410, N6411,
         N6412, N6413, N6414, N6415, N6416, N6417, N6418, N6419, N6420, N6421,
         N6422, N6423, N6424, N6425, N6426, N6427, N6428, N6429, N6430, N6431,
         N6432, N6433, N6434, N6435, N6436, N6437, N6438, N6439, N6440, N6624,
         N6625, N6626, N6627, N6628, N6629, N6630, N6631, N6632, N6633, N6634,
         N6635, N6636, N6637, N6638, N6639, N6640, N6641, N6642, N6643, N6644,
         N6645, N6646, N6647, N6648, N6649, N6650, N6651, N6652, N6653, N6654,
         N6655, N6656, N6840, N6841, N6842, N6843, N6844, N6845, N6846, N6847,
         N6848, N6849, N6850, N6851, N6852, N6853, N6854, N6855, N6856, N6857,
         N6858, N6859, N6860, N6861, N6862, N6863, N6864, N6865, N6866, N6867,
         N6868, N6869, N6870, N6871, N6872, N7056, N7057, N7058, N7059, N7060,
         N7061, N7062, N7063, N7064, N7065, N7066, N7067, N7068, N7069, N7070,
         N7071, N7072, N7073, N7074, N7075, N7076, N7077, N7078, N7079, N7080,
         N7081, N7082, N7083, N7084, N7085, N7086, N7087, N7088, N7272, N7273,
         N7274, N7275, N7276, N7277, N7278, N7279, N7280, N7281, N7282, N7283,
         N7284, N7285, N7286, N7287, N7288, N7289, N7290, N7291, N7292, N7293,
         N7294, N7295, N7296, N7297, N7298, N7299, N7300, N7301, N7302, N7303,
         N7304, N7488, N7489, N7490, N7491, N7492, N7493, N7494, N7495, N7496,
         N7497, N7498, N7499, N7500, N7501, N7502, N7503, N7504, N7505, N7506,
         N7507, N7508, N7509, N7510, N7511, N7512, N7513, N7514, N7515, N7516,
         N7517, N7518, N7519, N7520, N7704, N7705, N7706, N7707, N7708, N7709,
         N7710, N7711, N7712, N7713, N7714, N7715, N7716, N7717, N7718, N7719,
         N7720, N7721, N7722, N7723, N7724, N7725, N7726, N7727, N7728, N7729,
         N7730, N7731, N7732, N7733, N7734, N7735, N7736, N7850, N7851, N7852,
         N7853, N7854, N7855, N7856, N7857, N7858, N7859, N7860, N7861, N7862,
         N7863, N7864, N7865, N7866, N7867, N7868, N7869, N7870, N7871, N7872,
         N7873, N7874, N7875, N7876, N7877, N7878, N7879, N7880, N7881, N7882,
         N8066, N8067, N8068, N8069, N8070, N8071, N8072, N8073, N8074, N8075,
         N8076, N8077, N8078, N8079, N8080, N8081, N8082, N8083, N8084, N8085,
         N8086, N8087, N8088, N8089, N8090, N8091, N8092, N8093, N8094, N8095,
         N8096, N8097, N8098, N8282, N8283, N8284, N8285, N8286, N8287, N8288,
         N8289, N8290, N8291, N8292, N8293, N8294, N8295, N8296, N8297, N8298,
         N8299, N8300, N8301, N8302, N8303, N8304, N8305, N8306, N8307, N8308,
         N8309, N8310, N8311, N8312, N8313, N8314, N8498, N8499, N8500, N8501,
         N8502, N8503, N8504, N8505, N8506, N8507, N8508, N8509, N8510, N8511,
         N8512, N8513, N8514, N8515, N8516, N8517, N8518, N8519, N8520, N8521,
         N8522, N8523, N8524, N8525, N8526, N8527, N8528, N8529, N8530, N8714,
         N8715, N8716, N8717, N8718, N8719, N8720, N8721, N8722, N8723, N8724,
         N8725, N8726, N8727, N8728, N8729, N8730, N8731, N8732, N8733, N8734,
         N8735, N8736, N8737, N8738, N8739, N8740, N8741, N8742, N8743, N8744,
         N8745, N8746, N8930, N8931, N8932, N8933, N8934, N8935, N8936, N8937,
         N8938, N8939, N8940, N8941, N8942, N8943, N8944, N8945, N8946, N8947,
         N8948, N8949, N8950, N8951, N8952, N8953, N8954, N8955, N8956, N8957,
         N8958, N8959, N8960, N8961, N8962, N9146, N9147, N9148, N9149, N9150,
         N9151, N9152, N9153, N9154, N9155, N9156, N9157, N9158, N9159, N9160,
         N9161, N9162, N9163, N9164, N9165, N9166, N9167, N9168, N9169, N9170,
         N9171, N9172, N9173, N9174, N9175, N9176, N9177, N9178, N9362, N9363,
         N9364, N9365, N9366, N9367, N9368, N9369, N9370, N9371, N9372, N9373,
         N9374, N9375, N9376, N9377, N9378, N9379, N9380, N9381, N9382, N9383,
         N9384, N9385, N9386, N9387, N9388, N9389, N9390, N9391, N9392, N9393,
         N9394, N9578, N9579, N9580, N9581, N9582, N9583, N9584, N9585, N9586,
         N9587, N9588, N9589, N9590, N9591, N9592, N9593, N9594, N9595, N9596,
         N9597, N9598, N9599, N9600, N9601, N9602, N9603, N9604, N9605, N9606,
         N9607, N9608, N9609, N9610, N9724, N9725, N9726, N9727, N9728, N9729,
         N9730, N9731, N9732, N9733, N9734, N9735, N9736, N9737, N9738, N9739,
         N9740, N9741, N9742, N9743, N9744, N9745, N9746, N9747, N9748, N9749,
         N9750, N9751, N9752, N9753, N9754, N9755, N9756, N9940, N9941, N9942,
         N9943, N9944, N9945, N9946, N9947, N9948, N9949, N9950, N9951, N9952,
         N9953, N9954, N9955, N9956, N9957, N9958, N9959, N9960, N9961, N9962,
         N9963, N9964, N9965, N9966, N9967, N9968, N9969, N9970, N9971, N9972,
         N10156, N10157, N10158, N10159, N10160, N10161, N10162, N10163,
         N10164, N10165, N10166, N10167, N10168, N10169, N10170, N10171,
         N10172, N10173, N10174, N10175, N10176, N10177, N10178, N10179,
         N10180, N10181, N10182, N10183, N10184, N10185, N10186, N10187,
         N10188, N10372, N10373, N10374, N10375, N10376, N10377, N10378,
         N10379, N10380, N10381, N10382, N10383, N10384, N10385, N10386,
         N10387, N10388, N10389, N10390, N10391, N10392, N10393, N10394,
         N10395, N10396, N10397, N10398, N10399, N10400, N10401, N10402,
         N10403, N10404, N10588, N10589, N10590, N10591, N10592, N10593,
         N10594, N10595, N10596, N10597, N10598, N10599, N10600, N10601,
         N10602, N10603, N10604, N10605, N10606, N10607, N10608, N10609,
         N10610, N10611, N10612, N10613, N10614, N10615, N10616, N10617,
         N10618, N10619, N10620, N10804, N10805, N10806, N10807, N10808,
         N10809, N10810, N10811, N10812, N10813, N10814, N10815, N10816,
         N10817, N10818, N10819, N10820, N10821, N10822, N10823, N10824,
         N10825, N10826, N10827, N10828, N10829, N10830, N10831, N10832,
         N10833, N10834, N10835, N10836, N11020, N11021, N11022, N11023,
         N11024, N11025, N11026, N11027, N11028, N11029, N11030, N11031,
         N11032, N11033, N11034, N11035, N11036, N11037, N11038, N11039,
         N11040, N11041, N11042, N11043, N11044, N11045, N11046, N11047,
         N11048, N11049, N11050, N11051, N11052, N11236, N11237, N11238,
         N11239, N11240, N11241, N11242, N11243, N11244, N11245, N11246,
         N11247, N11248, N11249, N11250, N11251, N11252, N11253, N11254,
         N11255, N11256, N11257, N11258, N11259, N11260, N11261, N11262,
         N11263, N11264, N11265, N11266, N11267, N11268, N11452, N11453,
         N11454, N11455, N11456, N11457, N11458, N11459, N11460, N11461,
         N11462, N11463, N11464, N11465, N11466, N11467, N11468, N11469,
         N11470, N11471, N11472, N11473, N11474, N11475, N11476, N11477,
         N11478, N11479, N11480, N11481, N11482, N11483, N11484, N11598,
         N11599, N11600, N11601, N11602, N11603, N11604, N11605, N11606,
         N11607, N11608, N11609, N11610, N11611, N11612, N11613, N11614,
         N11615, N11616, N11617, N11618, N11619, N11620, N11621, N11622,
         N11623, N11624, N11625, N11626, N11627, N11628, N11629, N11630,
         N11814, N11815, N11816, N11817, N11818, N11819, N11820, N11821,
         N11822, N11823, N11824, N11825, N11826, N11827, N11828, N11829,
         N11830, N11831, N11832, N11833, N11834, N11835, N11836, N11837,
         N11838, N11839, N11840, N11841, N11842, N11843, N11844, N11845,
         N11846, N12030, N12031, N12032, N12033, N12034, N12035, N12036,
         N12037, N12038, N12039, N12040, N12041, N12042, N12043, N12044,
         N12045, N12046, N12047, N12048, N12049, N12050, N12051, N12052,
         N12053, N12054, N12055, N12056, N12057, N12058, N12059, N12060,
         N12061, N12062, N12246, N12247, N12248, N12249, N12250, N12251,
         N12252, N12253, N12254, N12255, N12256, N12257, N12258, N12259,
         N12260, N12261, N12262, N12263, N12264, N12265, N12266, N12267,
         N12268, N12269, N12270, N12271, N12272, N12273, N12274, N12275,
         N12276, N12277, N12278, N12462, N12463, N12464, N12465, N12466,
         N12467, N12468, N12469, N12470, N12471, N12472, N12473, N12474,
         N12475, N12476, N12477, N12478, N12479, N12480, N12481, N12482,
         N12483, N12484, N12485, N12486, N12487, N12488, N12489, N12490,
         N12491, N12492, N12493, N12494, N12678, N12679, N12680, N12681,
         N12682, N12683, N12684, N12685, N12686, N12687, N12688, N12689,
         N12690, N12691, N12692, N12693, N12694, N12695, N12696, N12697,
         N12698, N12699, N12700, N12701, N12702, N12703, N12704, N12705,
         N12706, N12707, N12708, N12709, N12710, N12894, N12895, N12896,
         N12897, N12898, N12899, N12900, N12901, N12902, N12903, N12904,
         N12905, N12906, N12907, N12908, N12909, N12910, N12911, N12912,
         N12913, N12914, N12915, N12916, N12917, N12918, N12919, N12920,
         N12921, N12922, N12923, N12924, N12925, N12926, N13110, N13111,
         N13112, N13113, N13114, N13115, N13116, N13117, N13118, N13119,
         N13120, N13121, N13122, N13123, N13124, N13125, N13126, N13127,
         N13128, N13129, N13130, N13131, N13132, N13133, N13134, N13135,
         N13136, N13137, N13138, N13139, N13140, N13141, N13142, N13326,
         N13327, N13328, N13329, N13330, N13331, N13332, N13333, N13334,
         N13335, N13336, N13337, N13338, N13339, N13340, N13341, N13342,
         N13343, N13344, N13345, N13346, N13347, N13348, N13349, N13350,
         N13351, N13352, N13353, N13354, N13355, N13356, N13357, N13358,
         N13472, N13473, N13474, N13475, N13476, N13477, N13478, N13479,
         N13480, N13481, N13482, N13483, N13484, N13485, N13486, N13487,
         N13488, N13489, N13490, N13491, N13492, N13493, N13494, N13495,
         N13496, N13497, N13498, N13499, N13500, N13501, N13502, N13503,
         N13504, N13688, N13689, N13690, N13691, N13692, N13693, N13694,
         N13695, N13696, N13697, N13698, N13699, N13700, N13701, N13702,
         N13703, N13704, N13705, N13706, N13707, N13708, N13709, N13710,
         N13711, N13712, N13713, N13714, N13715, N13716, N13717, N13718,
         N13719, N13720, N13904, N13905, N13906, N13907, N13908, N13909,
         N13910, N13911, N13912, N13913, N13914, N13915, N13916, N13917,
         N13918, N13919, N13920, N13921, N13922, N13923, N13924, N13925,
         N13926, N13927, N13928, N13929, N13930, N13931, N13932, N13933,
         N13934, N13935, N13936, N14120, N14121, N14122, N14123, N14124,
         N14125, N14126, N14127, N14128, N14129, N14130, N14131, N14132,
         N14133, N14134, N14135, N14136, N14137, N14138, N14139, N14140,
         N14141, N14142, N14143, N14144, N14145, N14146, N14147, N14148,
         N14149, N14150, N14151, N14152, N14336, N14337, N14338, N14339,
         N14340, N14341, N14342, N14343, N14344, N14345, N14346, N14347,
         N14348, N14349, N14350, N14351, N14352, N14353, N14354, N14355,
         N14356, N14357, N14358, N14359, N14360, N14361, N14362, N14363,
         N14364, N14365, N14366, N14367, N14368, N14552, N14553, N14554,
         N14555, N14556, N14557, N14558, N14559, N14560, N14561, N14562,
         N14563, N14564, N14565, N14566, N14567, N14568, N14569, N14570,
         N14571, N14572, N14573, N14574, N14575, N14576, N14577, N14578,
         N14579, N14580, N14581, N14582, N14583, N14584, N14768, N14769,
         N14770, N14771, N14772, N14773, N14774, N14775, N14776, N14777,
         N14778, N14779, N14780, N14781, N14782, N14783, N14784, N14785,
         N14786, N14787, N14788, N14789, N14790, N14791, N14792, N14793,
         N14794, N14795, N14796, N14797, N14798, N14799, N14800, N14984,
         N14985, N14986, N14987, N14988, N14989, N14990, N14991, N14992,
         N14993, N14994, N14995, N14996, N14997, N14998, N14999, N15000,
         N15001, N15002, N15003, N15004, N15005, N15006, N15007, N15008,
         N15009, N15010, N15011, N15012, N15013, N15014, N15015, N15016,
         N15200, N15201, N15202, N15203, N15204, N15205, N15206, N15207,
         N15208, N15209, N15210, N15211, N15212, N15213, N15214, N15215,
         N15216, N15217, N15218, N15219, N15220, N15221, N15222, N15223,
         N15224, N15225, N15226, N15227, N15228, N15229, N15230, N15231,
         N15232, N15346, N15347, N15348, N15349, N15350, N15351, N15352,
         N15353, N15354, N15355, N15356, N15357, N15358, N15359, N15360,
         N15361, N15362, N15363, N15364, N15365, N15366, N15367, N15368,
         N15369, N15370, N15371, N15372, N15373, N15374, N15375, N15376,
         N15377, N15378, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767;
  wire   [2047:0] inner_first_stage_data_reg;
  wire   [63:0] inner_first_stage_valid_reg;

  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_31_ ( .D(N574), .CP(clk), 
        .Q(inner_first_stage_data_reg[31]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_30_ ( .D(N573), .CP(clk), 
        .Q(inner_first_stage_data_reg[30]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_29_ ( .D(N572), .CP(clk), 
        .Q(inner_first_stage_data_reg[29]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_28_ ( .D(N571), .CP(clk), 
        .Q(inner_first_stage_data_reg[28]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_27_ ( .D(N570), .CP(clk), 
        .Q(inner_first_stage_data_reg[27]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_26_ ( .D(N569), .CP(clk), 
        .Q(inner_first_stage_data_reg[26]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_25_ ( .D(N568), .CP(clk), 
        .Q(inner_first_stage_data_reg[25]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_24_ ( .D(N567), .CP(clk), 
        .Q(inner_first_stage_data_reg[24]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_23_ ( .D(N566), .CP(clk), 
        .Q(inner_first_stage_data_reg[23]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_22_ ( .D(N565), .CP(clk), 
        .Q(inner_first_stage_data_reg[22]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_21_ ( .D(N564), .CP(clk), 
        .Q(inner_first_stage_data_reg[21]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_20_ ( .D(N563), .CP(clk), 
        .Q(inner_first_stage_data_reg[20]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_19_ ( .D(N562), .CP(clk), 
        .Q(inner_first_stage_data_reg[19]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_18_ ( .D(N561), .CP(clk), 
        .Q(inner_first_stage_data_reg[18]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_17_ ( .D(N560), .CP(clk), 
        .Q(inner_first_stage_data_reg[17]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_16_ ( .D(N559), .CP(clk), 
        .Q(inner_first_stage_data_reg[16]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_15_ ( .D(N558), .CP(clk), 
        .Q(inner_first_stage_data_reg[15]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_14_ ( .D(N557), .CP(clk), 
        .Q(inner_first_stage_data_reg[14]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_13_ ( .D(N556), .CP(clk), 
        .Q(inner_first_stage_data_reg[13]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_12_ ( .D(N555), .CP(clk), 
        .Q(inner_first_stage_data_reg[12]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_11_ ( .D(N554), .CP(clk), 
        .Q(inner_first_stage_data_reg[11]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_10_ ( .D(N553), .CP(clk), 
        .Q(inner_first_stage_data_reg[10]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_9_ ( .D(N552), .CP(clk), 
        .Q(inner_first_stage_data_reg[9]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_8_ ( .D(N551), .CP(clk), 
        .Q(inner_first_stage_data_reg[8]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_7_ ( .D(N550), .CP(clk), 
        .Q(inner_first_stage_data_reg[7]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_6_ ( .D(N549), .CP(clk), 
        .Q(inner_first_stage_data_reg[6]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_5_ ( .D(N548), .CP(clk), 
        .Q(inner_first_stage_data_reg[5]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_4_ ( .D(N547), .CP(clk), 
        .Q(inner_first_stage_data_reg[4]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_3_ ( .D(N546), .CP(clk), 
        .Q(inner_first_stage_data_reg[3]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2_ ( .D(N545), .CP(clk), 
        .Q(inner_first_stage_data_reg[2]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1_ ( .D(N544), .CP(clk), 
        .Q(inner_first_stage_data_reg[1]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_0_ ( .D(N543), .CP(clk), 
        .Q(inner_first_stage_data_reg[0]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_0_ ( .D(N542), .CP(clk), 
        .Q(inner_first_stage_valid_reg[0]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_63_ ( .D(N794), .CP(clk), 
        .Q(inner_first_stage_data_reg[63]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_62_ ( .D(N793), .CP(clk), 
        .Q(inner_first_stage_data_reg[62]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_61_ ( .D(N792), .CP(clk), 
        .Q(inner_first_stage_data_reg[61]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_60_ ( .D(N791), .CP(clk), 
        .Q(inner_first_stage_data_reg[60]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_59_ ( .D(N790), .CP(clk), 
        .Q(inner_first_stage_data_reg[59]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_58_ ( .D(N789), .CP(clk), 
        .Q(inner_first_stage_data_reg[58]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_57_ ( .D(N788), .CP(clk), 
        .Q(inner_first_stage_data_reg[57]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_56_ ( .D(N787), .CP(clk), 
        .Q(inner_first_stage_data_reg[56]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_55_ ( .D(N786), .CP(clk), 
        .Q(inner_first_stage_data_reg[55]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_54_ ( .D(N785), .CP(clk), 
        .Q(inner_first_stage_data_reg[54]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_53_ ( .D(N784), .CP(clk), 
        .Q(inner_first_stage_data_reg[53]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_52_ ( .D(N783), .CP(clk), 
        .Q(inner_first_stage_data_reg[52]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_51_ ( .D(N782), .CP(clk), 
        .Q(inner_first_stage_data_reg[51]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_50_ ( .D(N781), .CP(clk), 
        .Q(inner_first_stage_data_reg[50]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_49_ ( .D(N780), .CP(clk), 
        .Q(inner_first_stage_data_reg[49]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_48_ ( .D(N779), .CP(clk), 
        .Q(inner_first_stage_data_reg[48]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_47_ ( .D(N778), .CP(clk), 
        .Q(inner_first_stage_data_reg[47]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_46_ ( .D(N777), .CP(clk), 
        .Q(inner_first_stage_data_reg[46]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_45_ ( .D(N776), .CP(clk), 
        .Q(inner_first_stage_data_reg[45]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_44_ ( .D(N775), .CP(clk), 
        .Q(inner_first_stage_data_reg[44]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_43_ ( .D(N774), .CP(clk), 
        .Q(inner_first_stage_data_reg[43]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_42_ ( .D(N773), .CP(clk), 
        .Q(inner_first_stage_data_reg[42]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_41_ ( .D(N772), .CP(clk), 
        .Q(inner_first_stage_data_reg[41]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_40_ ( .D(N771), .CP(clk), 
        .Q(inner_first_stage_data_reg[40]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_39_ ( .D(N770), .CP(clk), 
        .Q(inner_first_stage_data_reg[39]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_38_ ( .D(N769), .CP(clk), 
        .Q(inner_first_stage_data_reg[38]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_37_ ( .D(N768), .CP(clk), 
        .Q(inner_first_stage_data_reg[37]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_36_ ( .D(N767), .CP(clk), 
        .Q(inner_first_stage_data_reg[36]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_35_ ( .D(N766), .CP(clk), 
        .Q(inner_first_stage_data_reg[35]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_34_ ( .D(N765), .CP(clk), 
        .Q(inner_first_stage_data_reg[34]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_33_ ( .D(N764), .CP(clk), 
        .Q(inner_first_stage_data_reg[33]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_32_ ( .D(N763), .CP(clk), 
        .Q(inner_first_stage_data_reg[32]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_1_ ( .D(N762), .CP(clk), 
        .Q(inner_first_stage_valid_reg[1]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_95_ ( .D(N1014), .CP(clk), 
        .Q(inner_first_stage_data_reg[95]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_94_ ( .D(N1013), .CP(clk), 
        .Q(inner_first_stage_data_reg[94]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_93_ ( .D(N1012), .CP(clk), 
        .Q(inner_first_stage_data_reg[93]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_92_ ( .D(N1011), .CP(clk), 
        .Q(inner_first_stage_data_reg[92]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_91_ ( .D(N1010), .CP(clk), 
        .Q(inner_first_stage_data_reg[91]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_90_ ( .D(N1009), .CP(clk), 
        .Q(inner_first_stage_data_reg[90]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_89_ ( .D(N1008), .CP(clk), 
        .Q(inner_first_stage_data_reg[89]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_88_ ( .D(N1007), .CP(clk), 
        .Q(inner_first_stage_data_reg[88]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_87_ ( .D(N1006), .CP(clk), 
        .Q(inner_first_stage_data_reg[87]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_86_ ( .D(N1005), .CP(clk), 
        .Q(inner_first_stage_data_reg[86]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_85_ ( .D(N1004), .CP(clk), 
        .Q(inner_first_stage_data_reg[85]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_84_ ( .D(N1003), .CP(clk), 
        .Q(inner_first_stage_data_reg[84]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_83_ ( .D(N1002), .CP(clk), 
        .Q(inner_first_stage_data_reg[83]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_82_ ( .D(N1001), .CP(clk), 
        .Q(inner_first_stage_data_reg[82]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_81_ ( .D(N1000), .CP(clk), 
        .Q(inner_first_stage_data_reg[81]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_80_ ( .D(N999), .CP(clk), 
        .Q(inner_first_stage_data_reg[80]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_79_ ( .D(N998), .CP(clk), 
        .Q(inner_first_stage_data_reg[79]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_78_ ( .D(N997), .CP(clk), 
        .Q(inner_first_stage_data_reg[78]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_77_ ( .D(N996), .CP(clk), 
        .Q(inner_first_stage_data_reg[77]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_76_ ( .D(N995), .CP(clk), 
        .Q(inner_first_stage_data_reg[76]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_75_ ( .D(N994), .CP(clk), 
        .Q(inner_first_stage_data_reg[75]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_74_ ( .D(N993), .CP(clk), 
        .Q(inner_first_stage_data_reg[74]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_73_ ( .D(N992), .CP(clk), 
        .Q(inner_first_stage_data_reg[73]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_72_ ( .D(N991), .CP(clk), 
        .Q(inner_first_stage_data_reg[72]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_71_ ( .D(N990), .CP(clk), 
        .Q(inner_first_stage_data_reg[71]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_70_ ( .D(N989), .CP(clk), 
        .Q(inner_first_stage_data_reg[70]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_69_ ( .D(N988), .CP(clk), 
        .Q(inner_first_stage_data_reg[69]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_68_ ( .D(N987), .CP(clk), 
        .Q(inner_first_stage_data_reg[68]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_67_ ( .D(N986), .CP(clk), 
        .Q(inner_first_stage_data_reg[67]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_66_ ( .D(N985), .CP(clk), 
        .Q(inner_first_stage_data_reg[66]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_65_ ( .D(N984), .CP(clk), 
        .Q(inner_first_stage_data_reg[65]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_64_ ( .D(N983), .CP(clk), 
        .Q(inner_first_stage_data_reg[64]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_2_ ( .D(N982), .CP(clk), 
        .Q(inner_first_stage_valid_reg[2]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_127_ ( .D(N1234), .CP(clk), 
        .Q(inner_first_stage_data_reg[127]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_126_ ( .D(N1233), .CP(clk), 
        .Q(inner_first_stage_data_reg[126]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_125_ ( .D(N1232), .CP(clk), 
        .Q(inner_first_stage_data_reg[125]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_124_ ( .D(N1231), .CP(clk), 
        .Q(inner_first_stage_data_reg[124]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_123_ ( .D(N1230), .CP(clk), 
        .Q(inner_first_stage_data_reg[123]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_122_ ( .D(N1229), .CP(clk), 
        .Q(inner_first_stage_data_reg[122]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_121_ ( .D(N1228), .CP(clk), 
        .Q(inner_first_stage_data_reg[121]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_120_ ( .D(N1227), .CP(clk), 
        .Q(inner_first_stage_data_reg[120]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_119_ ( .D(N1226), .CP(clk), 
        .Q(inner_first_stage_data_reg[119]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_118_ ( .D(N1225), .CP(clk), 
        .Q(inner_first_stage_data_reg[118]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_117_ ( .D(N1224), .CP(clk), 
        .Q(inner_first_stage_data_reg[117]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_116_ ( .D(N1223), .CP(clk), 
        .Q(inner_first_stage_data_reg[116]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_115_ ( .D(N1222), .CP(clk), 
        .Q(inner_first_stage_data_reg[115]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_114_ ( .D(N1221), .CP(clk), 
        .Q(inner_first_stage_data_reg[114]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_113_ ( .D(N1220), .CP(clk), 
        .Q(inner_first_stage_data_reg[113]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_112_ ( .D(N1219), .CP(clk), 
        .Q(inner_first_stage_data_reg[112]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_111_ ( .D(N1218), .CP(clk), 
        .Q(inner_first_stage_data_reg[111]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_110_ ( .D(N1217), .CP(clk), 
        .Q(inner_first_stage_data_reg[110]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_109_ ( .D(N1216), .CP(clk), 
        .Q(inner_first_stage_data_reg[109]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_108_ ( .D(N1215), .CP(clk), 
        .Q(inner_first_stage_data_reg[108]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_107_ ( .D(N1214), .CP(clk), 
        .Q(inner_first_stage_data_reg[107]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_106_ ( .D(N1213), .CP(clk), 
        .Q(inner_first_stage_data_reg[106]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_105_ ( .D(N1212), .CP(clk), 
        .Q(inner_first_stage_data_reg[105]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_104_ ( .D(N1211), .CP(clk), 
        .Q(inner_first_stage_data_reg[104]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_103_ ( .D(N1210), .CP(clk), 
        .Q(inner_first_stage_data_reg[103]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_102_ ( .D(N1209), .CP(clk), 
        .Q(inner_first_stage_data_reg[102]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_101_ ( .D(N1208), .CP(clk), 
        .Q(inner_first_stage_data_reg[101]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_100_ ( .D(N1207), .CP(clk), 
        .Q(inner_first_stage_data_reg[100]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_99_ ( .D(N1206), .CP(clk), 
        .Q(inner_first_stage_data_reg[99]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_98_ ( .D(N1205), .CP(clk), 
        .Q(inner_first_stage_data_reg[98]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_97_ ( .D(N1204), .CP(clk), 
        .Q(inner_first_stage_data_reg[97]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_96_ ( .D(N1203), .CP(clk), 
        .Q(inner_first_stage_data_reg[96]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_3_ ( .D(N1202), .CP(clk), 
        .Q(inner_first_stage_valid_reg[3]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_159_ ( .D(N1454), .CP(clk), 
        .Q(inner_first_stage_data_reg[159]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_158_ ( .D(N1453), .CP(clk), 
        .Q(inner_first_stage_data_reg[158]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_157_ ( .D(N1452), .CP(clk), 
        .Q(inner_first_stage_data_reg[157]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_156_ ( .D(N1451), .CP(clk), 
        .Q(inner_first_stage_data_reg[156]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_155_ ( .D(N1450), .CP(clk), 
        .Q(inner_first_stage_data_reg[155]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_154_ ( .D(N1449), .CP(clk), 
        .Q(inner_first_stage_data_reg[154]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_153_ ( .D(N1448), .CP(clk), 
        .Q(inner_first_stage_data_reg[153]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_152_ ( .D(N1447), .CP(clk), 
        .Q(inner_first_stage_data_reg[152]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_151_ ( .D(N1446), .CP(clk), 
        .Q(inner_first_stage_data_reg[151]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_150_ ( .D(N1445), .CP(clk), 
        .Q(inner_first_stage_data_reg[150]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_149_ ( .D(N1444), .CP(clk), 
        .Q(inner_first_stage_data_reg[149]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_148_ ( .D(N1443), .CP(clk), 
        .Q(inner_first_stage_data_reg[148]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_147_ ( .D(N1442), .CP(clk), 
        .Q(inner_first_stage_data_reg[147]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_146_ ( .D(N1441), .CP(clk), 
        .Q(inner_first_stage_data_reg[146]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_145_ ( .D(N1440), .CP(clk), 
        .Q(inner_first_stage_data_reg[145]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_144_ ( .D(N1439), .CP(clk), 
        .Q(inner_first_stage_data_reg[144]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_143_ ( .D(N1438), .CP(clk), 
        .Q(inner_first_stage_data_reg[143]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_142_ ( .D(N1437), .CP(clk), 
        .Q(inner_first_stage_data_reg[142]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_141_ ( .D(N1436), .CP(clk), 
        .Q(inner_first_stage_data_reg[141]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_140_ ( .D(N1435), .CP(clk), 
        .Q(inner_first_stage_data_reg[140]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_139_ ( .D(N1434), .CP(clk), 
        .Q(inner_first_stage_data_reg[139]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_138_ ( .D(N1433), .CP(clk), 
        .Q(inner_first_stage_data_reg[138]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_137_ ( .D(N1432), .CP(clk), 
        .Q(inner_first_stage_data_reg[137]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_136_ ( .D(N1431), .CP(clk), 
        .Q(inner_first_stage_data_reg[136]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_135_ ( .D(N1430), .CP(clk), 
        .Q(inner_first_stage_data_reg[135]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_134_ ( .D(N1429), .CP(clk), 
        .Q(inner_first_stage_data_reg[134]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_133_ ( .D(N1428), .CP(clk), 
        .Q(inner_first_stage_data_reg[133]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_132_ ( .D(N1427), .CP(clk), 
        .Q(inner_first_stage_data_reg[132]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_131_ ( .D(N1426), .CP(clk), 
        .Q(inner_first_stage_data_reg[131]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_130_ ( .D(N1425), .CP(clk), 
        .Q(inner_first_stage_data_reg[130]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_129_ ( .D(N1424), .CP(clk), 
        .Q(inner_first_stage_data_reg[129]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_128_ ( .D(N1423), .CP(clk), 
        .Q(inner_first_stage_data_reg[128]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_4_ ( .D(N1422), .CP(clk), 
        .Q(inner_first_stage_valid_reg[4]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_191_ ( .D(N1674), .CP(clk), 
        .Q(inner_first_stage_data_reg[191]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_190_ ( .D(N1673), .CP(clk), 
        .Q(inner_first_stage_data_reg[190]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_189_ ( .D(N1672), .CP(clk), 
        .Q(inner_first_stage_data_reg[189]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_188_ ( .D(N1671), .CP(clk), 
        .Q(inner_first_stage_data_reg[188]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_187_ ( .D(N1670), .CP(clk), 
        .Q(inner_first_stage_data_reg[187]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_186_ ( .D(N1669), .CP(clk), 
        .Q(inner_first_stage_data_reg[186]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_185_ ( .D(N1668), .CP(clk), 
        .Q(inner_first_stage_data_reg[185]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_184_ ( .D(N1667), .CP(clk), 
        .Q(inner_first_stage_data_reg[184]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_183_ ( .D(N1666), .CP(clk), 
        .Q(inner_first_stage_data_reg[183]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_182_ ( .D(N1665), .CP(clk), 
        .Q(inner_first_stage_data_reg[182]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_181_ ( .D(N1664), .CP(clk), 
        .Q(inner_first_stage_data_reg[181]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_180_ ( .D(N1663), .CP(clk), 
        .Q(inner_first_stage_data_reg[180]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_179_ ( .D(N1662), .CP(clk), 
        .Q(inner_first_stage_data_reg[179]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_178_ ( .D(N1661), .CP(clk), 
        .Q(inner_first_stage_data_reg[178]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_177_ ( .D(N1660), .CP(clk), 
        .Q(inner_first_stage_data_reg[177]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_176_ ( .D(N1659), .CP(clk), 
        .Q(inner_first_stage_data_reg[176]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_175_ ( .D(N1658), .CP(clk), 
        .Q(inner_first_stage_data_reg[175]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_174_ ( .D(N1657), .CP(clk), 
        .Q(inner_first_stage_data_reg[174]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_173_ ( .D(N1656), .CP(clk), 
        .Q(inner_first_stage_data_reg[173]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_172_ ( .D(N1655), .CP(clk), 
        .Q(inner_first_stage_data_reg[172]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_171_ ( .D(N1654), .CP(clk), 
        .Q(inner_first_stage_data_reg[171]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_170_ ( .D(N1653), .CP(clk), 
        .Q(inner_first_stage_data_reg[170]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_169_ ( .D(N1652), .CP(clk), 
        .Q(inner_first_stage_data_reg[169]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_168_ ( .D(N1651), .CP(clk), 
        .Q(inner_first_stage_data_reg[168]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_167_ ( .D(N1650), .CP(clk), 
        .Q(inner_first_stage_data_reg[167]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_166_ ( .D(N1649), .CP(clk), 
        .Q(inner_first_stage_data_reg[166]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_165_ ( .D(N1648), .CP(clk), 
        .Q(inner_first_stage_data_reg[165]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_164_ ( .D(N1647), .CP(clk), 
        .Q(inner_first_stage_data_reg[164]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_163_ ( .D(N1646), .CP(clk), 
        .Q(inner_first_stage_data_reg[163]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_162_ ( .D(N1645), .CP(clk), 
        .Q(inner_first_stage_data_reg[162]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_161_ ( .D(N1644), .CP(clk), 
        .Q(inner_first_stage_data_reg[161]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_160_ ( .D(N1643), .CP(clk), 
        .Q(inner_first_stage_data_reg[160]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_5_ ( .D(N1642), .CP(clk), 
        .Q(inner_first_stage_valid_reg[5]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_223_ ( .D(N1894), .CP(clk), 
        .Q(inner_first_stage_data_reg[223]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_222_ ( .D(N1893), .CP(clk), 
        .Q(inner_first_stage_data_reg[222]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_221_ ( .D(N1892), .CP(clk), 
        .Q(inner_first_stage_data_reg[221]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_220_ ( .D(N1891), .CP(clk), 
        .Q(inner_first_stage_data_reg[220]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_219_ ( .D(N1890), .CP(clk), 
        .Q(inner_first_stage_data_reg[219]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_218_ ( .D(N1889), .CP(clk), 
        .Q(inner_first_stage_data_reg[218]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_217_ ( .D(N1888), .CP(clk), 
        .Q(inner_first_stage_data_reg[217]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_216_ ( .D(N1887), .CP(clk), 
        .Q(inner_first_stage_data_reg[216]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_215_ ( .D(N1886), .CP(clk), 
        .Q(inner_first_stage_data_reg[215]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_214_ ( .D(N1885), .CP(clk), 
        .Q(inner_first_stage_data_reg[214]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_213_ ( .D(N1884), .CP(clk), 
        .Q(inner_first_stage_data_reg[213]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_212_ ( .D(N1883), .CP(clk), 
        .Q(inner_first_stage_data_reg[212]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_211_ ( .D(N1882), .CP(clk), 
        .Q(inner_first_stage_data_reg[211]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_210_ ( .D(N1881), .CP(clk), 
        .Q(inner_first_stage_data_reg[210]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_209_ ( .D(N1880), .CP(clk), 
        .Q(inner_first_stage_data_reg[209]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_208_ ( .D(N1879), .CP(clk), 
        .Q(inner_first_stage_data_reg[208]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_207_ ( .D(N1878), .CP(clk), 
        .Q(inner_first_stage_data_reg[207]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_206_ ( .D(N1877), .CP(clk), 
        .Q(inner_first_stage_data_reg[206]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_205_ ( .D(N1876), .CP(clk), 
        .Q(inner_first_stage_data_reg[205]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_204_ ( .D(N1875), .CP(clk), 
        .Q(inner_first_stage_data_reg[204]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_203_ ( .D(N1874), .CP(clk), 
        .Q(inner_first_stage_data_reg[203]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_202_ ( .D(N1873), .CP(clk), 
        .Q(inner_first_stage_data_reg[202]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_201_ ( .D(N1872), .CP(clk), 
        .Q(inner_first_stage_data_reg[201]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_200_ ( .D(N1871), .CP(clk), 
        .Q(inner_first_stage_data_reg[200]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_199_ ( .D(N1870), .CP(clk), 
        .Q(inner_first_stage_data_reg[199]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_198_ ( .D(N1869), .CP(clk), 
        .Q(inner_first_stage_data_reg[198]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_197_ ( .D(N1868), .CP(clk), 
        .Q(inner_first_stage_data_reg[197]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_196_ ( .D(N1867), .CP(clk), 
        .Q(inner_first_stage_data_reg[196]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_195_ ( .D(N1866), .CP(clk), 
        .Q(inner_first_stage_data_reg[195]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_194_ ( .D(N1865), .CP(clk), 
        .Q(inner_first_stage_data_reg[194]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_193_ ( .D(N1864), .CP(clk), 
        .Q(inner_first_stage_data_reg[193]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_192_ ( .D(N1863), .CP(clk), 
        .Q(inner_first_stage_data_reg[192]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_6_ ( .D(N1862), .CP(clk), 
        .Q(inner_first_stage_valid_reg[6]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_255_ ( .D(N2114), .CP(clk), 
        .Q(inner_first_stage_data_reg[255]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_254_ ( .D(N2113), .CP(clk), 
        .Q(inner_first_stage_data_reg[254]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_253_ ( .D(N2112), .CP(clk), 
        .Q(inner_first_stage_data_reg[253]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_252_ ( .D(N2111), .CP(clk), 
        .Q(inner_first_stage_data_reg[252]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_251_ ( .D(N2110), .CP(clk), 
        .Q(inner_first_stage_data_reg[251]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_250_ ( .D(N2109), .CP(clk), 
        .Q(inner_first_stage_data_reg[250]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_249_ ( .D(N2108), .CP(clk), 
        .Q(inner_first_stage_data_reg[249]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_248_ ( .D(N2107), .CP(clk), 
        .Q(inner_first_stage_data_reg[248]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_247_ ( .D(N2106), .CP(clk), 
        .Q(inner_first_stage_data_reg[247]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_246_ ( .D(N2105), .CP(clk), 
        .Q(inner_first_stage_data_reg[246]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_245_ ( .D(N2104), .CP(clk), 
        .Q(inner_first_stage_data_reg[245]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_244_ ( .D(N2103), .CP(clk), 
        .Q(inner_first_stage_data_reg[244]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_243_ ( .D(N2102), .CP(clk), 
        .Q(inner_first_stage_data_reg[243]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_242_ ( .D(N2101), .CP(clk), 
        .Q(inner_first_stage_data_reg[242]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_241_ ( .D(N2100), .CP(clk), 
        .Q(inner_first_stage_data_reg[241]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_240_ ( .D(N2099), .CP(clk), 
        .Q(inner_first_stage_data_reg[240]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_239_ ( .D(N2098), .CP(clk), 
        .Q(inner_first_stage_data_reg[239]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_238_ ( .D(N2097), .CP(clk), 
        .Q(inner_first_stage_data_reg[238]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_237_ ( .D(N2096), .CP(clk), 
        .Q(inner_first_stage_data_reg[237]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_236_ ( .D(N2095), .CP(clk), 
        .Q(inner_first_stage_data_reg[236]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_235_ ( .D(N2094), .CP(clk), 
        .Q(inner_first_stage_data_reg[235]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_234_ ( .D(N2093), .CP(clk), 
        .Q(inner_first_stage_data_reg[234]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_233_ ( .D(N2092), .CP(clk), 
        .Q(inner_first_stage_data_reg[233]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_232_ ( .D(N2091), .CP(clk), 
        .Q(inner_first_stage_data_reg[232]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_231_ ( .D(N2090), .CP(clk), 
        .Q(inner_first_stage_data_reg[231]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_230_ ( .D(N2089), .CP(clk), 
        .Q(inner_first_stage_data_reg[230]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_229_ ( .D(N2088), .CP(clk), 
        .Q(inner_first_stage_data_reg[229]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_228_ ( .D(N2087), .CP(clk), 
        .Q(inner_first_stage_data_reg[228]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_227_ ( .D(N2086), .CP(clk), 
        .Q(inner_first_stage_data_reg[227]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_226_ ( .D(N2085), .CP(clk), 
        .Q(inner_first_stage_data_reg[226]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_225_ ( .D(N2084), .CP(clk), 
        .Q(inner_first_stage_data_reg[225]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_224_ ( .D(N2083), .CP(clk), 
        .Q(inner_first_stage_data_reg[224]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_7_ ( .D(N2082), .CP(clk), 
        .Q(inner_first_stage_valid_reg[7]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_287_ ( .D(N2476), .CP(clk), 
        .Q(inner_first_stage_data_reg[287]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_286_ ( .D(N2475), .CP(clk), 
        .Q(inner_first_stage_data_reg[286]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_285_ ( .D(N2474), .CP(clk), 
        .Q(inner_first_stage_data_reg[285]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_284_ ( .D(N2473), .CP(clk), 
        .Q(inner_first_stage_data_reg[284]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_283_ ( .D(N2472), .CP(clk), 
        .Q(inner_first_stage_data_reg[283]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_282_ ( .D(N2471), .CP(clk), 
        .Q(inner_first_stage_data_reg[282]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_281_ ( .D(N2470), .CP(clk), 
        .Q(inner_first_stage_data_reg[281]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_280_ ( .D(N2469), .CP(clk), 
        .Q(inner_first_stage_data_reg[280]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_279_ ( .D(N2468), .CP(clk), 
        .Q(inner_first_stage_data_reg[279]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_278_ ( .D(N2467), .CP(clk), 
        .Q(inner_first_stage_data_reg[278]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_277_ ( .D(N2466), .CP(clk), 
        .Q(inner_first_stage_data_reg[277]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_276_ ( .D(N2465), .CP(clk), 
        .Q(inner_first_stage_data_reg[276]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_275_ ( .D(N2464), .CP(clk), 
        .Q(inner_first_stage_data_reg[275]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_274_ ( .D(N2463), .CP(clk), 
        .Q(inner_first_stage_data_reg[274]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_273_ ( .D(N2462), .CP(clk), 
        .Q(inner_first_stage_data_reg[273]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_272_ ( .D(N2461), .CP(clk), 
        .Q(inner_first_stage_data_reg[272]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_271_ ( .D(N2460), .CP(clk), 
        .Q(inner_first_stage_data_reg[271]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_270_ ( .D(N2459), .CP(clk), 
        .Q(inner_first_stage_data_reg[270]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_269_ ( .D(N2458), .CP(clk), 
        .Q(inner_first_stage_data_reg[269]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_268_ ( .D(N2457), .CP(clk), 
        .Q(inner_first_stage_data_reg[268]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_267_ ( .D(N2456), .CP(clk), 
        .Q(inner_first_stage_data_reg[267]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_266_ ( .D(N2455), .CP(clk), 
        .Q(inner_first_stage_data_reg[266]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_265_ ( .D(N2454), .CP(clk), 
        .Q(inner_first_stage_data_reg[265]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_264_ ( .D(N2453), .CP(clk), 
        .Q(inner_first_stage_data_reg[264]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_263_ ( .D(N2452), .CP(clk), 
        .Q(inner_first_stage_data_reg[263]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_262_ ( .D(N2451), .CP(clk), 
        .Q(inner_first_stage_data_reg[262]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_261_ ( .D(N2450), .CP(clk), 
        .Q(inner_first_stage_data_reg[261]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_260_ ( .D(N2449), .CP(clk), 
        .Q(inner_first_stage_data_reg[260]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_259_ ( .D(N2448), .CP(clk), 
        .Q(inner_first_stage_data_reg[259]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_258_ ( .D(N2447), .CP(clk), 
        .Q(inner_first_stage_data_reg[258]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_257_ ( .D(N2446), .CP(clk), 
        .Q(inner_first_stage_data_reg[257]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_256_ ( .D(N2445), .CP(clk), 
        .Q(inner_first_stage_data_reg[256]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_8_ ( .D(N2444), .CP(clk), 
        .Q(inner_first_stage_valid_reg[8]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_319_ ( .D(N2692), .CP(clk), 
        .Q(inner_first_stage_data_reg[319]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_318_ ( .D(N2691), .CP(clk), 
        .Q(inner_first_stage_data_reg[318]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_317_ ( .D(N2690), .CP(clk), 
        .Q(inner_first_stage_data_reg[317]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_316_ ( .D(N2689), .CP(clk), 
        .Q(inner_first_stage_data_reg[316]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_315_ ( .D(N2688), .CP(clk), 
        .Q(inner_first_stage_data_reg[315]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_314_ ( .D(N2687), .CP(clk), 
        .Q(inner_first_stage_data_reg[314]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_313_ ( .D(N2686), .CP(clk), 
        .Q(inner_first_stage_data_reg[313]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_312_ ( .D(N2685), .CP(clk), 
        .Q(inner_first_stage_data_reg[312]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_311_ ( .D(N2684), .CP(clk), 
        .Q(inner_first_stage_data_reg[311]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_310_ ( .D(N2683), .CP(clk), 
        .Q(inner_first_stage_data_reg[310]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_309_ ( .D(N2682), .CP(clk), 
        .Q(inner_first_stage_data_reg[309]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_308_ ( .D(N2681), .CP(clk), 
        .Q(inner_first_stage_data_reg[308]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_307_ ( .D(N2680), .CP(clk), 
        .Q(inner_first_stage_data_reg[307]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_306_ ( .D(N2679), .CP(clk), 
        .Q(inner_first_stage_data_reg[306]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_305_ ( .D(N2678), .CP(clk), 
        .Q(inner_first_stage_data_reg[305]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_304_ ( .D(N2677), .CP(clk), 
        .Q(inner_first_stage_data_reg[304]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_303_ ( .D(N2676), .CP(clk), 
        .Q(inner_first_stage_data_reg[303]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_302_ ( .D(N2675), .CP(clk), 
        .Q(inner_first_stage_data_reg[302]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_301_ ( .D(N2674), .CP(clk), 
        .Q(inner_first_stage_data_reg[301]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_300_ ( .D(N2673), .CP(clk), 
        .Q(inner_first_stage_data_reg[300]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_299_ ( .D(N2672), .CP(clk), 
        .Q(inner_first_stage_data_reg[299]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_298_ ( .D(N2671), .CP(clk), 
        .Q(inner_first_stage_data_reg[298]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_297_ ( .D(N2670), .CP(clk), 
        .Q(inner_first_stage_data_reg[297]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_296_ ( .D(N2669), .CP(clk), 
        .Q(inner_first_stage_data_reg[296]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_295_ ( .D(N2668), .CP(clk), 
        .Q(inner_first_stage_data_reg[295]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_294_ ( .D(N2667), .CP(clk), 
        .Q(inner_first_stage_data_reg[294]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_293_ ( .D(N2666), .CP(clk), 
        .Q(inner_first_stage_data_reg[293]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_292_ ( .D(N2665), .CP(clk), 
        .Q(inner_first_stage_data_reg[292]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_291_ ( .D(N2664), .CP(clk), 
        .Q(inner_first_stage_data_reg[291]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_290_ ( .D(N2663), .CP(clk), 
        .Q(inner_first_stage_data_reg[290]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_289_ ( .D(N2662), .CP(clk), 
        .Q(inner_first_stage_data_reg[289]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_288_ ( .D(N2661), .CP(clk), 
        .Q(inner_first_stage_data_reg[288]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_9_ ( .D(N2660), .CP(clk), 
        .Q(inner_first_stage_valid_reg[9]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_351_ ( .D(N2908), .CP(clk), 
        .Q(inner_first_stage_data_reg[351]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_350_ ( .D(N2907), .CP(clk), 
        .Q(inner_first_stage_data_reg[350]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_349_ ( .D(N2906), .CP(clk), 
        .Q(inner_first_stage_data_reg[349]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_348_ ( .D(N2905), .CP(clk), 
        .Q(inner_first_stage_data_reg[348]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_347_ ( .D(N2904), .CP(clk), 
        .Q(inner_first_stage_data_reg[347]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_346_ ( .D(N2903), .CP(clk), 
        .Q(inner_first_stage_data_reg[346]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_345_ ( .D(N2902), .CP(clk), 
        .Q(inner_first_stage_data_reg[345]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_344_ ( .D(N2901), .CP(clk), 
        .Q(inner_first_stage_data_reg[344]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_343_ ( .D(N2900), .CP(clk), 
        .Q(inner_first_stage_data_reg[343]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_342_ ( .D(N2899), .CP(clk), 
        .Q(inner_first_stage_data_reg[342]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_341_ ( .D(N2898), .CP(clk), 
        .Q(inner_first_stage_data_reg[341]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_340_ ( .D(N2897), .CP(clk), 
        .Q(inner_first_stage_data_reg[340]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_339_ ( .D(N2896), .CP(clk), 
        .Q(inner_first_stage_data_reg[339]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_338_ ( .D(N2895), .CP(clk), 
        .Q(inner_first_stage_data_reg[338]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_337_ ( .D(N2894), .CP(clk), 
        .Q(inner_first_stage_data_reg[337]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_336_ ( .D(N2893), .CP(clk), 
        .Q(inner_first_stage_data_reg[336]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_335_ ( .D(N2892), .CP(clk), 
        .Q(inner_first_stage_data_reg[335]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_334_ ( .D(N2891), .CP(clk), 
        .Q(inner_first_stage_data_reg[334]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_333_ ( .D(N2890), .CP(clk), 
        .Q(inner_first_stage_data_reg[333]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_332_ ( .D(N2889), .CP(clk), 
        .Q(inner_first_stage_data_reg[332]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_331_ ( .D(N2888), .CP(clk), 
        .Q(inner_first_stage_data_reg[331]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_330_ ( .D(N2887), .CP(clk), 
        .Q(inner_first_stage_data_reg[330]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_329_ ( .D(N2886), .CP(clk), 
        .Q(inner_first_stage_data_reg[329]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_328_ ( .D(N2885), .CP(clk), 
        .Q(inner_first_stage_data_reg[328]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_327_ ( .D(N2884), .CP(clk), 
        .Q(inner_first_stage_data_reg[327]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_326_ ( .D(N2883), .CP(clk), 
        .Q(inner_first_stage_data_reg[326]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_325_ ( .D(N2882), .CP(clk), 
        .Q(inner_first_stage_data_reg[325]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_324_ ( .D(N2881), .CP(clk), 
        .Q(inner_first_stage_data_reg[324]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_323_ ( .D(N2880), .CP(clk), 
        .Q(inner_first_stage_data_reg[323]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_322_ ( .D(N2879), .CP(clk), 
        .Q(inner_first_stage_data_reg[322]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_321_ ( .D(N2878), .CP(clk), 
        .Q(inner_first_stage_data_reg[321]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_320_ ( .D(N2877), .CP(clk), 
        .Q(inner_first_stage_data_reg[320]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_10_ ( .D(N2876), .CP(clk), 
        .Q(inner_first_stage_valid_reg[10]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_383_ ( .D(N3124), .CP(clk), 
        .Q(inner_first_stage_data_reg[383]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_382_ ( .D(N3123), .CP(clk), 
        .Q(inner_first_stage_data_reg[382]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_381_ ( .D(N3122), .CP(clk), 
        .Q(inner_first_stage_data_reg[381]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_380_ ( .D(N3121), .CP(clk), 
        .Q(inner_first_stage_data_reg[380]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_379_ ( .D(N3120), .CP(clk), 
        .Q(inner_first_stage_data_reg[379]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_378_ ( .D(N3119), .CP(clk), 
        .Q(inner_first_stage_data_reg[378]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_377_ ( .D(N3118), .CP(clk), 
        .Q(inner_first_stage_data_reg[377]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_376_ ( .D(N3117), .CP(clk), 
        .Q(inner_first_stage_data_reg[376]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_375_ ( .D(N3116), .CP(clk), 
        .Q(inner_first_stage_data_reg[375]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_374_ ( .D(N3115), .CP(clk), 
        .Q(inner_first_stage_data_reg[374]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_373_ ( .D(N3114), .CP(clk), 
        .Q(inner_first_stage_data_reg[373]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_372_ ( .D(N3113), .CP(clk), 
        .Q(inner_first_stage_data_reg[372]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_371_ ( .D(N3112), .CP(clk), 
        .Q(inner_first_stage_data_reg[371]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_370_ ( .D(N3111), .CP(clk), 
        .Q(inner_first_stage_data_reg[370]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_369_ ( .D(N3110), .CP(clk), 
        .Q(inner_first_stage_data_reg[369]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_368_ ( .D(N3109), .CP(clk), 
        .Q(inner_first_stage_data_reg[368]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_367_ ( .D(N3108), .CP(clk), 
        .Q(inner_first_stage_data_reg[367]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_366_ ( .D(N3107), .CP(clk), 
        .Q(inner_first_stage_data_reg[366]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_365_ ( .D(N3106), .CP(clk), 
        .Q(inner_first_stage_data_reg[365]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_364_ ( .D(N3105), .CP(clk), 
        .Q(inner_first_stage_data_reg[364]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_363_ ( .D(N3104), .CP(clk), 
        .Q(inner_first_stage_data_reg[363]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_362_ ( .D(N3103), .CP(clk), 
        .Q(inner_first_stage_data_reg[362]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_361_ ( .D(N3102), .CP(clk), 
        .Q(inner_first_stage_data_reg[361]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_360_ ( .D(N3101), .CP(clk), 
        .Q(inner_first_stage_data_reg[360]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_359_ ( .D(N3100), .CP(clk), 
        .Q(inner_first_stage_data_reg[359]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_358_ ( .D(N3099), .CP(clk), 
        .Q(inner_first_stage_data_reg[358]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_357_ ( .D(N3098), .CP(clk), 
        .Q(inner_first_stage_data_reg[357]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_356_ ( .D(N3097), .CP(clk), 
        .Q(inner_first_stage_data_reg[356]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_355_ ( .D(N3096), .CP(clk), 
        .Q(inner_first_stage_data_reg[355]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_354_ ( .D(N3095), .CP(clk), 
        .Q(inner_first_stage_data_reg[354]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_353_ ( .D(N3094), .CP(clk), 
        .Q(inner_first_stage_data_reg[353]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_352_ ( .D(N3093), .CP(clk), 
        .Q(inner_first_stage_data_reg[352]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_11_ ( .D(N3092), .CP(clk), 
        .Q(inner_first_stage_valid_reg[11]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_415_ ( .D(N3340), .CP(clk), 
        .Q(inner_first_stage_data_reg[415]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_414_ ( .D(N3339), .CP(clk), 
        .Q(inner_first_stage_data_reg[414]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_413_ ( .D(N3338), .CP(clk), 
        .Q(inner_first_stage_data_reg[413]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_412_ ( .D(N3337), .CP(clk), 
        .Q(inner_first_stage_data_reg[412]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_411_ ( .D(N3336), .CP(clk), 
        .Q(inner_first_stage_data_reg[411]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_410_ ( .D(N3335), .CP(clk), 
        .Q(inner_first_stage_data_reg[410]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_409_ ( .D(N3334), .CP(clk), 
        .Q(inner_first_stage_data_reg[409]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_408_ ( .D(N3333), .CP(clk), 
        .Q(inner_first_stage_data_reg[408]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_407_ ( .D(N3332), .CP(clk), 
        .Q(inner_first_stage_data_reg[407]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_406_ ( .D(N3331), .CP(clk), 
        .Q(inner_first_stage_data_reg[406]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_405_ ( .D(N3330), .CP(clk), 
        .Q(inner_first_stage_data_reg[405]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_404_ ( .D(N3329), .CP(clk), 
        .Q(inner_first_stage_data_reg[404]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_403_ ( .D(N3328), .CP(clk), 
        .Q(inner_first_stage_data_reg[403]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_402_ ( .D(N3327), .CP(clk), 
        .Q(inner_first_stage_data_reg[402]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_401_ ( .D(N3326), .CP(clk), 
        .Q(inner_first_stage_data_reg[401]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_400_ ( .D(N3325), .CP(clk), 
        .Q(inner_first_stage_data_reg[400]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_399_ ( .D(N3324), .CP(clk), 
        .Q(inner_first_stage_data_reg[399]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_398_ ( .D(N3323), .CP(clk), 
        .Q(inner_first_stage_data_reg[398]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_397_ ( .D(N3322), .CP(clk), 
        .Q(inner_first_stage_data_reg[397]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_396_ ( .D(N3321), .CP(clk), 
        .Q(inner_first_stage_data_reg[396]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_395_ ( .D(N3320), .CP(clk), 
        .Q(inner_first_stage_data_reg[395]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_394_ ( .D(N3319), .CP(clk), 
        .Q(inner_first_stage_data_reg[394]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_393_ ( .D(N3318), .CP(clk), 
        .Q(inner_first_stage_data_reg[393]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_392_ ( .D(N3317), .CP(clk), 
        .Q(inner_first_stage_data_reg[392]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_391_ ( .D(N3316), .CP(clk), 
        .Q(inner_first_stage_data_reg[391]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_390_ ( .D(N3315), .CP(clk), 
        .Q(inner_first_stage_data_reg[390]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_389_ ( .D(N3314), .CP(clk), 
        .Q(inner_first_stage_data_reg[389]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_388_ ( .D(N3313), .CP(clk), 
        .Q(inner_first_stage_data_reg[388]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_387_ ( .D(N3312), .CP(clk), 
        .Q(inner_first_stage_data_reg[387]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_386_ ( .D(N3311), .CP(clk), 
        .Q(inner_first_stage_data_reg[386]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_385_ ( .D(N3310), .CP(clk), 
        .Q(inner_first_stage_data_reg[385]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_384_ ( .D(N3309), .CP(clk), 
        .Q(inner_first_stage_data_reg[384]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_12_ ( .D(N3308), .CP(clk), 
        .Q(inner_first_stage_valid_reg[12]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_447_ ( .D(N3556), .CP(clk), 
        .Q(inner_first_stage_data_reg[447]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_446_ ( .D(N3555), .CP(clk), 
        .Q(inner_first_stage_data_reg[446]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_445_ ( .D(N3554), .CP(clk), 
        .Q(inner_first_stage_data_reg[445]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_444_ ( .D(N3553), .CP(clk), 
        .Q(inner_first_stage_data_reg[444]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_443_ ( .D(N3552), .CP(clk), 
        .Q(inner_first_stage_data_reg[443]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_442_ ( .D(N3551), .CP(clk), 
        .Q(inner_first_stage_data_reg[442]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_441_ ( .D(N3550), .CP(clk), 
        .Q(inner_first_stage_data_reg[441]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_440_ ( .D(N3549), .CP(clk), 
        .Q(inner_first_stage_data_reg[440]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_439_ ( .D(N3548), .CP(clk), 
        .Q(inner_first_stage_data_reg[439]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_438_ ( .D(N3547), .CP(clk), 
        .Q(inner_first_stage_data_reg[438]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_437_ ( .D(N3546), .CP(clk), 
        .Q(inner_first_stage_data_reg[437]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_436_ ( .D(N3545), .CP(clk), 
        .Q(inner_first_stage_data_reg[436]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_435_ ( .D(N3544), .CP(clk), 
        .Q(inner_first_stage_data_reg[435]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_434_ ( .D(N3543), .CP(clk), 
        .Q(inner_first_stage_data_reg[434]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_433_ ( .D(N3542), .CP(clk), 
        .Q(inner_first_stage_data_reg[433]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_432_ ( .D(N3541), .CP(clk), 
        .Q(inner_first_stage_data_reg[432]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_431_ ( .D(N3540), .CP(clk), 
        .Q(inner_first_stage_data_reg[431]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_430_ ( .D(N3539), .CP(clk), 
        .Q(inner_first_stage_data_reg[430]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_429_ ( .D(N3538), .CP(clk), 
        .Q(inner_first_stage_data_reg[429]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_428_ ( .D(N3537), .CP(clk), 
        .Q(inner_first_stage_data_reg[428]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_427_ ( .D(N3536), .CP(clk), 
        .Q(inner_first_stage_data_reg[427]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_426_ ( .D(N3535), .CP(clk), 
        .Q(inner_first_stage_data_reg[426]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_425_ ( .D(N3534), .CP(clk), 
        .Q(inner_first_stage_data_reg[425]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_424_ ( .D(N3533), .CP(clk), 
        .Q(inner_first_stage_data_reg[424]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_423_ ( .D(N3532), .CP(clk), 
        .Q(inner_first_stage_data_reg[423]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_422_ ( .D(N3531), .CP(clk), 
        .Q(inner_first_stage_data_reg[422]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_421_ ( .D(N3530), .CP(clk), 
        .Q(inner_first_stage_data_reg[421]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_420_ ( .D(N3529), .CP(clk), 
        .Q(inner_first_stage_data_reg[420]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_419_ ( .D(N3528), .CP(clk), 
        .Q(inner_first_stage_data_reg[419]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_418_ ( .D(N3527), .CP(clk), 
        .Q(inner_first_stage_data_reg[418]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_417_ ( .D(N3526), .CP(clk), 
        .Q(inner_first_stage_data_reg[417]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_416_ ( .D(N3525), .CP(clk), 
        .Q(inner_first_stage_data_reg[416]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_13_ ( .D(N3524), .CP(clk), 
        .Q(inner_first_stage_valid_reg[13]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_479_ ( .D(N3772), .CP(clk), 
        .Q(inner_first_stage_data_reg[479]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_478_ ( .D(N3771), .CP(clk), 
        .Q(inner_first_stage_data_reg[478]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_477_ ( .D(N3770), .CP(clk), 
        .Q(inner_first_stage_data_reg[477]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_476_ ( .D(N3769), .CP(clk), 
        .Q(inner_first_stage_data_reg[476]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_475_ ( .D(N3768), .CP(clk), 
        .Q(inner_first_stage_data_reg[475]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_474_ ( .D(N3767), .CP(clk), 
        .Q(inner_first_stage_data_reg[474]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_473_ ( .D(N3766), .CP(clk), 
        .Q(inner_first_stage_data_reg[473]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_472_ ( .D(N3765), .CP(clk), 
        .Q(inner_first_stage_data_reg[472]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_471_ ( .D(N3764), .CP(clk), 
        .Q(inner_first_stage_data_reg[471]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_470_ ( .D(N3763), .CP(clk), 
        .Q(inner_first_stage_data_reg[470]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_469_ ( .D(N3762), .CP(clk), 
        .Q(inner_first_stage_data_reg[469]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_468_ ( .D(N3761), .CP(clk), 
        .Q(inner_first_stage_data_reg[468]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_467_ ( .D(N3760), .CP(clk), 
        .Q(inner_first_stage_data_reg[467]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_466_ ( .D(N3759), .CP(clk), 
        .Q(inner_first_stage_data_reg[466]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_465_ ( .D(N3758), .CP(clk), 
        .Q(inner_first_stage_data_reg[465]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_464_ ( .D(N3757), .CP(clk), 
        .Q(inner_first_stage_data_reg[464]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_463_ ( .D(N3756), .CP(clk), 
        .Q(inner_first_stage_data_reg[463]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_462_ ( .D(N3755), .CP(clk), 
        .Q(inner_first_stage_data_reg[462]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_461_ ( .D(N3754), .CP(clk), 
        .Q(inner_first_stage_data_reg[461]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_460_ ( .D(N3753), .CP(clk), 
        .Q(inner_first_stage_data_reg[460]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_459_ ( .D(N3752), .CP(clk), 
        .Q(inner_first_stage_data_reg[459]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_458_ ( .D(N3751), .CP(clk), 
        .Q(inner_first_stage_data_reg[458]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_457_ ( .D(N3750), .CP(clk), 
        .Q(inner_first_stage_data_reg[457]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_456_ ( .D(N3749), .CP(clk), 
        .Q(inner_first_stage_data_reg[456]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_455_ ( .D(N3748), .CP(clk), 
        .Q(inner_first_stage_data_reg[455]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_454_ ( .D(N3747), .CP(clk), 
        .Q(inner_first_stage_data_reg[454]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_453_ ( .D(N3746), .CP(clk), 
        .Q(inner_first_stage_data_reg[453]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_452_ ( .D(N3745), .CP(clk), 
        .Q(inner_first_stage_data_reg[452]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_451_ ( .D(N3744), .CP(clk), 
        .Q(inner_first_stage_data_reg[451]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_450_ ( .D(N3743), .CP(clk), 
        .Q(inner_first_stage_data_reg[450]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_449_ ( .D(N3742), .CP(clk), 
        .Q(inner_first_stage_data_reg[449]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_448_ ( .D(N3741), .CP(clk), 
        .Q(inner_first_stage_data_reg[448]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_14_ ( .D(N3740), .CP(clk), 
        .Q(inner_first_stage_valid_reg[14]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_511_ ( .D(N3988), .CP(clk), 
        .Q(inner_first_stage_data_reg[511]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_510_ ( .D(N3987), .CP(clk), 
        .Q(inner_first_stage_data_reg[510]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_509_ ( .D(N3986), .CP(clk), 
        .Q(inner_first_stage_data_reg[509]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_508_ ( .D(N3985), .CP(clk), 
        .Q(inner_first_stage_data_reg[508]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_507_ ( .D(N3984), .CP(clk), 
        .Q(inner_first_stage_data_reg[507]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_506_ ( .D(N3983), .CP(clk), 
        .Q(inner_first_stage_data_reg[506]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_505_ ( .D(N3982), .CP(clk), 
        .Q(inner_first_stage_data_reg[505]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_504_ ( .D(N3981), .CP(clk), 
        .Q(inner_first_stage_data_reg[504]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_503_ ( .D(N3980), .CP(clk), 
        .Q(inner_first_stage_data_reg[503]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_502_ ( .D(N3979), .CP(clk), 
        .Q(inner_first_stage_data_reg[502]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_501_ ( .D(N3978), .CP(clk), 
        .Q(inner_first_stage_data_reg[501]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_500_ ( .D(N3977), .CP(clk), 
        .Q(inner_first_stage_data_reg[500]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_499_ ( .D(N3976), .CP(clk), 
        .Q(inner_first_stage_data_reg[499]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_498_ ( .D(N3975), .CP(clk), 
        .Q(inner_first_stage_data_reg[498]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_497_ ( .D(N3974), .CP(clk), 
        .Q(inner_first_stage_data_reg[497]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_496_ ( .D(N3973), .CP(clk), 
        .Q(inner_first_stage_data_reg[496]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_495_ ( .D(N3972), .CP(clk), 
        .Q(inner_first_stage_data_reg[495]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_494_ ( .D(N3971), .CP(clk), 
        .Q(inner_first_stage_data_reg[494]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_493_ ( .D(N3970), .CP(clk), 
        .Q(inner_first_stage_data_reg[493]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_492_ ( .D(N3969), .CP(clk), 
        .Q(inner_first_stage_data_reg[492]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_491_ ( .D(N3968), .CP(clk), 
        .Q(inner_first_stage_data_reg[491]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_490_ ( .D(N3967), .CP(clk), 
        .Q(inner_first_stage_data_reg[490]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_489_ ( .D(N3966), .CP(clk), 
        .Q(inner_first_stage_data_reg[489]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_488_ ( .D(N3965), .CP(clk), 
        .Q(inner_first_stage_data_reg[488]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_487_ ( .D(N3964), .CP(clk), 
        .Q(inner_first_stage_data_reg[487]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_486_ ( .D(N3963), .CP(clk), 
        .Q(inner_first_stage_data_reg[486]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_485_ ( .D(N3962), .CP(clk), 
        .Q(inner_first_stage_data_reg[485]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_484_ ( .D(N3961), .CP(clk), 
        .Q(inner_first_stage_data_reg[484]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_483_ ( .D(N3960), .CP(clk), 
        .Q(inner_first_stage_data_reg[483]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_482_ ( .D(N3959), .CP(clk), 
        .Q(inner_first_stage_data_reg[482]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_481_ ( .D(N3958), .CP(clk), 
        .Q(inner_first_stage_data_reg[481]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_480_ ( .D(N3957), .CP(clk), 
        .Q(inner_first_stage_data_reg[480]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_15_ ( .D(N3956), .CP(clk), 
        .Q(inner_first_stage_valid_reg[15]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_543_ ( .D(N4350), .CP(clk), 
        .Q(inner_first_stage_data_reg[543]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_542_ ( .D(N4349), .CP(clk), 
        .Q(inner_first_stage_data_reg[542]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_541_ ( .D(N4348), .CP(clk), 
        .Q(inner_first_stage_data_reg[541]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_540_ ( .D(N4347), .CP(clk), 
        .Q(inner_first_stage_data_reg[540]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_539_ ( .D(N4346), .CP(clk), 
        .Q(inner_first_stage_data_reg[539]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_538_ ( .D(N4345), .CP(clk), 
        .Q(inner_first_stage_data_reg[538]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_537_ ( .D(N4344), .CP(clk), 
        .Q(inner_first_stage_data_reg[537]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_536_ ( .D(N4343), .CP(clk), 
        .Q(inner_first_stage_data_reg[536]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_535_ ( .D(N4342), .CP(clk), 
        .Q(inner_first_stage_data_reg[535]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_534_ ( .D(N4341), .CP(clk), 
        .Q(inner_first_stage_data_reg[534]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_533_ ( .D(N4340), .CP(clk), 
        .Q(inner_first_stage_data_reg[533]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_532_ ( .D(N4339), .CP(clk), 
        .Q(inner_first_stage_data_reg[532]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_531_ ( .D(N4338), .CP(clk), 
        .Q(inner_first_stage_data_reg[531]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_530_ ( .D(N4337), .CP(clk), 
        .Q(inner_first_stage_data_reg[530]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_529_ ( .D(N4336), .CP(clk), 
        .Q(inner_first_stage_data_reg[529]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_528_ ( .D(N4335), .CP(clk), 
        .Q(inner_first_stage_data_reg[528]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_527_ ( .D(N4334), .CP(clk), 
        .Q(inner_first_stage_data_reg[527]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_526_ ( .D(N4333), .CP(clk), 
        .Q(inner_first_stage_data_reg[526]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_525_ ( .D(N4332), .CP(clk), 
        .Q(inner_first_stage_data_reg[525]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_524_ ( .D(N4331), .CP(clk), 
        .Q(inner_first_stage_data_reg[524]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_523_ ( .D(N4330), .CP(clk), 
        .Q(inner_first_stage_data_reg[523]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_522_ ( .D(N4329), .CP(clk), 
        .Q(inner_first_stage_data_reg[522]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_521_ ( .D(N4328), .CP(clk), 
        .Q(inner_first_stage_data_reg[521]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_520_ ( .D(N4327), .CP(clk), 
        .Q(inner_first_stage_data_reg[520]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_519_ ( .D(N4326), .CP(clk), 
        .Q(inner_first_stage_data_reg[519]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_518_ ( .D(N4325), .CP(clk), 
        .Q(inner_first_stage_data_reg[518]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_517_ ( .D(N4324), .CP(clk), 
        .Q(inner_first_stage_data_reg[517]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_516_ ( .D(N4323), .CP(clk), 
        .Q(inner_first_stage_data_reg[516]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_515_ ( .D(N4322), .CP(clk), 
        .Q(inner_first_stage_data_reg[515]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_514_ ( .D(N4321), .CP(clk), 
        .Q(inner_first_stage_data_reg[514]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_513_ ( .D(N4320), .CP(clk), 
        .Q(inner_first_stage_data_reg[513]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_512_ ( .D(N4319), .CP(clk), 
        .Q(inner_first_stage_data_reg[512]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_16_ ( .D(N4318), .CP(clk), 
        .Q(inner_first_stage_valid_reg[16]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_575_ ( .D(N4566), .CP(clk), 
        .Q(inner_first_stage_data_reg[575]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_574_ ( .D(N4565), .CP(clk), 
        .Q(inner_first_stage_data_reg[574]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_573_ ( .D(N4564), .CP(clk), 
        .Q(inner_first_stage_data_reg[573]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_572_ ( .D(N4563), .CP(clk), 
        .Q(inner_first_stage_data_reg[572]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_571_ ( .D(N4562), .CP(clk), 
        .Q(inner_first_stage_data_reg[571]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_570_ ( .D(N4561), .CP(clk), 
        .Q(inner_first_stage_data_reg[570]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_569_ ( .D(N4560), .CP(clk), 
        .Q(inner_first_stage_data_reg[569]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_568_ ( .D(N4559), .CP(clk), 
        .Q(inner_first_stage_data_reg[568]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_567_ ( .D(N4558), .CP(clk), 
        .Q(inner_first_stage_data_reg[567]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_566_ ( .D(N4557), .CP(clk), 
        .Q(inner_first_stage_data_reg[566]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_565_ ( .D(N4556), .CP(clk), 
        .Q(inner_first_stage_data_reg[565]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_564_ ( .D(N4555), .CP(clk), 
        .Q(inner_first_stage_data_reg[564]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_563_ ( .D(N4554), .CP(clk), 
        .Q(inner_first_stage_data_reg[563]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_562_ ( .D(N4553), .CP(clk), 
        .Q(inner_first_stage_data_reg[562]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_561_ ( .D(N4552), .CP(clk), 
        .Q(inner_first_stage_data_reg[561]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_560_ ( .D(N4551), .CP(clk), 
        .Q(inner_first_stage_data_reg[560]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_559_ ( .D(N4550), .CP(clk), 
        .Q(inner_first_stage_data_reg[559]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_558_ ( .D(N4549), .CP(clk), 
        .Q(inner_first_stage_data_reg[558]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_557_ ( .D(N4548), .CP(clk), 
        .Q(inner_first_stage_data_reg[557]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_556_ ( .D(N4547), .CP(clk), 
        .Q(inner_first_stage_data_reg[556]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_555_ ( .D(N4546), .CP(clk), 
        .Q(inner_first_stage_data_reg[555]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_554_ ( .D(N4545), .CP(clk), 
        .Q(inner_first_stage_data_reg[554]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_553_ ( .D(N4544), .CP(clk), 
        .Q(inner_first_stage_data_reg[553]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_552_ ( .D(N4543), .CP(clk), 
        .Q(inner_first_stage_data_reg[552]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_551_ ( .D(N4542), .CP(clk), 
        .Q(inner_first_stage_data_reg[551]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_550_ ( .D(N4541), .CP(clk), 
        .Q(inner_first_stage_data_reg[550]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_549_ ( .D(N4540), .CP(clk), 
        .Q(inner_first_stage_data_reg[549]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_548_ ( .D(N4539), .CP(clk), 
        .Q(inner_first_stage_data_reg[548]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_547_ ( .D(N4538), .CP(clk), 
        .Q(inner_first_stage_data_reg[547]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_546_ ( .D(N4537), .CP(clk), 
        .Q(inner_first_stage_data_reg[546]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_545_ ( .D(N4536), .CP(clk), 
        .Q(inner_first_stage_data_reg[545]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_544_ ( .D(N4535), .CP(clk), 
        .Q(inner_first_stage_data_reg[544]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_17_ ( .D(N4534), .CP(clk), 
        .Q(inner_first_stage_valid_reg[17]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_607_ ( .D(N4782), .CP(clk), 
        .Q(inner_first_stage_data_reg[607]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_606_ ( .D(N4781), .CP(clk), 
        .Q(inner_first_stage_data_reg[606]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_605_ ( .D(N4780), .CP(clk), 
        .Q(inner_first_stage_data_reg[605]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_604_ ( .D(N4779), .CP(clk), 
        .Q(inner_first_stage_data_reg[604]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_603_ ( .D(N4778), .CP(clk), 
        .Q(inner_first_stage_data_reg[603]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_602_ ( .D(N4777), .CP(clk), 
        .Q(inner_first_stage_data_reg[602]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_601_ ( .D(N4776), .CP(clk), 
        .Q(inner_first_stage_data_reg[601]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_600_ ( .D(N4775), .CP(clk), 
        .Q(inner_first_stage_data_reg[600]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_599_ ( .D(N4774), .CP(clk), 
        .Q(inner_first_stage_data_reg[599]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_598_ ( .D(N4773), .CP(clk), 
        .Q(inner_first_stage_data_reg[598]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_597_ ( .D(N4772), .CP(clk), 
        .Q(inner_first_stage_data_reg[597]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_596_ ( .D(N4771), .CP(clk), 
        .Q(inner_first_stage_data_reg[596]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_595_ ( .D(N4770), .CP(clk), 
        .Q(inner_first_stage_data_reg[595]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_594_ ( .D(N4769), .CP(clk), 
        .Q(inner_first_stage_data_reg[594]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_593_ ( .D(N4768), .CP(clk), 
        .Q(inner_first_stage_data_reg[593]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_592_ ( .D(N4767), .CP(clk), 
        .Q(inner_first_stage_data_reg[592]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_591_ ( .D(N4766), .CP(clk), 
        .Q(inner_first_stage_data_reg[591]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_590_ ( .D(N4765), .CP(clk), 
        .Q(inner_first_stage_data_reg[590]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_589_ ( .D(N4764), .CP(clk), 
        .Q(inner_first_stage_data_reg[589]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_588_ ( .D(N4763), .CP(clk), 
        .Q(inner_first_stage_data_reg[588]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_587_ ( .D(N4762), .CP(clk), 
        .Q(inner_first_stage_data_reg[587]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_586_ ( .D(N4761), .CP(clk), 
        .Q(inner_first_stage_data_reg[586]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_585_ ( .D(N4760), .CP(clk), 
        .Q(inner_first_stage_data_reg[585]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_584_ ( .D(N4759), .CP(clk), 
        .Q(inner_first_stage_data_reg[584]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_583_ ( .D(N4758), .CP(clk), 
        .Q(inner_first_stage_data_reg[583]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_582_ ( .D(N4757), .CP(clk), 
        .Q(inner_first_stage_data_reg[582]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_581_ ( .D(N4756), .CP(clk), 
        .Q(inner_first_stage_data_reg[581]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_580_ ( .D(N4755), .CP(clk), 
        .Q(inner_first_stage_data_reg[580]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_579_ ( .D(N4754), .CP(clk), 
        .Q(inner_first_stage_data_reg[579]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_578_ ( .D(N4753), .CP(clk), 
        .Q(inner_first_stage_data_reg[578]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_577_ ( .D(N4752), .CP(clk), 
        .Q(inner_first_stage_data_reg[577]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_576_ ( .D(N4751), .CP(clk), 
        .Q(inner_first_stage_data_reg[576]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_639_ ( .D(N4998), .CP(clk), 
        .Q(inner_first_stage_data_reg[639]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_638_ ( .D(N4997), .CP(clk), 
        .Q(inner_first_stage_data_reg[638]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_637_ ( .D(N4996), .CP(clk), 
        .Q(inner_first_stage_data_reg[637]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_636_ ( .D(N4995), .CP(clk), 
        .Q(inner_first_stage_data_reg[636]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_635_ ( .D(N4994), .CP(clk), 
        .Q(inner_first_stage_data_reg[635]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_634_ ( .D(N4993), .CP(clk), 
        .Q(inner_first_stage_data_reg[634]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_633_ ( .D(N4992), .CP(clk), 
        .Q(inner_first_stage_data_reg[633]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_632_ ( .D(N4991), .CP(clk), 
        .Q(inner_first_stage_data_reg[632]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_631_ ( .D(N4990), .CP(clk), 
        .Q(inner_first_stage_data_reg[631]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_630_ ( .D(N4989), .CP(clk), 
        .Q(inner_first_stage_data_reg[630]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_629_ ( .D(N4988), .CP(clk), 
        .Q(inner_first_stage_data_reg[629]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_628_ ( .D(N4987), .CP(clk), 
        .Q(inner_first_stage_data_reg[628]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_627_ ( .D(N4986), .CP(clk), 
        .Q(inner_first_stage_data_reg[627]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_626_ ( .D(N4985), .CP(clk), 
        .Q(inner_first_stage_data_reg[626]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_625_ ( .D(N4984), .CP(clk), 
        .Q(inner_first_stage_data_reg[625]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_624_ ( .D(N4983), .CP(clk), 
        .Q(inner_first_stage_data_reg[624]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_623_ ( .D(N4982), .CP(clk), 
        .Q(inner_first_stage_data_reg[623]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_622_ ( .D(N4981), .CP(clk), 
        .Q(inner_first_stage_data_reg[622]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_621_ ( .D(N4980), .CP(clk), 
        .Q(inner_first_stage_data_reg[621]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_620_ ( .D(N4979), .CP(clk), 
        .Q(inner_first_stage_data_reg[620]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_619_ ( .D(N4978), .CP(clk), 
        .Q(inner_first_stage_data_reg[619]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_618_ ( .D(N4977), .CP(clk), 
        .Q(inner_first_stage_data_reg[618]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_617_ ( .D(N4976), .CP(clk), 
        .Q(inner_first_stage_data_reg[617]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_616_ ( .D(N4975), .CP(clk), 
        .Q(inner_first_stage_data_reg[616]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_615_ ( .D(N4974), .CP(clk), 
        .Q(inner_first_stage_data_reg[615]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_614_ ( .D(N4973), .CP(clk), 
        .Q(inner_first_stage_data_reg[614]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_613_ ( .D(N4972), .CP(clk), 
        .Q(inner_first_stage_data_reg[613]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_612_ ( .D(N4971), .CP(clk), 
        .Q(inner_first_stage_data_reg[612]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_611_ ( .D(N4970), .CP(clk), 
        .Q(inner_first_stage_data_reg[611]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_610_ ( .D(N4969), .CP(clk), 
        .Q(inner_first_stage_data_reg[610]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_609_ ( .D(N4968), .CP(clk), 
        .Q(inner_first_stage_data_reg[609]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_608_ ( .D(N4967), .CP(clk), 
        .Q(inner_first_stage_data_reg[608]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_19_ ( .D(N4966), .CP(clk), 
        .Q(inner_first_stage_valid_reg[19]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_671_ ( .D(N5214), .CP(clk), 
        .Q(inner_first_stage_data_reg[671]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_670_ ( .D(N5213), .CP(clk), 
        .Q(inner_first_stage_data_reg[670]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_669_ ( .D(N5212), .CP(clk), 
        .Q(inner_first_stage_data_reg[669]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_668_ ( .D(N5211), .CP(clk), 
        .Q(inner_first_stage_data_reg[668]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_667_ ( .D(N5210), .CP(clk), 
        .Q(inner_first_stage_data_reg[667]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_666_ ( .D(N5209), .CP(clk), 
        .Q(inner_first_stage_data_reg[666]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_665_ ( .D(N5208), .CP(clk), 
        .Q(inner_first_stage_data_reg[665]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_664_ ( .D(N5207), .CP(clk), 
        .Q(inner_first_stage_data_reg[664]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_663_ ( .D(N5206), .CP(clk), 
        .Q(inner_first_stage_data_reg[663]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_662_ ( .D(N5205), .CP(clk), 
        .Q(inner_first_stage_data_reg[662]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_661_ ( .D(N5204), .CP(clk), 
        .Q(inner_first_stage_data_reg[661]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_660_ ( .D(N5203), .CP(clk), 
        .Q(inner_first_stage_data_reg[660]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_659_ ( .D(N5202), .CP(clk), 
        .Q(inner_first_stage_data_reg[659]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_658_ ( .D(N5201), .CP(clk), 
        .Q(inner_first_stage_data_reg[658]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_657_ ( .D(N5200), .CP(clk), 
        .Q(inner_first_stage_data_reg[657]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_656_ ( .D(N5199), .CP(clk), 
        .Q(inner_first_stage_data_reg[656]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_655_ ( .D(N5198), .CP(clk), 
        .Q(inner_first_stage_data_reg[655]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_654_ ( .D(N5197), .CP(clk), 
        .Q(inner_first_stage_data_reg[654]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_653_ ( .D(N5196), .CP(clk), 
        .Q(inner_first_stage_data_reg[653]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_652_ ( .D(N5195), .CP(clk), 
        .Q(inner_first_stage_data_reg[652]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_651_ ( .D(N5194), .CP(clk), 
        .Q(inner_first_stage_data_reg[651]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_650_ ( .D(N5193), .CP(clk), 
        .Q(inner_first_stage_data_reg[650]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_649_ ( .D(N5192), .CP(clk), 
        .Q(inner_first_stage_data_reg[649]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_648_ ( .D(N5191), .CP(clk), 
        .Q(inner_first_stage_data_reg[648]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_647_ ( .D(N5190), .CP(clk), 
        .Q(inner_first_stage_data_reg[647]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_646_ ( .D(N5189), .CP(clk), 
        .Q(inner_first_stage_data_reg[646]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_645_ ( .D(N5188), .CP(clk), 
        .Q(inner_first_stage_data_reg[645]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_644_ ( .D(N5187), .CP(clk), 
        .Q(inner_first_stage_data_reg[644]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_643_ ( .D(N5186), .CP(clk), 
        .Q(inner_first_stage_data_reg[643]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_642_ ( .D(N5185), .CP(clk), 
        .Q(inner_first_stage_data_reg[642]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_641_ ( .D(N5184), .CP(clk), 
        .Q(inner_first_stage_data_reg[641]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_640_ ( .D(N5183), .CP(clk), 
        .Q(inner_first_stage_data_reg[640]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_20_ ( .D(N5182), .CP(clk), 
        .Q(inner_first_stage_valid_reg[20]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_703_ ( .D(N5430), .CP(clk), 
        .Q(inner_first_stage_data_reg[703]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_702_ ( .D(N5429), .CP(clk), 
        .Q(inner_first_stage_data_reg[702]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_701_ ( .D(N5428), .CP(clk), 
        .Q(inner_first_stage_data_reg[701]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_700_ ( .D(N5427), .CP(clk), 
        .Q(inner_first_stage_data_reg[700]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_699_ ( .D(N5426), .CP(clk), 
        .Q(inner_first_stage_data_reg[699]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_698_ ( .D(N5425), .CP(clk), 
        .Q(inner_first_stage_data_reg[698]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_697_ ( .D(N5424), .CP(clk), 
        .Q(inner_first_stage_data_reg[697]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_696_ ( .D(N5423), .CP(clk), 
        .Q(inner_first_stage_data_reg[696]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_695_ ( .D(N5422), .CP(clk), 
        .Q(inner_first_stage_data_reg[695]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_694_ ( .D(N5421), .CP(clk), 
        .Q(inner_first_stage_data_reg[694]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_693_ ( .D(N5420), .CP(clk), 
        .Q(inner_first_stage_data_reg[693]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_692_ ( .D(N5419), .CP(clk), 
        .Q(inner_first_stage_data_reg[692]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_691_ ( .D(N5418), .CP(clk), 
        .Q(inner_first_stage_data_reg[691]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_690_ ( .D(N5417), .CP(clk), 
        .Q(inner_first_stage_data_reg[690]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_689_ ( .D(N5416), .CP(clk), 
        .Q(inner_first_stage_data_reg[689]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_688_ ( .D(N5415), .CP(clk), 
        .Q(inner_first_stage_data_reg[688]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_687_ ( .D(N5414), .CP(clk), 
        .Q(inner_first_stage_data_reg[687]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_686_ ( .D(N5413), .CP(clk), 
        .Q(inner_first_stage_data_reg[686]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_685_ ( .D(N5412), .CP(clk), 
        .Q(inner_first_stage_data_reg[685]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_684_ ( .D(N5411), .CP(clk), 
        .Q(inner_first_stage_data_reg[684]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_683_ ( .D(N5410), .CP(clk), 
        .Q(inner_first_stage_data_reg[683]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_682_ ( .D(N5409), .CP(clk), 
        .Q(inner_first_stage_data_reg[682]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_681_ ( .D(N5408), .CP(clk), 
        .Q(inner_first_stage_data_reg[681]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_680_ ( .D(N5407), .CP(clk), 
        .Q(inner_first_stage_data_reg[680]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_679_ ( .D(N5406), .CP(clk), 
        .Q(inner_first_stage_data_reg[679]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_678_ ( .D(N5405), .CP(clk), 
        .Q(inner_first_stage_data_reg[678]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_677_ ( .D(N5404), .CP(clk), 
        .Q(inner_first_stage_data_reg[677]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_676_ ( .D(N5403), .CP(clk), 
        .Q(inner_first_stage_data_reg[676]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_675_ ( .D(N5402), .CP(clk), 
        .Q(inner_first_stage_data_reg[675]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_674_ ( .D(N5401), .CP(clk), 
        .Q(inner_first_stage_data_reg[674]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_673_ ( .D(N5400), .CP(clk), 
        .Q(inner_first_stage_data_reg[673]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_672_ ( .D(N5399), .CP(clk), 
        .Q(inner_first_stage_data_reg[672]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_21_ ( .D(N5398), .CP(clk), 
        .Q(inner_first_stage_valid_reg[21]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_735_ ( .D(N5646), .CP(clk), 
        .Q(inner_first_stage_data_reg[735]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_734_ ( .D(N5645), .CP(clk), 
        .Q(inner_first_stage_data_reg[734]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_733_ ( .D(N5644), .CP(clk), 
        .Q(inner_first_stage_data_reg[733]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_732_ ( .D(N5643), .CP(clk), 
        .Q(inner_first_stage_data_reg[732]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_731_ ( .D(N5642), .CP(clk), 
        .Q(inner_first_stage_data_reg[731]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_730_ ( .D(N5641), .CP(clk), 
        .Q(inner_first_stage_data_reg[730]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_729_ ( .D(N5640), .CP(clk), 
        .Q(inner_first_stage_data_reg[729]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_728_ ( .D(N5639), .CP(clk), 
        .Q(inner_first_stage_data_reg[728]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_727_ ( .D(N5638), .CP(clk), 
        .Q(inner_first_stage_data_reg[727]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_726_ ( .D(N5637), .CP(clk), 
        .Q(inner_first_stage_data_reg[726]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_725_ ( .D(N5636), .CP(clk), 
        .Q(inner_first_stage_data_reg[725]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_724_ ( .D(N5635), .CP(clk), 
        .Q(inner_first_stage_data_reg[724]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_723_ ( .D(N5634), .CP(clk), 
        .Q(inner_first_stage_data_reg[723]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_722_ ( .D(N5633), .CP(clk), 
        .Q(inner_first_stage_data_reg[722]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_721_ ( .D(N5632), .CP(clk), 
        .Q(inner_first_stage_data_reg[721]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_720_ ( .D(N5631), .CP(clk), 
        .Q(inner_first_stage_data_reg[720]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_719_ ( .D(N5630), .CP(clk), 
        .Q(inner_first_stage_data_reg[719]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_718_ ( .D(N5629), .CP(clk), 
        .Q(inner_first_stage_data_reg[718]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_717_ ( .D(N5628), .CP(clk), 
        .Q(inner_first_stage_data_reg[717]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_716_ ( .D(N5627), .CP(clk), 
        .Q(inner_first_stage_data_reg[716]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_715_ ( .D(N5626), .CP(clk), 
        .Q(inner_first_stage_data_reg[715]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_714_ ( .D(N5625), .CP(clk), 
        .Q(inner_first_stage_data_reg[714]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_713_ ( .D(N5624), .CP(clk), 
        .Q(inner_first_stage_data_reg[713]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_712_ ( .D(N5623), .CP(clk), 
        .Q(inner_first_stage_data_reg[712]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_711_ ( .D(N5622), .CP(clk), 
        .Q(inner_first_stage_data_reg[711]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_710_ ( .D(N5621), .CP(clk), 
        .Q(inner_first_stage_data_reg[710]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_709_ ( .D(N5620), .CP(clk), 
        .Q(inner_first_stage_data_reg[709]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_708_ ( .D(N5619), .CP(clk), 
        .Q(inner_first_stage_data_reg[708]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_707_ ( .D(N5618), .CP(clk), 
        .Q(inner_first_stage_data_reg[707]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_706_ ( .D(N5617), .CP(clk), 
        .Q(inner_first_stage_data_reg[706]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_705_ ( .D(N5616), .CP(clk), 
        .Q(inner_first_stage_data_reg[705]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_704_ ( .D(N5615), .CP(clk), 
        .Q(inner_first_stage_data_reg[704]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_22_ ( .D(N5614), .CP(clk), 
        .Q(inner_first_stage_valid_reg[22]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_767_ ( .D(N5862), .CP(clk), 
        .Q(inner_first_stage_data_reg[767]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_766_ ( .D(N5861), .CP(clk), 
        .Q(inner_first_stage_data_reg[766]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_765_ ( .D(N5860), .CP(clk), 
        .Q(inner_first_stage_data_reg[765]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_764_ ( .D(N5859), .CP(clk), 
        .Q(inner_first_stage_data_reg[764]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_763_ ( .D(N5858), .CP(clk), 
        .Q(inner_first_stage_data_reg[763]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_762_ ( .D(N5857), .CP(clk), 
        .Q(inner_first_stage_data_reg[762]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_761_ ( .D(N5856), .CP(clk), 
        .Q(inner_first_stage_data_reg[761]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_760_ ( .D(N5855), .CP(clk), 
        .Q(inner_first_stage_data_reg[760]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_759_ ( .D(N5854), .CP(clk), 
        .Q(inner_first_stage_data_reg[759]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_758_ ( .D(N5853), .CP(clk), 
        .Q(inner_first_stage_data_reg[758]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_757_ ( .D(N5852), .CP(clk), 
        .Q(inner_first_stage_data_reg[757]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_756_ ( .D(N5851), .CP(clk), 
        .Q(inner_first_stage_data_reg[756]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_755_ ( .D(N5850), .CP(clk), 
        .Q(inner_first_stage_data_reg[755]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_754_ ( .D(N5849), .CP(clk), 
        .Q(inner_first_stage_data_reg[754]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_753_ ( .D(N5848), .CP(clk), 
        .Q(inner_first_stage_data_reg[753]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_752_ ( .D(N5847), .CP(clk), 
        .Q(inner_first_stage_data_reg[752]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_751_ ( .D(N5846), .CP(clk), 
        .Q(inner_first_stage_data_reg[751]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_750_ ( .D(N5845), .CP(clk), 
        .Q(inner_first_stage_data_reg[750]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_749_ ( .D(N5844), .CP(clk), 
        .Q(inner_first_stage_data_reg[749]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_748_ ( .D(N5843), .CP(clk), 
        .Q(inner_first_stage_data_reg[748]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_747_ ( .D(N5842), .CP(clk), 
        .Q(inner_first_stage_data_reg[747]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_746_ ( .D(N5841), .CP(clk), 
        .Q(inner_first_stage_data_reg[746]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_745_ ( .D(N5840), .CP(clk), 
        .Q(inner_first_stage_data_reg[745]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_744_ ( .D(N5839), .CP(clk), 
        .Q(inner_first_stage_data_reg[744]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_743_ ( .D(N5838), .CP(clk), 
        .Q(inner_first_stage_data_reg[743]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_742_ ( .D(N5837), .CP(clk), 
        .Q(inner_first_stage_data_reg[742]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_741_ ( .D(N5836), .CP(clk), 
        .Q(inner_first_stage_data_reg[741]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_740_ ( .D(N5835), .CP(clk), 
        .Q(inner_first_stage_data_reg[740]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_739_ ( .D(N5834), .CP(clk), 
        .Q(inner_first_stage_data_reg[739]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_738_ ( .D(N5833), .CP(clk), 
        .Q(inner_first_stage_data_reg[738]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_737_ ( .D(N5832), .CP(clk), 
        .Q(inner_first_stage_data_reg[737]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_736_ ( .D(N5831), .CP(clk), 
        .Q(inner_first_stage_data_reg[736]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_23_ ( .D(N5830), .CP(clk), 
        .Q(inner_first_stage_valid_reg[23]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_799_ ( .D(N6224), .CP(clk), 
        .Q(inner_first_stage_data_reg[799]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_798_ ( .D(N6223), .CP(clk), 
        .Q(inner_first_stage_data_reg[798]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_797_ ( .D(N6222), .CP(clk), 
        .Q(inner_first_stage_data_reg[797]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_796_ ( .D(N6221), .CP(clk), 
        .Q(inner_first_stage_data_reg[796]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_795_ ( .D(N6220), .CP(clk), 
        .Q(inner_first_stage_data_reg[795]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_794_ ( .D(N6219), .CP(clk), 
        .Q(inner_first_stage_data_reg[794]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_793_ ( .D(N6218), .CP(clk), 
        .Q(inner_first_stage_data_reg[793]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_792_ ( .D(N6217), .CP(clk), 
        .Q(inner_first_stage_data_reg[792]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_791_ ( .D(N6216), .CP(clk), 
        .Q(inner_first_stage_data_reg[791]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_790_ ( .D(N6215), .CP(clk), 
        .Q(inner_first_stage_data_reg[790]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_789_ ( .D(N6214), .CP(clk), 
        .Q(inner_first_stage_data_reg[789]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_788_ ( .D(N6213), .CP(clk), 
        .Q(inner_first_stage_data_reg[788]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_787_ ( .D(N6212), .CP(clk), 
        .Q(inner_first_stage_data_reg[787]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_786_ ( .D(N6211), .CP(clk), 
        .Q(inner_first_stage_data_reg[786]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_785_ ( .D(N6210), .CP(clk), 
        .Q(inner_first_stage_data_reg[785]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_784_ ( .D(N6209), .CP(clk), 
        .Q(inner_first_stage_data_reg[784]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_783_ ( .D(N6208), .CP(clk), 
        .Q(inner_first_stage_data_reg[783]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_782_ ( .D(N6207), .CP(clk), 
        .Q(inner_first_stage_data_reg[782]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_781_ ( .D(N6206), .CP(clk), 
        .Q(inner_first_stage_data_reg[781]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_780_ ( .D(N6205), .CP(clk), 
        .Q(inner_first_stage_data_reg[780]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_779_ ( .D(N6204), .CP(clk), 
        .Q(inner_first_stage_data_reg[779]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_778_ ( .D(N6203), .CP(clk), 
        .Q(inner_first_stage_data_reg[778]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_777_ ( .D(N6202), .CP(clk), 
        .Q(inner_first_stage_data_reg[777]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_776_ ( .D(N6201), .CP(clk), 
        .Q(inner_first_stage_data_reg[776]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_775_ ( .D(N6200), .CP(clk), 
        .Q(inner_first_stage_data_reg[775]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_774_ ( .D(N6199), .CP(clk), 
        .Q(inner_first_stage_data_reg[774]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_773_ ( .D(N6198), .CP(clk), 
        .Q(inner_first_stage_data_reg[773]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_772_ ( .D(N6197), .CP(clk), 
        .Q(inner_first_stage_data_reg[772]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_771_ ( .D(N6196), .CP(clk), 
        .Q(inner_first_stage_data_reg[771]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_770_ ( .D(N6195), .CP(clk), 
        .Q(inner_first_stage_data_reg[770]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_769_ ( .D(N6194), .CP(clk), 
        .Q(inner_first_stage_data_reg[769]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_768_ ( .D(N6193), .CP(clk), 
        .Q(inner_first_stage_data_reg[768]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_24_ ( .D(N6192), .CP(clk), 
        .Q(inner_first_stage_valid_reg[24]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_831_ ( .D(N6440), .CP(clk), 
        .Q(inner_first_stage_data_reg[831]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_830_ ( .D(N6439), .CP(clk), 
        .Q(inner_first_stage_data_reg[830]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_829_ ( .D(N6438), .CP(clk), 
        .Q(inner_first_stage_data_reg[829]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_828_ ( .D(N6437), .CP(clk), 
        .Q(inner_first_stage_data_reg[828]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_827_ ( .D(N6436), .CP(clk), 
        .Q(inner_first_stage_data_reg[827]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_826_ ( .D(N6435), .CP(clk), 
        .Q(inner_first_stage_data_reg[826]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_825_ ( .D(N6434), .CP(clk), 
        .Q(inner_first_stage_data_reg[825]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_824_ ( .D(N6433), .CP(clk), 
        .Q(inner_first_stage_data_reg[824]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_823_ ( .D(N6432), .CP(clk), 
        .Q(inner_first_stage_data_reg[823]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_822_ ( .D(N6431), .CP(clk), 
        .Q(inner_first_stage_data_reg[822]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_821_ ( .D(N6430), .CP(clk), 
        .Q(inner_first_stage_data_reg[821]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_820_ ( .D(N6429), .CP(clk), 
        .Q(inner_first_stage_data_reg[820]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_819_ ( .D(N6428), .CP(clk), 
        .Q(inner_first_stage_data_reg[819]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_818_ ( .D(N6427), .CP(clk), 
        .Q(inner_first_stage_data_reg[818]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_817_ ( .D(N6426), .CP(clk), 
        .Q(inner_first_stage_data_reg[817]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_816_ ( .D(N6425), .CP(clk), 
        .Q(inner_first_stage_data_reg[816]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_815_ ( .D(N6424), .CP(clk), 
        .Q(inner_first_stage_data_reg[815]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_814_ ( .D(N6423), .CP(clk), 
        .Q(inner_first_stage_data_reg[814]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_813_ ( .D(N6422), .CP(clk), 
        .Q(inner_first_stage_data_reg[813]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_812_ ( .D(N6421), .CP(clk), 
        .Q(inner_first_stage_data_reg[812]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_811_ ( .D(N6420), .CP(clk), 
        .Q(inner_first_stage_data_reg[811]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_810_ ( .D(N6419), .CP(clk), 
        .Q(inner_first_stage_data_reg[810]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_809_ ( .D(N6418), .CP(clk), 
        .Q(inner_first_stage_data_reg[809]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_808_ ( .D(N6417), .CP(clk), 
        .Q(inner_first_stage_data_reg[808]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_807_ ( .D(N6416), .CP(clk), 
        .Q(inner_first_stage_data_reg[807]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_806_ ( .D(N6415), .CP(clk), 
        .Q(inner_first_stage_data_reg[806]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_805_ ( .D(N6414), .CP(clk), 
        .Q(inner_first_stage_data_reg[805]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_804_ ( .D(N6413), .CP(clk), 
        .Q(inner_first_stage_data_reg[804]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_803_ ( .D(N6412), .CP(clk), 
        .Q(inner_first_stage_data_reg[803]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_802_ ( .D(N6411), .CP(clk), 
        .Q(inner_first_stage_data_reg[802]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_801_ ( .D(N6410), .CP(clk), 
        .Q(inner_first_stage_data_reg[801]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_800_ ( .D(N6409), .CP(clk), 
        .Q(inner_first_stage_data_reg[800]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_25_ ( .D(N6408), .CP(clk), 
        .Q(inner_first_stage_valid_reg[25]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_863_ ( .D(N6656), .CP(clk), 
        .Q(inner_first_stage_data_reg[863]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_862_ ( .D(N6655), .CP(clk), 
        .Q(inner_first_stage_data_reg[862]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_861_ ( .D(N6654), .CP(clk), 
        .Q(inner_first_stage_data_reg[861]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_860_ ( .D(N6653), .CP(clk), 
        .Q(inner_first_stage_data_reg[860]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_859_ ( .D(N6652), .CP(clk), 
        .Q(inner_first_stage_data_reg[859]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_858_ ( .D(N6651), .CP(clk), 
        .Q(inner_first_stage_data_reg[858]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_857_ ( .D(N6650), .CP(clk), 
        .Q(inner_first_stage_data_reg[857]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_856_ ( .D(N6649), .CP(clk), 
        .Q(inner_first_stage_data_reg[856]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_855_ ( .D(N6648), .CP(clk), 
        .Q(inner_first_stage_data_reg[855]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_854_ ( .D(N6647), .CP(clk), 
        .Q(inner_first_stage_data_reg[854]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_853_ ( .D(N6646), .CP(clk), 
        .Q(inner_first_stage_data_reg[853]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_852_ ( .D(N6645), .CP(clk), 
        .Q(inner_first_stage_data_reg[852]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_851_ ( .D(N6644), .CP(clk), 
        .Q(inner_first_stage_data_reg[851]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_850_ ( .D(N6643), .CP(clk), 
        .Q(inner_first_stage_data_reg[850]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_849_ ( .D(N6642), .CP(clk), 
        .Q(inner_first_stage_data_reg[849]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_848_ ( .D(N6641), .CP(clk), 
        .Q(inner_first_stage_data_reg[848]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_847_ ( .D(N6640), .CP(clk), 
        .Q(inner_first_stage_data_reg[847]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_846_ ( .D(N6639), .CP(clk), 
        .Q(inner_first_stage_data_reg[846]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_845_ ( .D(N6638), .CP(clk), 
        .Q(inner_first_stage_data_reg[845]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_844_ ( .D(N6637), .CP(clk), 
        .Q(inner_first_stage_data_reg[844]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_843_ ( .D(N6636), .CP(clk), 
        .Q(inner_first_stage_data_reg[843]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_842_ ( .D(N6635), .CP(clk), 
        .Q(inner_first_stage_data_reg[842]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_841_ ( .D(N6634), .CP(clk), 
        .Q(inner_first_stage_data_reg[841]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_840_ ( .D(N6633), .CP(clk), 
        .Q(inner_first_stage_data_reg[840]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_839_ ( .D(N6632), .CP(clk), 
        .Q(inner_first_stage_data_reg[839]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_838_ ( .D(N6631), .CP(clk), 
        .Q(inner_first_stage_data_reg[838]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_837_ ( .D(N6630), .CP(clk), 
        .Q(inner_first_stage_data_reg[837]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_836_ ( .D(N6629), .CP(clk), 
        .Q(inner_first_stage_data_reg[836]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_835_ ( .D(N6628), .CP(clk), 
        .Q(inner_first_stage_data_reg[835]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_834_ ( .D(N6627), .CP(clk), 
        .Q(inner_first_stage_data_reg[834]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_833_ ( .D(N6626), .CP(clk), 
        .Q(inner_first_stage_data_reg[833]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_832_ ( .D(N6625), .CP(clk), 
        .Q(inner_first_stage_data_reg[832]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_26_ ( .D(N6624), .CP(clk), 
        .Q(inner_first_stage_valid_reg[26]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_895_ ( .D(N6872), .CP(clk), 
        .Q(inner_first_stage_data_reg[895]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_894_ ( .D(N6871), .CP(clk), 
        .Q(inner_first_stage_data_reg[894]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_893_ ( .D(N6870), .CP(clk), 
        .Q(inner_first_stage_data_reg[893]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_892_ ( .D(N6869), .CP(clk), 
        .Q(inner_first_stage_data_reg[892]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_891_ ( .D(N6868), .CP(clk), 
        .Q(inner_first_stage_data_reg[891]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_890_ ( .D(N6867), .CP(clk), 
        .Q(inner_first_stage_data_reg[890]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_889_ ( .D(N6866), .CP(clk), 
        .Q(inner_first_stage_data_reg[889]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_888_ ( .D(N6865), .CP(clk), 
        .Q(inner_first_stage_data_reg[888]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_887_ ( .D(N6864), .CP(clk), 
        .Q(inner_first_stage_data_reg[887]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_886_ ( .D(N6863), .CP(clk), 
        .Q(inner_first_stage_data_reg[886]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_885_ ( .D(N6862), .CP(clk), 
        .Q(inner_first_stage_data_reg[885]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_884_ ( .D(N6861), .CP(clk), 
        .Q(inner_first_stage_data_reg[884]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_883_ ( .D(N6860), .CP(clk), 
        .Q(inner_first_stage_data_reg[883]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_882_ ( .D(N6859), .CP(clk), 
        .Q(inner_first_stage_data_reg[882]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_881_ ( .D(N6858), .CP(clk), 
        .Q(inner_first_stage_data_reg[881]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_880_ ( .D(N6857), .CP(clk), 
        .Q(inner_first_stage_data_reg[880]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_879_ ( .D(N6856), .CP(clk), 
        .Q(inner_first_stage_data_reg[879]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_878_ ( .D(N6855), .CP(clk), 
        .Q(inner_first_stage_data_reg[878]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_877_ ( .D(N6854), .CP(clk), 
        .Q(inner_first_stage_data_reg[877]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_876_ ( .D(N6853), .CP(clk), 
        .Q(inner_first_stage_data_reg[876]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_875_ ( .D(N6852), .CP(clk), 
        .Q(inner_first_stage_data_reg[875]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_874_ ( .D(N6851), .CP(clk), 
        .Q(inner_first_stage_data_reg[874]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_873_ ( .D(N6850), .CP(clk), 
        .Q(inner_first_stage_data_reg[873]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_872_ ( .D(N6849), .CP(clk), 
        .Q(inner_first_stage_data_reg[872]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_871_ ( .D(N6848), .CP(clk), 
        .Q(inner_first_stage_data_reg[871]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_870_ ( .D(N6847), .CP(clk), 
        .Q(inner_first_stage_data_reg[870]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_869_ ( .D(N6846), .CP(clk), 
        .Q(inner_first_stage_data_reg[869]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_868_ ( .D(N6845), .CP(clk), 
        .Q(inner_first_stage_data_reg[868]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_867_ ( .D(N6844), .CP(clk), 
        .Q(inner_first_stage_data_reg[867]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_866_ ( .D(N6843), .CP(clk), 
        .Q(inner_first_stage_data_reg[866]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_865_ ( .D(N6842), .CP(clk), 
        .Q(inner_first_stage_data_reg[865]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_864_ ( .D(N6841), .CP(clk), 
        .Q(inner_first_stage_data_reg[864]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_27_ ( .D(N6840), .CP(clk), 
        .Q(inner_first_stage_valid_reg[27]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_927_ ( .D(N7088), .CP(clk), 
        .Q(inner_first_stage_data_reg[927]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_926_ ( .D(N7087), .CP(clk), 
        .Q(inner_first_stage_data_reg[926]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_925_ ( .D(N7086), .CP(clk), 
        .Q(inner_first_stage_data_reg[925]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_924_ ( .D(N7085), .CP(clk), 
        .Q(inner_first_stage_data_reg[924]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_923_ ( .D(N7084), .CP(clk), 
        .Q(inner_first_stage_data_reg[923]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_922_ ( .D(N7083), .CP(clk), 
        .Q(inner_first_stage_data_reg[922]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_921_ ( .D(N7082), .CP(clk), 
        .Q(inner_first_stage_data_reg[921]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_920_ ( .D(N7081), .CP(clk), 
        .Q(inner_first_stage_data_reg[920]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_919_ ( .D(N7080), .CP(clk), 
        .Q(inner_first_stage_data_reg[919]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_918_ ( .D(N7079), .CP(clk), 
        .Q(inner_first_stage_data_reg[918]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_917_ ( .D(N7078), .CP(clk), 
        .Q(inner_first_stage_data_reg[917]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_916_ ( .D(N7077), .CP(clk), 
        .Q(inner_first_stage_data_reg[916]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_915_ ( .D(N7076), .CP(clk), 
        .Q(inner_first_stage_data_reg[915]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_914_ ( .D(N7075), .CP(clk), 
        .Q(inner_first_stage_data_reg[914]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_913_ ( .D(N7074), .CP(clk), 
        .Q(inner_first_stage_data_reg[913]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_912_ ( .D(N7073), .CP(clk), 
        .Q(inner_first_stage_data_reg[912]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_911_ ( .D(N7072), .CP(clk), 
        .Q(inner_first_stage_data_reg[911]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_910_ ( .D(N7071), .CP(clk), 
        .Q(inner_first_stage_data_reg[910]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_909_ ( .D(N7070), .CP(clk), 
        .Q(inner_first_stage_data_reg[909]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_908_ ( .D(N7069), .CP(clk), 
        .Q(inner_first_stage_data_reg[908]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_907_ ( .D(N7068), .CP(clk), 
        .Q(inner_first_stage_data_reg[907]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_906_ ( .D(N7067), .CP(clk), 
        .Q(inner_first_stage_data_reg[906]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_905_ ( .D(N7066), .CP(clk), 
        .Q(inner_first_stage_data_reg[905]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_904_ ( .D(N7065), .CP(clk), 
        .Q(inner_first_stage_data_reg[904]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_903_ ( .D(N7064), .CP(clk), 
        .Q(inner_first_stage_data_reg[903]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_902_ ( .D(N7063), .CP(clk), 
        .Q(inner_first_stage_data_reg[902]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_901_ ( .D(N7062), .CP(clk), 
        .Q(inner_first_stage_data_reg[901]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_900_ ( .D(N7061), .CP(clk), 
        .Q(inner_first_stage_data_reg[900]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_899_ ( .D(N7060), .CP(clk), 
        .Q(inner_first_stage_data_reg[899]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_898_ ( .D(N7059), .CP(clk), 
        .Q(inner_first_stage_data_reg[898]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_897_ ( .D(N7058), .CP(clk), 
        .Q(inner_first_stage_data_reg[897]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_896_ ( .D(N7057), .CP(clk), 
        .Q(inner_first_stage_data_reg[896]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_28_ ( .D(N7056), .CP(clk), 
        .Q(inner_first_stage_valid_reg[28]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_959_ ( .D(N7304), .CP(clk), 
        .Q(inner_first_stage_data_reg[959]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_958_ ( .D(N7303), .CP(clk), 
        .Q(inner_first_stage_data_reg[958]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_957_ ( .D(N7302), .CP(clk), 
        .Q(inner_first_stage_data_reg[957]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_956_ ( .D(N7301), .CP(clk), 
        .Q(inner_first_stage_data_reg[956]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_955_ ( .D(N7300), .CP(clk), 
        .Q(inner_first_stage_data_reg[955]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_954_ ( .D(N7299), .CP(clk), 
        .Q(inner_first_stage_data_reg[954]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_953_ ( .D(N7298), .CP(clk), 
        .Q(inner_first_stage_data_reg[953]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_952_ ( .D(N7297), .CP(clk), 
        .Q(inner_first_stage_data_reg[952]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_951_ ( .D(N7296), .CP(clk), 
        .Q(inner_first_stage_data_reg[951]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_950_ ( .D(N7295), .CP(clk), 
        .Q(inner_first_stage_data_reg[950]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_949_ ( .D(N7294), .CP(clk), 
        .Q(inner_first_stage_data_reg[949]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_948_ ( .D(N7293), .CP(clk), 
        .Q(inner_first_stage_data_reg[948]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_947_ ( .D(N7292), .CP(clk), 
        .Q(inner_first_stage_data_reg[947]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_946_ ( .D(N7291), .CP(clk), 
        .Q(inner_first_stage_data_reg[946]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_945_ ( .D(N7290), .CP(clk), 
        .Q(inner_first_stage_data_reg[945]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_944_ ( .D(N7289), .CP(clk), 
        .Q(inner_first_stage_data_reg[944]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_943_ ( .D(N7288), .CP(clk), 
        .Q(inner_first_stage_data_reg[943]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_942_ ( .D(N7287), .CP(clk), 
        .Q(inner_first_stage_data_reg[942]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_941_ ( .D(N7286), .CP(clk), 
        .Q(inner_first_stage_data_reg[941]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_940_ ( .D(N7285), .CP(clk), 
        .Q(inner_first_stage_data_reg[940]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_939_ ( .D(N7284), .CP(clk), 
        .Q(inner_first_stage_data_reg[939]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_938_ ( .D(N7283), .CP(clk), 
        .Q(inner_first_stage_data_reg[938]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_937_ ( .D(N7282), .CP(clk), 
        .Q(inner_first_stage_data_reg[937]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_936_ ( .D(N7281), .CP(clk), 
        .Q(inner_first_stage_data_reg[936]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_935_ ( .D(N7280), .CP(clk), 
        .Q(inner_first_stage_data_reg[935]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_934_ ( .D(N7279), .CP(clk), 
        .Q(inner_first_stage_data_reg[934]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_933_ ( .D(N7278), .CP(clk), 
        .Q(inner_first_stage_data_reg[933]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_932_ ( .D(N7277), .CP(clk), 
        .Q(inner_first_stage_data_reg[932]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_931_ ( .D(N7276), .CP(clk), 
        .Q(inner_first_stage_data_reg[931]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_930_ ( .D(N7275), .CP(clk), 
        .Q(inner_first_stage_data_reg[930]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_929_ ( .D(N7274), .CP(clk), 
        .Q(inner_first_stage_data_reg[929]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_928_ ( .D(N7273), .CP(clk), 
        .Q(inner_first_stage_data_reg[928]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_29_ ( .D(N7272), .CP(clk), 
        .Q(inner_first_stage_valid_reg[29]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_991_ ( .D(N7520), .CP(clk), 
        .Q(inner_first_stage_data_reg[991]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_990_ ( .D(N7519), .CP(clk), 
        .Q(inner_first_stage_data_reg[990]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_989_ ( .D(N7518), .CP(clk), 
        .Q(inner_first_stage_data_reg[989]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_988_ ( .D(N7517), .CP(clk), 
        .Q(inner_first_stage_data_reg[988]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_987_ ( .D(N7516), .CP(clk), 
        .Q(inner_first_stage_data_reg[987]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_986_ ( .D(N7515), .CP(clk), 
        .Q(inner_first_stage_data_reg[986]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_985_ ( .D(N7514), .CP(clk), 
        .Q(inner_first_stage_data_reg[985]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_984_ ( .D(N7513), .CP(clk), 
        .Q(inner_first_stage_data_reg[984]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_983_ ( .D(N7512), .CP(clk), 
        .Q(inner_first_stage_data_reg[983]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_982_ ( .D(N7511), .CP(clk), 
        .Q(inner_first_stage_data_reg[982]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_981_ ( .D(N7510), .CP(clk), 
        .Q(inner_first_stage_data_reg[981]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_980_ ( .D(N7509), .CP(clk), 
        .Q(inner_first_stage_data_reg[980]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_979_ ( .D(N7508), .CP(clk), 
        .Q(inner_first_stage_data_reg[979]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_978_ ( .D(N7507), .CP(clk), 
        .Q(inner_first_stage_data_reg[978]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_977_ ( .D(N7506), .CP(clk), 
        .Q(inner_first_stage_data_reg[977]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_976_ ( .D(N7505), .CP(clk), 
        .Q(inner_first_stage_data_reg[976]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_975_ ( .D(N7504), .CP(clk), 
        .Q(inner_first_stage_data_reg[975]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_974_ ( .D(N7503), .CP(clk), 
        .Q(inner_first_stage_data_reg[974]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_973_ ( .D(N7502), .CP(clk), 
        .Q(inner_first_stage_data_reg[973]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_972_ ( .D(N7501), .CP(clk), 
        .Q(inner_first_stage_data_reg[972]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_971_ ( .D(N7500), .CP(clk), 
        .Q(inner_first_stage_data_reg[971]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_970_ ( .D(N7499), .CP(clk), 
        .Q(inner_first_stage_data_reg[970]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_969_ ( .D(N7498), .CP(clk), 
        .Q(inner_first_stage_data_reg[969]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_968_ ( .D(N7497), .CP(clk), 
        .Q(inner_first_stage_data_reg[968]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_967_ ( .D(N7496), .CP(clk), 
        .Q(inner_first_stage_data_reg[967]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_966_ ( .D(N7495), .CP(clk), 
        .Q(inner_first_stage_data_reg[966]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_965_ ( .D(N7494), .CP(clk), 
        .Q(inner_first_stage_data_reg[965]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_964_ ( .D(N7493), .CP(clk), 
        .Q(inner_first_stage_data_reg[964]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_963_ ( .D(N7492), .CP(clk), 
        .Q(inner_first_stage_data_reg[963]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_962_ ( .D(N7491), .CP(clk), 
        .Q(inner_first_stage_data_reg[962]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_961_ ( .D(N7490), .CP(clk), 
        .Q(inner_first_stage_data_reg[961]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_960_ ( .D(N7489), .CP(clk), 
        .Q(inner_first_stage_data_reg[960]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_30_ ( .D(N7488), .CP(clk), 
        .Q(inner_first_stage_valid_reg[30]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1023_ ( .D(N7736), .CP(clk), 
        .Q(inner_first_stage_data_reg[1023]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1022_ ( .D(N7735), .CP(clk), 
        .Q(inner_first_stage_data_reg[1022]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1021_ ( .D(N7734), .CP(clk), 
        .Q(inner_first_stage_data_reg[1021]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1020_ ( .D(N7733), .CP(clk), 
        .Q(inner_first_stage_data_reg[1020]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1019_ ( .D(N7732), .CP(clk), 
        .Q(inner_first_stage_data_reg[1019]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1018_ ( .D(N7731), .CP(clk), 
        .Q(inner_first_stage_data_reg[1018]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1017_ ( .D(N7730), .CP(clk), 
        .Q(inner_first_stage_data_reg[1017]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1016_ ( .D(N7729), .CP(clk), 
        .Q(inner_first_stage_data_reg[1016]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1015_ ( .D(N7728), .CP(clk), 
        .Q(inner_first_stage_data_reg[1015]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1014_ ( .D(N7727), .CP(clk), 
        .Q(inner_first_stage_data_reg[1014]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1013_ ( .D(N7726), .CP(clk), 
        .Q(inner_first_stage_data_reg[1013]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1012_ ( .D(N7725), .CP(clk), 
        .Q(inner_first_stage_data_reg[1012]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1011_ ( .D(N7724), .CP(clk), 
        .Q(inner_first_stage_data_reg[1011]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1010_ ( .D(N7723), .CP(clk), 
        .Q(inner_first_stage_data_reg[1010]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1009_ ( .D(N7722), .CP(clk), 
        .Q(inner_first_stage_data_reg[1009]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1008_ ( .D(N7721), .CP(clk), 
        .Q(inner_first_stage_data_reg[1008]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1007_ ( .D(N7720), .CP(clk), 
        .Q(inner_first_stage_data_reg[1007]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1006_ ( .D(N7719), .CP(clk), 
        .Q(inner_first_stage_data_reg[1006]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1005_ ( .D(N7718), .CP(clk), 
        .Q(inner_first_stage_data_reg[1005]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1004_ ( .D(N7717), .CP(clk), 
        .Q(inner_first_stage_data_reg[1004]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1003_ ( .D(N7716), .CP(clk), 
        .Q(inner_first_stage_data_reg[1003]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1002_ ( .D(N7715), .CP(clk), 
        .Q(inner_first_stage_data_reg[1002]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1001_ ( .D(N7714), .CP(clk), 
        .Q(inner_first_stage_data_reg[1001]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1000_ ( .D(N7713), .CP(clk), 
        .Q(inner_first_stage_data_reg[1000]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_999_ ( .D(N7712), .CP(clk), 
        .Q(inner_first_stage_data_reg[999]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_998_ ( .D(N7711), .CP(clk), 
        .Q(inner_first_stage_data_reg[998]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_997_ ( .D(N7710), .CP(clk), 
        .Q(inner_first_stage_data_reg[997]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_996_ ( .D(N7709), .CP(clk), 
        .Q(inner_first_stage_data_reg[996]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_995_ ( .D(N7708), .CP(clk), 
        .Q(inner_first_stage_data_reg[995]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_994_ ( .D(N7707), .CP(clk), 
        .Q(inner_first_stage_data_reg[994]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_993_ ( .D(N7706), .CP(clk), 
        .Q(inner_first_stage_data_reg[993]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_992_ ( .D(N7705), .CP(clk), 
        .Q(inner_first_stage_data_reg[992]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_31_ ( .D(N7704), .CP(clk), 
        .Q(inner_first_stage_valid_reg[31]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1055_ ( .D(N8098), .CP(clk), 
        .Q(inner_first_stage_data_reg[1055]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1054_ ( .D(N8097), .CP(clk), 
        .Q(inner_first_stage_data_reg[1054]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1053_ ( .D(N8096), .CP(clk), 
        .Q(inner_first_stage_data_reg[1053]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1052_ ( .D(N8095), .CP(clk), 
        .Q(inner_first_stage_data_reg[1052]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1051_ ( .D(N8094), .CP(clk), 
        .Q(inner_first_stage_data_reg[1051]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1050_ ( .D(N8093), .CP(clk), 
        .Q(inner_first_stage_data_reg[1050]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1049_ ( .D(N8092), .CP(clk), 
        .Q(inner_first_stage_data_reg[1049]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1048_ ( .D(N8091), .CP(clk), 
        .Q(inner_first_stage_data_reg[1048]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1047_ ( .D(N8090), .CP(clk), 
        .Q(inner_first_stage_data_reg[1047]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1046_ ( .D(N8089), .CP(clk), 
        .Q(inner_first_stage_data_reg[1046]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1045_ ( .D(N8088), .CP(clk), 
        .Q(inner_first_stage_data_reg[1045]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1044_ ( .D(N8087), .CP(clk), 
        .Q(inner_first_stage_data_reg[1044]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1043_ ( .D(N8086), .CP(clk), 
        .Q(inner_first_stage_data_reg[1043]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1042_ ( .D(N8085), .CP(clk), 
        .Q(inner_first_stage_data_reg[1042]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1041_ ( .D(N8084), .CP(clk), 
        .Q(inner_first_stage_data_reg[1041]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1040_ ( .D(N8083), .CP(clk), 
        .Q(inner_first_stage_data_reg[1040]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1039_ ( .D(N8082), .CP(clk), 
        .Q(inner_first_stage_data_reg[1039]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1038_ ( .D(N8081), .CP(clk), 
        .Q(inner_first_stage_data_reg[1038]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1037_ ( .D(N8080), .CP(clk), 
        .Q(inner_first_stage_data_reg[1037]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1036_ ( .D(N8079), .CP(clk), 
        .Q(inner_first_stage_data_reg[1036]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1035_ ( .D(N8078), .CP(clk), 
        .Q(inner_first_stage_data_reg[1035]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1034_ ( .D(N8077), .CP(clk), 
        .Q(inner_first_stage_data_reg[1034]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1033_ ( .D(N8076), .CP(clk), 
        .Q(inner_first_stage_data_reg[1033]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1032_ ( .D(N8075), .CP(clk), 
        .Q(inner_first_stage_data_reg[1032]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1031_ ( .D(N8074), .CP(clk), 
        .Q(inner_first_stage_data_reg[1031]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1030_ ( .D(N8073), .CP(clk), 
        .Q(inner_first_stage_data_reg[1030]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1029_ ( .D(N8072), .CP(clk), 
        .Q(inner_first_stage_data_reg[1029]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1028_ ( .D(N8071), .CP(clk), 
        .Q(inner_first_stage_data_reg[1028]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1027_ ( .D(N8070), .CP(clk), 
        .Q(inner_first_stage_data_reg[1027]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1026_ ( .D(N8069), .CP(clk), 
        .Q(inner_first_stage_data_reg[1026]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1025_ ( .D(N8068), .CP(clk), 
        .Q(inner_first_stage_data_reg[1025]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1024_ ( .D(N8067), .CP(clk), 
        .Q(inner_first_stage_data_reg[1024]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_32_ ( .D(N8066), .CP(clk), 
        .Q(inner_first_stage_valid_reg[32]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1087_ ( .D(N8314), .CP(clk), 
        .Q(inner_first_stage_data_reg[1087]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1086_ ( .D(N8313), .CP(clk), 
        .Q(inner_first_stage_data_reg[1086]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1085_ ( .D(N8312), .CP(clk), 
        .Q(inner_first_stage_data_reg[1085]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1084_ ( .D(N8311), .CP(clk), 
        .Q(inner_first_stage_data_reg[1084]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1083_ ( .D(N8310), .CP(clk), 
        .Q(inner_first_stage_data_reg[1083]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1082_ ( .D(N8309), .CP(clk), 
        .Q(inner_first_stage_data_reg[1082]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1081_ ( .D(N8308), .CP(clk), 
        .Q(inner_first_stage_data_reg[1081]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1080_ ( .D(N8307), .CP(clk), 
        .Q(inner_first_stage_data_reg[1080]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1079_ ( .D(N8306), .CP(clk), 
        .Q(inner_first_stage_data_reg[1079]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1078_ ( .D(N8305), .CP(clk), 
        .Q(inner_first_stage_data_reg[1078]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1077_ ( .D(N8304), .CP(clk), 
        .Q(inner_first_stage_data_reg[1077]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1076_ ( .D(N8303), .CP(clk), 
        .Q(inner_first_stage_data_reg[1076]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1075_ ( .D(N8302), .CP(clk), 
        .Q(inner_first_stage_data_reg[1075]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1074_ ( .D(N8301), .CP(clk), 
        .Q(inner_first_stage_data_reg[1074]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1073_ ( .D(N8300), .CP(clk), 
        .Q(inner_first_stage_data_reg[1073]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1072_ ( .D(N8299), .CP(clk), 
        .Q(inner_first_stage_data_reg[1072]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1071_ ( .D(N8298), .CP(clk), 
        .Q(inner_first_stage_data_reg[1071]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1070_ ( .D(N8297), .CP(clk), 
        .Q(inner_first_stage_data_reg[1070]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1069_ ( .D(N8296), .CP(clk), 
        .Q(inner_first_stage_data_reg[1069]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1068_ ( .D(N8295), .CP(clk), 
        .Q(inner_first_stage_data_reg[1068]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1067_ ( .D(N8294), .CP(clk), 
        .Q(inner_first_stage_data_reg[1067]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1066_ ( .D(N8293), .CP(clk), 
        .Q(inner_first_stage_data_reg[1066]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1065_ ( .D(N8292), .CP(clk), 
        .Q(inner_first_stage_data_reg[1065]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1064_ ( .D(N8291), .CP(clk), 
        .Q(inner_first_stage_data_reg[1064]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1063_ ( .D(N8290), .CP(clk), 
        .Q(inner_first_stage_data_reg[1063]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1062_ ( .D(N8289), .CP(clk), 
        .Q(inner_first_stage_data_reg[1062]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1061_ ( .D(N8288), .CP(clk), 
        .Q(inner_first_stage_data_reg[1061]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1060_ ( .D(N8287), .CP(clk), 
        .Q(inner_first_stage_data_reg[1060]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1059_ ( .D(N8286), .CP(clk), 
        .Q(inner_first_stage_data_reg[1059]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1058_ ( .D(N8285), .CP(clk), 
        .Q(inner_first_stage_data_reg[1058]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1057_ ( .D(N8284), .CP(clk), 
        .Q(inner_first_stage_data_reg[1057]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1056_ ( .D(N8283), .CP(clk), 
        .Q(inner_first_stage_data_reg[1056]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_33_ ( .D(N8282), .CP(clk), 
        .Q(inner_first_stage_valid_reg[33]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1119_ ( .D(N8530), .CP(clk), 
        .Q(inner_first_stage_data_reg[1119]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1118_ ( .D(N8529), .CP(clk), 
        .Q(inner_first_stage_data_reg[1118]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1117_ ( .D(N8528), .CP(clk), 
        .Q(inner_first_stage_data_reg[1117]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1116_ ( .D(N8527), .CP(clk), 
        .Q(inner_first_stage_data_reg[1116]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1115_ ( .D(N8526), .CP(clk), 
        .Q(inner_first_stage_data_reg[1115]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1114_ ( .D(N8525), .CP(clk), 
        .Q(inner_first_stage_data_reg[1114]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1113_ ( .D(N8524), .CP(clk), 
        .Q(inner_first_stage_data_reg[1113]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1112_ ( .D(N8523), .CP(clk), 
        .Q(inner_first_stage_data_reg[1112]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1111_ ( .D(N8522), .CP(clk), 
        .Q(inner_first_stage_data_reg[1111]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1110_ ( .D(N8521), .CP(clk), 
        .Q(inner_first_stage_data_reg[1110]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1109_ ( .D(N8520), .CP(clk), 
        .Q(inner_first_stage_data_reg[1109]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1108_ ( .D(N8519), .CP(clk), 
        .Q(inner_first_stage_data_reg[1108]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1107_ ( .D(N8518), .CP(clk), 
        .Q(inner_first_stage_data_reg[1107]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1106_ ( .D(N8517), .CP(clk), 
        .Q(inner_first_stage_data_reg[1106]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1105_ ( .D(N8516), .CP(clk), 
        .Q(inner_first_stage_data_reg[1105]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1104_ ( .D(N8515), .CP(clk), 
        .Q(inner_first_stage_data_reg[1104]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1103_ ( .D(N8514), .CP(clk), 
        .Q(inner_first_stage_data_reg[1103]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1102_ ( .D(N8513), .CP(clk), 
        .Q(inner_first_stage_data_reg[1102]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1101_ ( .D(N8512), .CP(clk), 
        .Q(inner_first_stage_data_reg[1101]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1100_ ( .D(N8511), .CP(clk), 
        .Q(inner_first_stage_data_reg[1100]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1099_ ( .D(N8510), .CP(clk), 
        .Q(inner_first_stage_data_reg[1099]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1098_ ( .D(N8509), .CP(clk), 
        .Q(inner_first_stage_data_reg[1098]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1097_ ( .D(N8508), .CP(clk), 
        .Q(inner_first_stage_data_reg[1097]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1096_ ( .D(N8507), .CP(clk), 
        .Q(inner_first_stage_data_reg[1096]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1095_ ( .D(N8506), .CP(clk), 
        .Q(inner_first_stage_data_reg[1095]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1094_ ( .D(N8505), .CP(clk), 
        .Q(inner_first_stage_data_reg[1094]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1093_ ( .D(N8504), .CP(clk), 
        .Q(inner_first_stage_data_reg[1093]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1092_ ( .D(N8503), .CP(clk), 
        .Q(inner_first_stage_data_reg[1092]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1091_ ( .D(N8502), .CP(clk), 
        .Q(inner_first_stage_data_reg[1091]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1090_ ( .D(N8501), .CP(clk), 
        .Q(inner_first_stage_data_reg[1090]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1089_ ( .D(N8500), .CP(clk), 
        .Q(inner_first_stage_data_reg[1089]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1088_ ( .D(N8499), .CP(clk), 
        .Q(inner_first_stage_data_reg[1088]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_34_ ( .D(N8498), .CP(clk), 
        .Q(inner_first_stage_valid_reg[34]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1151_ ( .D(N8746), .CP(clk), 
        .Q(inner_first_stage_data_reg[1151]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1150_ ( .D(N8745), .CP(clk), 
        .Q(inner_first_stage_data_reg[1150]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1149_ ( .D(N8744), .CP(clk), 
        .Q(inner_first_stage_data_reg[1149]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1148_ ( .D(N8743), .CP(clk), 
        .Q(inner_first_stage_data_reg[1148]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1147_ ( .D(N8742), .CP(clk), 
        .Q(inner_first_stage_data_reg[1147]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1146_ ( .D(N8741), .CP(clk), 
        .Q(inner_first_stage_data_reg[1146]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1145_ ( .D(N8740), .CP(clk), 
        .Q(inner_first_stage_data_reg[1145]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1144_ ( .D(N8739), .CP(clk), 
        .Q(inner_first_stage_data_reg[1144]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1143_ ( .D(N8738), .CP(clk), 
        .Q(inner_first_stage_data_reg[1143]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1142_ ( .D(N8737), .CP(clk), 
        .Q(inner_first_stage_data_reg[1142]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1141_ ( .D(N8736), .CP(clk), 
        .Q(inner_first_stage_data_reg[1141]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1140_ ( .D(N8735), .CP(clk), 
        .Q(inner_first_stage_data_reg[1140]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1139_ ( .D(N8734), .CP(clk), 
        .Q(inner_first_stage_data_reg[1139]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1138_ ( .D(N8733), .CP(clk), 
        .Q(inner_first_stage_data_reg[1138]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1137_ ( .D(N8732), .CP(clk), 
        .Q(inner_first_stage_data_reg[1137]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1136_ ( .D(N8731), .CP(clk), 
        .Q(inner_first_stage_data_reg[1136]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1135_ ( .D(N8730), .CP(clk), 
        .Q(inner_first_stage_data_reg[1135]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1134_ ( .D(N8729), .CP(clk), 
        .Q(inner_first_stage_data_reg[1134]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1133_ ( .D(N8728), .CP(clk), 
        .Q(inner_first_stage_data_reg[1133]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1132_ ( .D(N8727), .CP(clk), 
        .Q(inner_first_stage_data_reg[1132]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1131_ ( .D(N8726), .CP(clk), 
        .Q(inner_first_stage_data_reg[1131]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1130_ ( .D(N8725), .CP(clk), 
        .Q(inner_first_stage_data_reg[1130]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1129_ ( .D(N8724), .CP(clk), 
        .Q(inner_first_stage_data_reg[1129]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1128_ ( .D(N8723), .CP(clk), 
        .Q(inner_first_stage_data_reg[1128]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1127_ ( .D(N8722), .CP(clk), 
        .Q(inner_first_stage_data_reg[1127]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1126_ ( .D(N8721), .CP(clk), 
        .Q(inner_first_stage_data_reg[1126]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1125_ ( .D(N8720), .CP(clk), 
        .Q(inner_first_stage_data_reg[1125]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1124_ ( .D(N8719), .CP(clk), 
        .Q(inner_first_stage_data_reg[1124]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1123_ ( .D(N8718), .CP(clk), 
        .Q(inner_first_stage_data_reg[1123]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1122_ ( .D(N8717), .CP(clk), 
        .Q(inner_first_stage_data_reg[1122]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1121_ ( .D(N8716), .CP(clk), 
        .Q(inner_first_stage_data_reg[1121]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1120_ ( .D(N8715), .CP(clk), 
        .Q(inner_first_stage_data_reg[1120]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_35_ ( .D(N8714), .CP(clk), 
        .Q(inner_first_stage_valid_reg[35]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1183_ ( .D(N8962), .CP(clk), 
        .Q(inner_first_stage_data_reg[1183]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1182_ ( .D(N8961), .CP(clk), 
        .Q(inner_first_stage_data_reg[1182]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1181_ ( .D(N8960), .CP(clk), 
        .Q(inner_first_stage_data_reg[1181]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1180_ ( .D(N8959), .CP(clk), 
        .Q(inner_first_stage_data_reg[1180]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1179_ ( .D(N8958), .CP(clk), 
        .Q(inner_first_stage_data_reg[1179]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1178_ ( .D(N8957), .CP(clk), 
        .Q(inner_first_stage_data_reg[1178]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1177_ ( .D(N8956), .CP(clk), 
        .Q(inner_first_stage_data_reg[1177]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1176_ ( .D(N8955), .CP(clk), 
        .Q(inner_first_stage_data_reg[1176]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1175_ ( .D(N8954), .CP(clk), 
        .Q(inner_first_stage_data_reg[1175]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1174_ ( .D(N8953), .CP(clk), 
        .Q(inner_first_stage_data_reg[1174]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1173_ ( .D(N8952), .CP(clk), 
        .Q(inner_first_stage_data_reg[1173]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1172_ ( .D(N8951), .CP(clk), 
        .Q(inner_first_stage_data_reg[1172]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1171_ ( .D(N8950), .CP(clk), 
        .Q(inner_first_stage_data_reg[1171]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1170_ ( .D(N8949), .CP(clk), 
        .Q(inner_first_stage_data_reg[1170]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1169_ ( .D(N8948), .CP(clk), 
        .Q(inner_first_stage_data_reg[1169]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1168_ ( .D(N8947), .CP(clk), 
        .Q(inner_first_stage_data_reg[1168]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1167_ ( .D(N8946), .CP(clk), 
        .Q(inner_first_stage_data_reg[1167]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1166_ ( .D(N8945), .CP(clk), 
        .Q(inner_first_stage_data_reg[1166]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1165_ ( .D(N8944), .CP(clk), 
        .Q(inner_first_stage_data_reg[1165]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1164_ ( .D(N8943), .CP(clk), 
        .Q(inner_first_stage_data_reg[1164]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1163_ ( .D(N8942), .CP(clk), 
        .Q(inner_first_stage_data_reg[1163]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1162_ ( .D(N8941), .CP(clk), 
        .Q(inner_first_stage_data_reg[1162]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1161_ ( .D(N8940), .CP(clk), 
        .Q(inner_first_stage_data_reg[1161]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1160_ ( .D(N8939), .CP(clk), 
        .Q(inner_first_stage_data_reg[1160]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1159_ ( .D(N8938), .CP(clk), 
        .Q(inner_first_stage_data_reg[1159]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1158_ ( .D(N8937), .CP(clk), 
        .Q(inner_first_stage_data_reg[1158]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1157_ ( .D(N8936), .CP(clk), 
        .Q(inner_first_stage_data_reg[1157]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1156_ ( .D(N8935), .CP(clk), 
        .Q(inner_first_stage_data_reg[1156]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1155_ ( .D(N8934), .CP(clk), 
        .Q(inner_first_stage_data_reg[1155]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1154_ ( .D(N8933), .CP(clk), 
        .Q(inner_first_stage_data_reg[1154]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1153_ ( .D(N8932), .CP(clk), 
        .Q(inner_first_stage_data_reg[1153]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1152_ ( .D(N8931), .CP(clk), 
        .Q(inner_first_stage_data_reg[1152]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_36_ ( .D(N8930), .CP(clk), 
        .Q(inner_first_stage_valid_reg[36]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1215_ ( .D(N9178), .CP(clk), 
        .Q(inner_first_stage_data_reg[1215]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1214_ ( .D(N9177), .CP(clk), 
        .Q(inner_first_stage_data_reg[1214]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1213_ ( .D(N9176), .CP(clk), 
        .Q(inner_first_stage_data_reg[1213]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1212_ ( .D(N9175), .CP(clk), 
        .Q(inner_first_stage_data_reg[1212]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1211_ ( .D(N9174), .CP(clk), 
        .Q(inner_first_stage_data_reg[1211]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1210_ ( .D(N9173), .CP(clk), 
        .Q(inner_first_stage_data_reg[1210]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1209_ ( .D(N9172), .CP(clk), 
        .Q(inner_first_stage_data_reg[1209]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1208_ ( .D(N9171), .CP(clk), 
        .Q(inner_first_stage_data_reg[1208]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1207_ ( .D(N9170), .CP(clk), 
        .Q(inner_first_stage_data_reg[1207]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1206_ ( .D(N9169), .CP(clk), 
        .Q(inner_first_stage_data_reg[1206]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1205_ ( .D(N9168), .CP(clk), 
        .Q(inner_first_stage_data_reg[1205]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1204_ ( .D(N9167), .CP(clk), 
        .Q(inner_first_stage_data_reg[1204]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1203_ ( .D(N9166), .CP(clk), 
        .Q(inner_first_stage_data_reg[1203]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1202_ ( .D(N9165), .CP(clk), 
        .Q(inner_first_stage_data_reg[1202]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1201_ ( .D(N9164), .CP(clk), 
        .Q(inner_first_stage_data_reg[1201]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1200_ ( .D(N9163), .CP(clk), 
        .Q(inner_first_stage_data_reg[1200]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1199_ ( .D(N9162), .CP(clk), 
        .Q(inner_first_stage_data_reg[1199]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1198_ ( .D(N9161), .CP(clk), 
        .Q(inner_first_stage_data_reg[1198]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1197_ ( .D(N9160), .CP(clk), 
        .Q(inner_first_stage_data_reg[1197]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1196_ ( .D(N9159), .CP(clk), 
        .Q(inner_first_stage_data_reg[1196]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1195_ ( .D(N9158), .CP(clk), 
        .Q(inner_first_stage_data_reg[1195]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1194_ ( .D(N9157), .CP(clk), 
        .Q(inner_first_stage_data_reg[1194]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1193_ ( .D(N9156), .CP(clk), 
        .Q(inner_first_stage_data_reg[1193]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1192_ ( .D(N9155), .CP(clk), 
        .Q(inner_first_stage_data_reg[1192]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1191_ ( .D(N9154), .CP(clk), 
        .Q(inner_first_stage_data_reg[1191]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1190_ ( .D(N9153), .CP(clk), 
        .Q(inner_first_stage_data_reg[1190]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1189_ ( .D(N9152), .CP(clk), 
        .Q(inner_first_stage_data_reg[1189]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1188_ ( .D(N9151), .CP(clk), 
        .Q(inner_first_stage_data_reg[1188]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1187_ ( .D(N9150), .CP(clk), 
        .Q(inner_first_stage_data_reg[1187]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1186_ ( .D(N9149), .CP(clk), 
        .Q(inner_first_stage_data_reg[1186]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1185_ ( .D(N9148), .CP(clk), 
        .Q(inner_first_stage_data_reg[1185]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1184_ ( .D(N9147), .CP(clk), 
        .Q(inner_first_stage_data_reg[1184]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_37_ ( .D(N9146), .CP(clk), 
        .Q(inner_first_stage_valid_reg[37]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1247_ ( .D(N9394), .CP(clk), 
        .Q(inner_first_stage_data_reg[1247]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1246_ ( .D(N9393), .CP(clk), 
        .Q(inner_first_stage_data_reg[1246]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1245_ ( .D(N9392), .CP(clk), 
        .Q(inner_first_stage_data_reg[1245]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1244_ ( .D(N9391), .CP(clk), 
        .Q(inner_first_stage_data_reg[1244]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1243_ ( .D(N9390), .CP(clk), 
        .Q(inner_first_stage_data_reg[1243]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1242_ ( .D(N9389), .CP(clk), 
        .Q(inner_first_stage_data_reg[1242]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1241_ ( .D(N9388), .CP(clk), 
        .Q(inner_first_stage_data_reg[1241]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1240_ ( .D(N9387), .CP(clk), 
        .Q(inner_first_stage_data_reg[1240]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1239_ ( .D(N9386), .CP(clk), 
        .Q(inner_first_stage_data_reg[1239]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1238_ ( .D(N9385), .CP(clk), 
        .Q(inner_first_stage_data_reg[1238]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1237_ ( .D(N9384), .CP(clk), 
        .Q(inner_first_stage_data_reg[1237]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1236_ ( .D(N9383), .CP(clk), 
        .Q(inner_first_stage_data_reg[1236]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1235_ ( .D(N9382), .CP(clk), 
        .Q(inner_first_stage_data_reg[1235]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1234_ ( .D(N9381), .CP(clk), 
        .Q(inner_first_stage_data_reg[1234]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1233_ ( .D(N9380), .CP(clk), 
        .Q(inner_first_stage_data_reg[1233]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1232_ ( .D(N9379), .CP(clk), 
        .Q(inner_first_stage_data_reg[1232]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1231_ ( .D(N9378), .CP(clk), 
        .Q(inner_first_stage_data_reg[1231]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1230_ ( .D(N9377), .CP(clk), 
        .Q(inner_first_stage_data_reg[1230]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1229_ ( .D(N9376), .CP(clk), 
        .Q(inner_first_stage_data_reg[1229]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1228_ ( .D(N9375), .CP(clk), 
        .Q(inner_first_stage_data_reg[1228]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1227_ ( .D(N9374), .CP(clk), 
        .Q(inner_first_stage_data_reg[1227]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1226_ ( .D(N9373), .CP(clk), 
        .Q(inner_first_stage_data_reg[1226]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1225_ ( .D(N9372), .CP(clk), 
        .Q(inner_first_stage_data_reg[1225]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1224_ ( .D(N9371), .CP(clk), 
        .Q(inner_first_stage_data_reg[1224]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1223_ ( .D(N9370), .CP(clk), 
        .Q(inner_first_stage_data_reg[1223]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1222_ ( .D(N9369), .CP(clk), 
        .Q(inner_first_stage_data_reg[1222]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1221_ ( .D(N9368), .CP(clk), 
        .Q(inner_first_stage_data_reg[1221]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1220_ ( .D(N9367), .CP(clk), 
        .Q(inner_first_stage_data_reg[1220]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1219_ ( .D(N9366), .CP(clk), 
        .Q(inner_first_stage_data_reg[1219]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1218_ ( .D(N9365), .CP(clk), 
        .Q(inner_first_stage_data_reg[1218]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1217_ ( .D(N9364), .CP(clk), 
        .Q(inner_first_stage_data_reg[1217]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1216_ ( .D(N9363), .CP(clk), 
        .Q(inner_first_stage_data_reg[1216]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_38_ ( .D(N9362), .CP(clk), 
        .Q(inner_first_stage_valid_reg[38]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1279_ ( .D(N9610), .CP(clk), 
        .Q(inner_first_stage_data_reg[1279]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1278_ ( .D(N9609), .CP(clk), 
        .Q(inner_first_stage_data_reg[1278]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1277_ ( .D(N9608), .CP(clk), 
        .Q(inner_first_stage_data_reg[1277]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1276_ ( .D(N9607), .CP(clk), 
        .Q(inner_first_stage_data_reg[1276]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1275_ ( .D(N9606), .CP(clk), 
        .Q(inner_first_stage_data_reg[1275]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1274_ ( .D(N9605), .CP(clk), 
        .Q(inner_first_stage_data_reg[1274]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1273_ ( .D(N9604), .CP(clk), 
        .Q(inner_first_stage_data_reg[1273]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1272_ ( .D(N9603), .CP(clk), 
        .Q(inner_first_stage_data_reg[1272]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1271_ ( .D(N9602), .CP(clk), 
        .Q(inner_first_stage_data_reg[1271]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1270_ ( .D(N9601), .CP(clk), 
        .Q(inner_first_stage_data_reg[1270]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1269_ ( .D(N9600), .CP(clk), 
        .Q(inner_first_stage_data_reg[1269]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1268_ ( .D(N9599), .CP(clk), 
        .Q(inner_first_stage_data_reg[1268]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1267_ ( .D(N9598), .CP(clk), 
        .Q(inner_first_stage_data_reg[1267]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1266_ ( .D(N9597), .CP(clk), 
        .Q(inner_first_stage_data_reg[1266]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1265_ ( .D(N9596), .CP(clk), 
        .Q(inner_first_stage_data_reg[1265]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1264_ ( .D(N9595), .CP(clk), 
        .Q(inner_first_stage_data_reg[1264]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1263_ ( .D(N9594), .CP(clk), 
        .Q(inner_first_stage_data_reg[1263]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1262_ ( .D(N9593), .CP(clk), 
        .Q(inner_first_stage_data_reg[1262]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1261_ ( .D(N9592), .CP(clk), 
        .Q(inner_first_stage_data_reg[1261]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1260_ ( .D(N9591), .CP(clk), 
        .Q(inner_first_stage_data_reg[1260]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1259_ ( .D(N9590), .CP(clk), 
        .Q(inner_first_stage_data_reg[1259]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1258_ ( .D(N9589), .CP(clk), 
        .Q(inner_first_stage_data_reg[1258]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1257_ ( .D(N9588), .CP(clk), 
        .Q(inner_first_stage_data_reg[1257]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1256_ ( .D(N9587), .CP(clk), 
        .Q(inner_first_stage_data_reg[1256]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1255_ ( .D(N9586), .CP(clk), 
        .Q(inner_first_stage_data_reg[1255]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1254_ ( .D(N9585), .CP(clk), 
        .Q(inner_first_stage_data_reg[1254]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1253_ ( .D(N9584), .CP(clk), 
        .Q(inner_first_stage_data_reg[1253]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1252_ ( .D(N9583), .CP(clk), 
        .Q(inner_first_stage_data_reg[1252]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1251_ ( .D(N9582), .CP(clk), 
        .Q(inner_first_stage_data_reg[1251]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1250_ ( .D(N9581), .CP(clk), 
        .Q(inner_first_stage_data_reg[1250]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1249_ ( .D(N9580), .CP(clk), 
        .Q(inner_first_stage_data_reg[1249]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1248_ ( .D(N9579), .CP(clk), 
        .Q(inner_first_stage_data_reg[1248]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_39_ ( .D(N9578), .CP(clk), 
        .Q(inner_first_stage_valid_reg[39]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1311_ ( .D(N9972), .CP(clk), 
        .Q(inner_first_stage_data_reg[1311]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1310_ ( .D(N9971), .CP(clk), 
        .Q(inner_first_stage_data_reg[1310]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1309_ ( .D(N9970), .CP(clk), 
        .Q(inner_first_stage_data_reg[1309]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1308_ ( .D(N9969), .CP(clk), 
        .Q(inner_first_stage_data_reg[1308]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1307_ ( .D(N9968), .CP(clk), 
        .Q(inner_first_stage_data_reg[1307]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1306_ ( .D(N9967), .CP(clk), 
        .Q(inner_first_stage_data_reg[1306]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1305_ ( .D(N9966), .CP(clk), 
        .Q(inner_first_stage_data_reg[1305]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1304_ ( .D(N9965), .CP(clk), 
        .Q(inner_first_stage_data_reg[1304]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1303_ ( .D(N9964), .CP(clk), 
        .Q(inner_first_stage_data_reg[1303]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1302_ ( .D(N9963), .CP(clk), 
        .Q(inner_first_stage_data_reg[1302]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1301_ ( .D(N9962), .CP(clk), 
        .Q(inner_first_stage_data_reg[1301]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1300_ ( .D(N9961), .CP(clk), 
        .Q(inner_first_stage_data_reg[1300]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1299_ ( .D(N9960), .CP(clk), 
        .Q(inner_first_stage_data_reg[1299]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1298_ ( .D(N9959), .CP(clk), 
        .Q(inner_first_stage_data_reg[1298]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1297_ ( .D(N9958), .CP(clk), 
        .Q(inner_first_stage_data_reg[1297]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1296_ ( .D(N9957), .CP(clk), 
        .Q(inner_first_stage_data_reg[1296]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1295_ ( .D(N9956), .CP(clk), 
        .Q(inner_first_stage_data_reg[1295]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1294_ ( .D(N9955), .CP(clk), 
        .Q(inner_first_stage_data_reg[1294]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1293_ ( .D(N9954), .CP(clk), 
        .Q(inner_first_stage_data_reg[1293]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1292_ ( .D(N9953), .CP(clk), 
        .Q(inner_first_stage_data_reg[1292]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1291_ ( .D(N9952), .CP(clk), 
        .Q(inner_first_stage_data_reg[1291]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1290_ ( .D(N9951), .CP(clk), 
        .Q(inner_first_stage_data_reg[1290]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1289_ ( .D(N9950), .CP(clk), 
        .Q(inner_first_stage_data_reg[1289]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1288_ ( .D(N9949), .CP(clk), 
        .Q(inner_first_stage_data_reg[1288]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1287_ ( .D(N9948), .CP(clk), 
        .Q(inner_first_stage_data_reg[1287]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1286_ ( .D(N9947), .CP(clk), 
        .Q(inner_first_stage_data_reg[1286]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1285_ ( .D(N9946), .CP(clk), 
        .Q(inner_first_stage_data_reg[1285]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1284_ ( .D(N9945), .CP(clk), 
        .Q(inner_first_stage_data_reg[1284]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1283_ ( .D(N9944), .CP(clk), 
        .Q(inner_first_stage_data_reg[1283]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1282_ ( .D(N9943), .CP(clk), 
        .Q(inner_first_stage_data_reg[1282]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1281_ ( .D(N9942), .CP(clk), 
        .Q(inner_first_stage_data_reg[1281]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1280_ ( .D(N9941), .CP(clk), 
        .Q(inner_first_stage_data_reg[1280]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_40_ ( .D(N9940), .CP(clk), 
        .Q(inner_first_stage_valid_reg[40]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1343_ ( .D(N10188), .CP(clk), .Q(inner_first_stage_data_reg[1343]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1342_ ( .D(N10187), .CP(clk), .Q(inner_first_stage_data_reg[1342]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1341_ ( .D(N10186), .CP(clk), .Q(inner_first_stage_data_reg[1341]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1340_ ( .D(N10185), .CP(clk), .Q(inner_first_stage_data_reg[1340]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1339_ ( .D(N10184), .CP(clk), .Q(inner_first_stage_data_reg[1339]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1338_ ( .D(N10183), .CP(clk), .Q(inner_first_stage_data_reg[1338]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1337_ ( .D(N10182), .CP(clk), .Q(inner_first_stage_data_reg[1337]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1336_ ( .D(N10181), .CP(clk), .Q(inner_first_stage_data_reg[1336]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1335_ ( .D(N10180), .CP(clk), .Q(inner_first_stage_data_reg[1335]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1334_ ( .D(N10179), .CP(clk), .Q(inner_first_stage_data_reg[1334]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1333_ ( .D(N10178), .CP(clk), .Q(inner_first_stage_data_reg[1333]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1332_ ( .D(N10177), .CP(clk), .Q(inner_first_stage_data_reg[1332]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1331_ ( .D(N10176), .CP(clk), .Q(inner_first_stage_data_reg[1331]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1330_ ( .D(N10175), .CP(clk), .Q(inner_first_stage_data_reg[1330]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1329_ ( .D(N10174), .CP(clk), .Q(inner_first_stage_data_reg[1329]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1328_ ( .D(N10173), .CP(clk), .Q(inner_first_stage_data_reg[1328]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1327_ ( .D(N10172), .CP(clk), .Q(inner_first_stage_data_reg[1327]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1326_ ( .D(N10171), .CP(clk), .Q(inner_first_stage_data_reg[1326]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1325_ ( .D(N10170), .CP(clk), .Q(inner_first_stage_data_reg[1325]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1324_ ( .D(N10169), .CP(clk), .Q(inner_first_stage_data_reg[1324]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1323_ ( .D(N10168), .CP(clk), .Q(inner_first_stage_data_reg[1323]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1322_ ( .D(N10167), .CP(clk), .Q(inner_first_stage_data_reg[1322]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1321_ ( .D(N10166), .CP(clk), .Q(inner_first_stage_data_reg[1321]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1320_ ( .D(N10165), .CP(clk), .Q(inner_first_stage_data_reg[1320]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1319_ ( .D(N10164), .CP(clk), .Q(inner_first_stage_data_reg[1319]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1318_ ( .D(N10163), .CP(clk), .Q(inner_first_stage_data_reg[1318]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1317_ ( .D(N10162), .CP(clk), .Q(inner_first_stage_data_reg[1317]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1316_ ( .D(N10161), .CP(clk), .Q(inner_first_stage_data_reg[1316]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1315_ ( .D(N10160), .CP(clk), .Q(inner_first_stage_data_reg[1315]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1314_ ( .D(N10159), .CP(clk), .Q(inner_first_stage_data_reg[1314]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1313_ ( .D(N10158), .CP(clk), .Q(inner_first_stage_data_reg[1313]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1312_ ( .D(N10157), .CP(clk), .Q(inner_first_stage_data_reg[1312]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_41_ ( .D(N10156), .CP(clk), 
        .Q(inner_first_stage_valid_reg[41]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1375_ ( .D(N10404), .CP(clk), .Q(inner_first_stage_data_reg[1375]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1374_ ( .D(N10403), .CP(clk), .Q(inner_first_stage_data_reg[1374]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1373_ ( .D(N10402), .CP(clk), .Q(inner_first_stage_data_reg[1373]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1372_ ( .D(N10401), .CP(clk), .Q(inner_first_stage_data_reg[1372]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1371_ ( .D(N10400), .CP(clk), .Q(inner_first_stage_data_reg[1371]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1370_ ( .D(N10399), .CP(clk), .Q(inner_first_stage_data_reg[1370]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1369_ ( .D(N10398), .CP(clk), .Q(inner_first_stage_data_reg[1369]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1368_ ( .D(N10397), .CP(clk), .Q(inner_first_stage_data_reg[1368]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1367_ ( .D(N10396), .CP(clk), .Q(inner_first_stage_data_reg[1367]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1366_ ( .D(N10395), .CP(clk), .Q(inner_first_stage_data_reg[1366]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1365_ ( .D(N10394), .CP(clk), .Q(inner_first_stage_data_reg[1365]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1364_ ( .D(N10393), .CP(clk), .Q(inner_first_stage_data_reg[1364]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1363_ ( .D(N10392), .CP(clk), .Q(inner_first_stage_data_reg[1363]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1362_ ( .D(N10391), .CP(clk), .Q(inner_first_stage_data_reg[1362]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1361_ ( .D(N10390), .CP(clk), .Q(inner_first_stage_data_reg[1361]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1360_ ( .D(N10389), .CP(clk), .Q(inner_first_stage_data_reg[1360]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1359_ ( .D(N10388), .CP(clk), .Q(inner_first_stage_data_reg[1359]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1358_ ( .D(N10387), .CP(clk), .Q(inner_first_stage_data_reg[1358]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1357_ ( .D(N10386), .CP(clk), .Q(inner_first_stage_data_reg[1357]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1356_ ( .D(N10385), .CP(clk), .Q(inner_first_stage_data_reg[1356]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1355_ ( .D(N10384), .CP(clk), .Q(inner_first_stage_data_reg[1355]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1354_ ( .D(N10383), .CP(clk), .Q(inner_first_stage_data_reg[1354]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1353_ ( .D(N10382), .CP(clk), .Q(inner_first_stage_data_reg[1353]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1352_ ( .D(N10381), .CP(clk), .Q(inner_first_stage_data_reg[1352]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1351_ ( .D(N10380), .CP(clk), .Q(inner_first_stage_data_reg[1351]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1350_ ( .D(N10379), .CP(clk), .Q(inner_first_stage_data_reg[1350]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1349_ ( .D(N10378), .CP(clk), .Q(inner_first_stage_data_reg[1349]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1348_ ( .D(N10377), .CP(clk), .Q(inner_first_stage_data_reg[1348]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1347_ ( .D(N10376), .CP(clk), .Q(inner_first_stage_data_reg[1347]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1346_ ( .D(N10375), .CP(clk), .Q(inner_first_stage_data_reg[1346]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1345_ ( .D(N10374), .CP(clk), .Q(inner_first_stage_data_reg[1345]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1344_ ( .D(N10373), .CP(clk), .Q(inner_first_stage_data_reg[1344]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_42_ ( .D(N10372), .CP(clk), 
        .Q(inner_first_stage_valid_reg[42]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1407_ ( .D(N10620), .CP(clk), .Q(inner_first_stage_data_reg[1407]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1406_ ( .D(N10619), .CP(clk), .Q(inner_first_stage_data_reg[1406]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1405_ ( .D(N10618), .CP(clk), .Q(inner_first_stage_data_reg[1405]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1404_ ( .D(N10617), .CP(clk), .Q(inner_first_stage_data_reg[1404]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1403_ ( .D(N10616), .CP(clk), .Q(inner_first_stage_data_reg[1403]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1402_ ( .D(N10615), .CP(clk), .Q(inner_first_stage_data_reg[1402]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1401_ ( .D(N10614), .CP(clk), .Q(inner_first_stage_data_reg[1401]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1400_ ( .D(N10613), .CP(clk), .Q(inner_first_stage_data_reg[1400]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1399_ ( .D(N10612), .CP(clk), .Q(inner_first_stage_data_reg[1399]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1398_ ( .D(N10611), .CP(clk), .Q(inner_first_stage_data_reg[1398]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1397_ ( .D(N10610), .CP(clk), .Q(inner_first_stage_data_reg[1397]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1396_ ( .D(N10609), .CP(clk), .Q(inner_first_stage_data_reg[1396]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1395_ ( .D(N10608), .CP(clk), .Q(inner_first_stage_data_reg[1395]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1394_ ( .D(N10607), .CP(clk), .Q(inner_first_stage_data_reg[1394]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1393_ ( .D(N10606), .CP(clk), .Q(inner_first_stage_data_reg[1393]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1392_ ( .D(N10605), .CP(clk), .Q(inner_first_stage_data_reg[1392]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1391_ ( .D(N10604), .CP(clk), .Q(inner_first_stage_data_reg[1391]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1390_ ( .D(N10603), .CP(clk), .Q(inner_first_stage_data_reg[1390]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1389_ ( .D(N10602), .CP(clk), .Q(inner_first_stage_data_reg[1389]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1388_ ( .D(N10601), .CP(clk), .Q(inner_first_stage_data_reg[1388]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1387_ ( .D(N10600), .CP(clk), .Q(inner_first_stage_data_reg[1387]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1386_ ( .D(N10599), .CP(clk), .Q(inner_first_stage_data_reg[1386]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1385_ ( .D(N10598), .CP(clk), .Q(inner_first_stage_data_reg[1385]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1384_ ( .D(N10597), .CP(clk), .Q(inner_first_stage_data_reg[1384]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1383_ ( .D(N10596), .CP(clk), .Q(inner_first_stage_data_reg[1383]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1382_ ( .D(N10595), .CP(clk), .Q(inner_first_stage_data_reg[1382]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1381_ ( .D(N10594), .CP(clk), .Q(inner_first_stage_data_reg[1381]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1380_ ( .D(N10593), .CP(clk), .Q(inner_first_stage_data_reg[1380]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1379_ ( .D(N10592), .CP(clk), .Q(inner_first_stage_data_reg[1379]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1378_ ( .D(N10591), .CP(clk), .Q(inner_first_stage_data_reg[1378]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1377_ ( .D(N10590), .CP(clk), .Q(inner_first_stage_data_reg[1377]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1376_ ( .D(N10589), .CP(clk), .Q(inner_first_stage_data_reg[1376]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_43_ ( .D(N10588), .CP(clk), 
        .Q(inner_first_stage_valid_reg[43]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1439_ ( .D(N10836), .CP(clk), .Q(inner_first_stage_data_reg[1439]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1438_ ( .D(N10835), .CP(clk), .Q(inner_first_stage_data_reg[1438]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1437_ ( .D(N10834), .CP(clk), .Q(inner_first_stage_data_reg[1437]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1436_ ( .D(N10833), .CP(clk), .Q(inner_first_stage_data_reg[1436]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1435_ ( .D(N10832), .CP(clk), .Q(inner_first_stage_data_reg[1435]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1434_ ( .D(N10831), .CP(clk), .Q(inner_first_stage_data_reg[1434]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1433_ ( .D(N10830), .CP(clk), .Q(inner_first_stage_data_reg[1433]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1432_ ( .D(N10829), .CP(clk), .Q(inner_first_stage_data_reg[1432]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1431_ ( .D(N10828), .CP(clk), .Q(inner_first_stage_data_reg[1431]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1430_ ( .D(N10827), .CP(clk), .Q(inner_first_stage_data_reg[1430]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1429_ ( .D(N10826), .CP(clk), .Q(inner_first_stage_data_reg[1429]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1428_ ( .D(N10825), .CP(clk), .Q(inner_first_stage_data_reg[1428]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1427_ ( .D(N10824), .CP(clk), .Q(inner_first_stage_data_reg[1427]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1426_ ( .D(N10823), .CP(clk), .Q(inner_first_stage_data_reg[1426]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1425_ ( .D(N10822), .CP(clk), .Q(inner_first_stage_data_reg[1425]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1424_ ( .D(N10821), .CP(clk), .Q(inner_first_stage_data_reg[1424]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1423_ ( .D(N10820), .CP(clk), .Q(inner_first_stage_data_reg[1423]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1422_ ( .D(N10819), .CP(clk), .Q(inner_first_stage_data_reg[1422]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1421_ ( .D(N10818), .CP(clk), .Q(inner_first_stage_data_reg[1421]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1420_ ( .D(N10817), .CP(clk), .Q(inner_first_stage_data_reg[1420]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1419_ ( .D(N10816), .CP(clk), .Q(inner_first_stage_data_reg[1419]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1418_ ( .D(N10815), .CP(clk), .Q(inner_first_stage_data_reg[1418]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1417_ ( .D(N10814), .CP(clk), .Q(inner_first_stage_data_reg[1417]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1416_ ( .D(N10813), .CP(clk), .Q(inner_first_stage_data_reg[1416]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1415_ ( .D(N10812), .CP(clk), .Q(inner_first_stage_data_reg[1415]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1414_ ( .D(N10811), .CP(clk), .Q(inner_first_stage_data_reg[1414]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1413_ ( .D(N10810), .CP(clk), .Q(inner_first_stage_data_reg[1413]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1412_ ( .D(N10809), .CP(clk), .Q(inner_first_stage_data_reg[1412]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1411_ ( .D(N10808), .CP(clk), .Q(inner_first_stage_data_reg[1411]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1410_ ( .D(N10807), .CP(clk), .Q(inner_first_stage_data_reg[1410]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1409_ ( .D(N10806), .CP(clk), .Q(inner_first_stage_data_reg[1409]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1408_ ( .D(N10805), .CP(clk), .Q(inner_first_stage_data_reg[1408]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_44_ ( .D(N10804), .CP(clk), 
        .Q(inner_first_stage_valid_reg[44]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1471_ ( .D(N11052), .CP(clk), .Q(inner_first_stage_data_reg[1471]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1470_ ( .D(N11051), .CP(clk), .Q(inner_first_stage_data_reg[1470]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1469_ ( .D(N11050), .CP(clk), .Q(inner_first_stage_data_reg[1469]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1468_ ( .D(N11049), .CP(clk), .Q(inner_first_stage_data_reg[1468]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1467_ ( .D(N11048), .CP(clk), .Q(inner_first_stage_data_reg[1467]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1466_ ( .D(N11047), .CP(clk), .Q(inner_first_stage_data_reg[1466]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1465_ ( .D(N11046), .CP(clk), .Q(inner_first_stage_data_reg[1465]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1464_ ( .D(N11045), .CP(clk), .Q(inner_first_stage_data_reg[1464]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1463_ ( .D(N11044), .CP(clk), .Q(inner_first_stage_data_reg[1463]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1462_ ( .D(N11043), .CP(clk), .Q(inner_first_stage_data_reg[1462]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1461_ ( .D(N11042), .CP(clk), .Q(inner_first_stage_data_reg[1461]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1460_ ( .D(N11041), .CP(clk), .Q(inner_first_stage_data_reg[1460]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1459_ ( .D(N11040), .CP(clk), .Q(inner_first_stage_data_reg[1459]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1458_ ( .D(N11039), .CP(clk), .Q(inner_first_stage_data_reg[1458]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1457_ ( .D(N11038), .CP(clk), .Q(inner_first_stage_data_reg[1457]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1456_ ( .D(N11037), .CP(clk), .Q(inner_first_stage_data_reg[1456]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1455_ ( .D(N11036), .CP(clk), .Q(inner_first_stage_data_reg[1455]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1454_ ( .D(N11035), .CP(clk), .Q(inner_first_stage_data_reg[1454]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1453_ ( .D(N11034), .CP(clk), .Q(inner_first_stage_data_reg[1453]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1452_ ( .D(N11033), .CP(clk), .Q(inner_first_stage_data_reg[1452]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1451_ ( .D(N11032), .CP(clk), .Q(inner_first_stage_data_reg[1451]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1450_ ( .D(N11031), .CP(clk), .Q(inner_first_stage_data_reg[1450]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1449_ ( .D(N11030), .CP(clk), .Q(inner_first_stage_data_reg[1449]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1448_ ( .D(N11029), .CP(clk), .Q(inner_first_stage_data_reg[1448]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1447_ ( .D(N11028), .CP(clk), .Q(inner_first_stage_data_reg[1447]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1446_ ( .D(N11027), .CP(clk), .Q(inner_first_stage_data_reg[1446]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1445_ ( .D(N11026), .CP(clk), .Q(inner_first_stage_data_reg[1445]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1444_ ( .D(N11025), .CP(clk), .Q(inner_first_stage_data_reg[1444]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1443_ ( .D(N11024), .CP(clk), .Q(inner_first_stage_data_reg[1443]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1442_ ( .D(N11023), .CP(clk), .Q(inner_first_stage_data_reg[1442]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1441_ ( .D(N11022), .CP(clk), .Q(inner_first_stage_data_reg[1441]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1440_ ( .D(N11021), .CP(clk), .Q(inner_first_stage_data_reg[1440]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_45_ ( .D(N11020), .CP(clk), 
        .Q(inner_first_stage_valid_reg[45]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1503_ ( .D(N11268), .CP(clk), .Q(inner_first_stage_data_reg[1503]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1502_ ( .D(N11267), .CP(clk), .Q(inner_first_stage_data_reg[1502]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1501_ ( .D(N11266), .CP(clk), .Q(inner_first_stage_data_reg[1501]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1500_ ( .D(N11265), .CP(clk), .Q(inner_first_stage_data_reg[1500]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1499_ ( .D(N11264), .CP(clk), .Q(inner_first_stage_data_reg[1499]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1498_ ( .D(N11263), .CP(clk), .Q(inner_first_stage_data_reg[1498]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1497_ ( .D(N11262), .CP(clk), .Q(inner_first_stage_data_reg[1497]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1496_ ( .D(N11261), .CP(clk), .Q(inner_first_stage_data_reg[1496]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1495_ ( .D(N11260), .CP(clk), .Q(inner_first_stage_data_reg[1495]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1494_ ( .D(N11259), .CP(clk), .Q(inner_first_stage_data_reg[1494]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1493_ ( .D(N11258), .CP(clk), .Q(inner_first_stage_data_reg[1493]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1492_ ( .D(N11257), .CP(clk), .Q(inner_first_stage_data_reg[1492]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1491_ ( .D(N11256), .CP(clk), .Q(inner_first_stage_data_reg[1491]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1490_ ( .D(N11255), .CP(clk), .Q(inner_first_stage_data_reg[1490]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1489_ ( .D(N11254), .CP(clk), .Q(inner_first_stage_data_reg[1489]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1488_ ( .D(N11253), .CP(clk), .Q(inner_first_stage_data_reg[1488]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1487_ ( .D(N11252), .CP(clk), .Q(inner_first_stage_data_reg[1487]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1486_ ( .D(N11251), .CP(clk), .Q(inner_first_stage_data_reg[1486]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1485_ ( .D(N11250), .CP(clk), .Q(inner_first_stage_data_reg[1485]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1484_ ( .D(N11249), .CP(clk), .Q(inner_first_stage_data_reg[1484]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1483_ ( .D(N11248), .CP(clk), .Q(inner_first_stage_data_reg[1483]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1482_ ( .D(N11247), .CP(clk), .Q(inner_first_stage_data_reg[1482]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1481_ ( .D(N11246), .CP(clk), .Q(inner_first_stage_data_reg[1481]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1480_ ( .D(N11245), .CP(clk), .Q(inner_first_stage_data_reg[1480]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1479_ ( .D(N11244), .CP(clk), .Q(inner_first_stage_data_reg[1479]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1478_ ( .D(N11243), .CP(clk), .Q(inner_first_stage_data_reg[1478]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1477_ ( .D(N11242), .CP(clk), .Q(inner_first_stage_data_reg[1477]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1476_ ( .D(N11241), .CP(clk), .Q(inner_first_stage_data_reg[1476]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1475_ ( .D(N11240), .CP(clk), .Q(inner_first_stage_data_reg[1475]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1474_ ( .D(N11239), .CP(clk), .Q(inner_first_stage_data_reg[1474]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1473_ ( .D(N11238), .CP(clk), .Q(inner_first_stage_data_reg[1473]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1472_ ( .D(N11237), .CP(clk), .Q(inner_first_stage_data_reg[1472]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_46_ ( .D(N11236), .CP(clk), 
        .Q(inner_first_stage_valid_reg[46]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1535_ ( .D(N11484), .CP(clk), .Q(inner_first_stage_data_reg[1535]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1534_ ( .D(N11483), .CP(clk), .Q(inner_first_stage_data_reg[1534]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1533_ ( .D(N11482), .CP(clk), .Q(inner_first_stage_data_reg[1533]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1532_ ( .D(N11481), .CP(clk), .Q(inner_first_stage_data_reg[1532]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1531_ ( .D(N11480), .CP(clk), .Q(inner_first_stage_data_reg[1531]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1530_ ( .D(N11479), .CP(clk), .Q(inner_first_stage_data_reg[1530]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1529_ ( .D(N11478), .CP(clk), .Q(inner_first_stage_data_reg[1529]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1528_ ( .D(N11477), .CP(clk), .Q(inner_first_stage_data_reg[1528]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1527_ ( .D(N11476), .CP(clk), .Q(inner_first_stage_data_reg[1527]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1526_ ( .D(N11475), .CP(clk), .Q(inner_first_stage_data_reg[1526]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1525_ ( .D(N11474), .CP(clk), .Q(inner_first_stage_data_reg[1525]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1524_ ( .D(N11473), .CP(clk), .Q(inner_first_stage_data_reg[1524]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1523_ ( .D(N11472), .CP(clk), .Q(inner_first_stage_data_reg[1523]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1522_ ( .D(N11471), .CP(clk), .Q(inner_first_stage_data_reg[1522]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1521_ ( .D(N11470), .CP(clk), .Q(inner_first_stage_data_reg[1521]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1520_ ( .D(N11469), .CP(clk), .Q(inner_first_stage_data_reg[1520]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1519_ ( .D(N11468), .CP(clk), .Q(inner_first_stage_data_reg[1519]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1518_ ( .D(N11467), .CP(clk), .Q(inner_first_stage_data_reg[1518]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1517_ ( .D(N11466), .CP(clk), .Q(inner_first_stage_data_reg[1517]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1516_ ( .D(N11465), .CP(clk), .Q(inner_first_stage_data_reg[1516]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1515_ ( .D(N11464), .CP(clk), .Q(inner_first_stage_data_reg[1515]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1514_ ( .D(N11463), .CP(clk), .Q(inner_first_stage_data_reg[1514]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1513_ ( .D(N11462), .CP(clk), .Q(inner_first_stage_data_reg[1513]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1512_ ( .D(N11461), .CP(clk), .Q(inner_first_stage_data_reg[1512]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1511_ ( .D(N11460), .CP(clk), .Q(inner_first_stage_data_reg[1511]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1510_ ( .D(N11459), .CP(clk), .Q(inner_first_stage_data_reg[1510]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1509_ ( .D(N11458), .CP(clk), .Q(inner_first_stage_data_reg[1509]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1508_ ( .D(N11457), .CP(clk), .Q(inner_first_stage_data_reg[1508]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1507_ ( .D(N11456), .CP(clk), .Q(inner_first_stage_data_reg[1507]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1506_ ( .D(N11455), .CP(clk), .Q(inner_first_stage_data_reg[1506]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1505_ ( .D(N11454), .CP(clk), .Q(inner_first_stage_data_reg[1505]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1504_ ( .D(N11453), .CP(clk), .Q(inner_first_stage_data_reg[1504]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_47_ ( .D(N11452), .CP(clk), 
        .Q(inner_first_stage_valid_reg[47]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1567_ ( .D(N11846), .CP(clk), .Q(inner_first_stage_data_reg[1567]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1566_ ( .D(N11845), .CP(clk), .Q(inner_first_stage_data_reg[1566]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1565_ ( .D(N11844), .CP(clk), .Q(inner_first_stage_data_reg[1565]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1564_ ( .D(N11843), .CP(clk), .Q(inner_first_stage_data_reg[1564]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1563_ ( .D(N11842), .CP(clk), .Q(inner_first_stage_data_reg[1563]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1562_ ( .D(N11841), .CP(clk), .Q(inner_first_stage_data_reg[1562]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1561_ ( .D(N11840), .CP(clk), .Q(inner_first_stage_data_reg[1561]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1560_ ( .D(N11839), .CP(clk), .Q(inner_first_stage_data_reg[1560]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1559_ ( .D(N11838), .CP(clk), .Q(inner_first_stage_data_reg[1559]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1558_ ( .D(N11837), .CP(clk), .Q(inner_first_stage_data_reg[1558]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1557_ ( .D(N11836), .CP(clk), .Q(inner_first_stage_data_reg[1557]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1556_ ( .D(N11835), .CP(clk), .Q(inner_first_stage_data_reg[1556]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1555_ ( .D(N11834), .CP(clk), .Q(inner_first_stage_data_reg[1555]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1554_ ( .D(N11833), .CP(clk), .Q(inner_first_stage_data_reg[1554]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1553_ ( .D(N11832), .CP(clk), .Q(inner_first_stage_data_reg[1553]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1552_ ( .D(N11831), .CP(clk), .Q(inner_first_stage_data_reg[1552]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1551_ ( .D(N11830), .CP(clk), .Q(inner_first_stage_data_reg[1551]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1550_ ( .D(N11829), .CP(clk), .Q(inner_first_stage_data_reg[1550]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1549_ ( .D(N11828), .CP(clk), .Q(inner_first_stage_data_reg[1549]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1548_ ( .D(N11827), .CP(clk), .Q(inner_first_stage_data_reg[1548]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1547_ ( .D(N11826), .CP(clk), .Q(inner_first_stage_data_reg[1547]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1546_ ( .D(N11825), .CP(clk), .Q(inner_first_stage_data_reg[1546]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1545_ ( .D(N11824), .CP(clk), .Q(inner_first_stage_data_reg[1545]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1544_ ( .D(N11823), .CP(clk), .Q(inner_first_stage_data_reg[1544]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1543_ ( .D(N11822), .CP(clk), .Q(inner_first_stage_data_reg[1543]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1542_ ( .D(N11821), .CP(clk), .Q(inner_first_stage_data_reg[1542]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1541_ ( .D(N11820), .CP(clk), .Q(inner_first_stage_data_reg[1541]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1540_ ( .D(N11819), .CP(clk), .Q(inner_first_stage_data_reg[1540]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1539_ ( .D(N11818), .CP(clk), .Q(inner_first_stage_data_reg[1539]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1538_ ( .D(N11817), .CP(clk), .Q(inner_first_stage_data_reg[1538]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1537_ ( .D(N11816), .CP(clk), .Q(inner_first_stage_data_reg[1537]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1536_ ( .D(N11815), .CP(clk), .Q(inner_first_stage_data_reg[1536]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_48_ ( .D(N11814), .CP(clk), 
        .Q(inner_first_stage_valid_reg[48]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1599_ ( .D(N12062), .CP(clk), .Q(inner_first_stage_data_reg[1599]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1598_ ( .D(N12061), .CP(clk), .Q(inner_first_stage_data_reg[1598]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1597_ ( .D(N12060), .CP(clk), .Q(inner_first_stage_data_reg[1597]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1596_ ( .D(N12059), .CP(clk), .Q(inner_first_stage_data_reg[1596]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1595_ ( .D(N12058), .CP(clk), .Q(inner_first_stage_data_reg[1595]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1594_ ( .D(N12057), .CP(clk), .Q(inner_first_stage_data_reg[1594]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1593_ ( .D(N12056), .CP(clk), .Q(inner_first_stage_data_reg[1593]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1592_ ( .D(N12055), .CP(clk), .Q(inner_first_stage_data_reg[1592]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1591_ ( .D(N12054), .CP(clk), .Q(inner_first_stage_data_reg[1591]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1590_ ( .D(N12053), .CP(clk), .Q(inner_first_stage_data_reg[1590]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1589_ ( .D(N12052), .CP(clk), .Q(inner_first_stage_data_reg[1589]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1588_ ( .D(N12051), .CP(clk), .Q(inner_first_stage_data_reg[1588]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1587_ ( .D(N12050), .CP(clk), .Q(inner_first_stage_data_reg[1587]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1586_ ( .D(N12049), .CP(clk), .Q(inner_first_stage_data_reg[1586]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1585_ ( .D(N12048), .CP(clk), .Q(inner_first_stage_data_reg[1585]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1584_ ( .D(N12047), .CP(clk), .Q(inner_first_stage_data_reg[1584]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1583_ ( .D(N12046), .CP(clk), .Q(inner_first_stage_data_reg[1583]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1582_ ( .D(N12045), .CP(clk), .Q(inner_first_stage_data_reg[1582]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1581_ ( .D(N12044), .CP(clk), .Q(inner_first_stage_data_reg[1581]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1580_ ( .D(N12043), .CP(clk), .Q(inner_first_stage_data_reg[1580]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1579_ ( .D(N12042), .CP(clk), .Q(inner_first_stage_data_reg[1579]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1578_ ( .D(N12041), .CP(clk), .Q(inner_first_stage_data_reg[1578]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1577_ ( .D(N12040), .CP(clk), .Q(inner_first_stage_data_reg[1577]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1576_ ( .D(N12039), .CP(clk), .Q(inner_first_stage_data_reg[1576]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1575_ ( .D(N12038), .CP(clk), .Q(inner_first_stage_data_reg[1575]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1574_ ( .D(N12037), .CP(clk), .Q(inner_first_stage_data_reg[1574]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1573_ ( .D(N12036), .CP(clk), .Q(inner_first_stage_data_reg[1573]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1572_ ( .D(N12035), .CP(clk), .Q(inner_first_stage_data_reg[1572]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1571_ ( .D(N12034), .CP(clk), .Q(inner_first_stage_data_reg[1571]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1570_ ( .D(N12033), .CP(clk), .Q(inner_first_stage_data_reg[1570]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1569_ ( .D(N12032), .CP(clk), .Q(inner_first_stage_data_reg[1569]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1568_ ( .D(N12031), .CP(clk), .Q(inner_first_stage_data_reg[1568]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_49_ ( .D(N12030), .CP(clk), 
        .Q(inner_first_stage_valid_reg[49]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1631_ ( .D(N12278), .CP(clk), .Q(inner_first_stage_data_reg[1631]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1630_ ( .D(N12277), .CP(clk), .Q(inner_first_stage_data_reg[1630]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1629_ ( .D(N12276), .CP(clk), .Q(inner_first_stage_data_reg[1629]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1628_ ( .D(N12275), .CP(clk), .Q(inner_first_stage_data_reg[1628]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1627_ ( .D(N12274), .CP(clk), .Q(inner_first_stage_data_reg[1627]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1626_ ( .D(N12273), .CP(clk), .Q(inner_first_stage_data_reg[1626]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1625_ ( .D(N12272), .CP(clk), .Q(inner_first_stage_data_reg[1625]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1624_ ( .D(N12271), .CP(clk), .Q(inner_first_stage_data_reg[1624]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1623_ ( .D(N12270), .CP(clk), .Q(inner_first_stage_data_reg[1623]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1622_ ( .D(N12269), .CP(clk), .Q(inner_first_stage_data_reg[1622]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1621_ ( .D(N12268), .CP(clk), .Q(inner_first_stage_data_reg[1621]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1620_ ( .D(N12267), .CP(clk), .Q(inner_first_stage_data_reg[1620]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1619_ ( .D(N12266), .CP(clk), .Q(inner_first_stage_data_reg[1619]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1618_ ( .D(N12265), .CP(clk), .Q(inner_first_stage_data_reg[1618]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1617_ ( .D(N12264), .CP(clk), .Q(inner_first_stage_data_reg[1617]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1616_ ( .D(N12263), .CP(clk), .Q(inner_first_stage_data_reg[1616]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1615_ ( .D(N12262), .CP(clk), .Q(inner_first_stage_data_reg[1615]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1614_ ( .D(N12261), .CP(clk), .Q(inner_first_stage_data_reg[1614]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1613_ ( .D(N12260), .CP(clk), .Q(inner_first_stage_data_reg[1613]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1612_ ( .D(N12259), .CP(clk), .Q(inner_first_stage_data_reg[1612]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1611_ ( .D(N12258), .CP(clk), .Q(inner_first_stage_data_reg[1611]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1610_ ( .D(N12257), .CP(clk), .Q(inner_first_stage_data_reg[1610]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1609_ ( .D(N12256), .CP(clk), .Q(inner_first_stage_data_reg[1609]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1608_ ( .D(N12255), .CP(clk), .Q(inner_first_stage_data_reg[1608]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1607_ ( .D(N12254), .CP(clk), .Q(inner_first_stage_data_reg[1607]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1606_ ( .D(N12253), .CP(clk), .Q(inner_first_stage_data_reg[1606]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1605_ ( .D(N12252), .CP(clk), .Q(inner_first_stage_data_reg[1605]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1604_ ( .D(N12251), .CP(clk), .Q(inner_first_stage_data_reg[1604]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1603_ ( .D(N12250), .CP(clk), .Q(inner_first_stage_data_reg[1603]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1602_ ( .D(N12249), .CP(clk), .Q(inner_first_stage_data_reg[1602]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1601_ ( .D(N12248), .CP(clk), .Q(inner_first_stage_data_reg[1601]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1600_ ( .D(N12247), .CP(clk), .Q(inner_first_stage_data_reg[1600]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_50_ ( .D(N12246), .CP(clk), 
        .Q(inner_first_stage_valid_reg[50]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1663_ ( .D(N12494), .CP(clk), .Q(inner_first_stage_data_reg[1663]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1662_ ( .D(N12493), .CP(clk), .Q(inner_first_stage_data_reg[1662]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1661_ ( .D(N12492), .CP(clk), .Q(inner_first_stage_data_reg[1661]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1660_ ( .D(N12491), .CP(clk), .Q(inner_first_stage_data_reg[1660]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1659_ ( .D(N12490), .CP(clk), .Q(inner_first_stage_data_reg[1659]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1658_ ( .D(N12489), .CP(clk), .Q(inner_first_stage_data_reg[1658]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1657_ ( .D(N12488), .CP(clk), .Q(inner_first_stage_data_reg[1657]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1656_ ( .D(N12487), .CP(clk), .Q(inner_first_stage_data_reg[1656]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1655_ ( .D(N12486), .CP(clk), .Q(inner_first_stage_data_reg[1655]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1654_ ( .D(N12485), .CP(clk), .Q(inner_first_stage_data_reg[1654]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1653_ ( .D(N12484), .CP(clk), .Q(inner_first_stage_data_reg[1653]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1652_ ( .D(N12483), .CP(clk), .Q(inner_first_stage_data_reg[1652]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1651_ ( .D(N12482), .CP(clk), .Q(inner_first_stage_data_reg[1651]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1650_ ( .D(N12481), .CP(clk), .Q(inner_first_stage_data_reg[1650]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1649_ ( .D(N12480), .CP(clk), .Q(inner_first_stage_data_reg[1649]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1648_ ( .D(N12479), .CP(clk), .Q(inner_first_stage_data_reg[1648]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1647_ ( .D(N12478), .CP(clk), .Q(inner_first_stage_data_reg[1647]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1646_ ( .D(N12477), .CP(clk), .Q(inner_first_stage_data_reg[1646]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1645_ ( .D(N12476), .CP(clk), .Q(inner_first_stage_data_reg[1645]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1644_ ( .D(N12475), .CP(clk), .Q(inner_first_stage_data_reg[1644]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1643_ ( .D(N12474), .CP(clk), .Q(inner_first_stage_data_reg[1643]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1642_ ( .D(N12473), .CP(clk), .Q(inner_first_stage_data_reg[1642]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1641_ ( .D(N12472), .CP(clk), .Q(inner_first_stage_data_reg[1641]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1640_ ( .D(N12471), .CP(clk), .Q(inner_first_stage_data_reg[1640]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1639_ ( .D(N12470), .CP(clk), .Q(inner_first_stage_data_reg[1639]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1638_ ( .D(N12469), .CP(clk), .Q(inner_first_stage_data_reg[1638]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1637_ ( .D(N12468), .CP(clk), .Q(inner_first_stage_data_reg[1637]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1636_ ( .D(N12467), .CP(clk), .Q(inner_first_stage_data_reg[1636]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1635_ ( .D(N12466), .CP(clk), .Q(inner_first_stage_data_reg[1635]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1634_ ( .D(N12465), .CP(clk), .Q(inner_first_stage_data_reg[1634]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1633_ ( .D(N12464), .CP(clk), .Q(inner_first_stage_data_reg[1633]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1632_ ( .D(N12463), .CP(clk), .Q(inner_first_stage_data_reg[1632]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_51_ ( .D(N12462), .CP(clk), 
        .Q(inner_first_stage_valid_reg[51]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1695_ ( .D(N12710), .CP(clk), .Q(inner_first_stage_data_reg[1695]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1694_ ( .D(N12709), .CP(clk), .Q(inner_first_stage_data_reg[1694]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1693_ ( .D(N12708), .CP(clk), .Q(inner_first_stage_data_reg[1693]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1692_ ( .D(N12707), .CP(clk), .Q(inner_first_stage_data_reg[1692]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1691_ ( .D(N12706), .CP(clk), .Q(inner_first_stage_data_reg[1691]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1690_ ( .D(N12705), .CP(clk), .Q(inner_first_stage_data_reg[1690]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1689_ ( .D(N12704), .CP(clk), .Q(inner_first_stage_data_reg[1689]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1688_ ( .D(N12703), .CP(clk), .Q(inner_first_stage_data_reg[1688]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1687_ ( .D(N12702), .CP(clk), .Q(inner_first_stage_data_reg[1687]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1686_ ( .D(N12701), .CP(clk), .Q(inner_first_stage_data_reg[1686]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1685_ ( .D(N12700), .CP(clk), .Q(inner_first_stage_data_reg[1685]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1684_ ( .D(N12699), .CP(clk), .Q(inner_first_stage_data_reg[1684]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1683_ ( .D(N12698), .CP(clk), .Q(inner_first_stage_data_reg[1683]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1682_ ( .D(N12697), .CP(clk), .Q(inner_first_stage_data_reg[1682]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1681_ ( .D(N12696), .CP(clk), .Q(inner_first_stage_data_reg[1681]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1680_ ( .D(N12695), .CP(clk), .Q(inner_first_stage_data_reg[1680]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1679_ ( .D(N12694), .CP(clk), .Q(inner_first_stage_data_reg[1679]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1678_ ( .D(N12693), .CP(clk), .Q(inner_first_stage_data_reg[1678]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1677_ ( .D(N12692), .CP(clk), .Q(inner_first_stage_data_reg[1677]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1676_ ( .D(N12691), .CP(clk), .Q(inner_first_stage_data_reg[1676]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1675_ ( .D(N12690), .CP(clk), .Q(inner_first_stage_data_reg[1675]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1674_ ( .D(N12689), .CP(clk), .Q(inner_first_stage_data_reg[1674]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1673_ ( .D(N12688), .CP(clk), .Q(inner_first_stage_data_reg[1673]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1672_ ( .D(N12687), .CP(clk), .Q(inner_first_stage_data_reg[1672]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1671_ ( .D(N12686), .CP(clk), .Q(inner_first_stage_data_reg[1671]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1670_ ( .D(N12685), .CP(clk), .Q(inner_first_stage_data_reg[1670]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1669_ ( .D(N12684), .CP(clk), .Q(inner_first_stage_data_reg[1669]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1668_ ( .D(N12683), .CP(clk), .Q(inner_first_stage_data_reg[1668]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1667_ ( .D(N12682), .CP(clk), .Q(inner_first_stage_data_reg[1667]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1666_ ( .D(N12681), .CP(clk), .Q(inner_first_stage_data_reg[1666]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1665_ ( .D(N12680), .CP(clk), .Q(inner_first_stage_data_reg[1665]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1664_ ( .D(N12679), .CP(clk), .Q(inner_first_stage_data_reg[1664]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_52_ ( .D(N12678), .CP(clk), 
        .Q(inner_first_stage_valid_reg[52]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1727_ ( .D(N12926), .CP(clk), .Q(inner_first_stage_data_reg[1727]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1726_ ( .D(N12925), .CP(clk), .Q(inner_first_stage_data_reg[1726]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1725_ ( .D(N12924), .CP(clk), .Q(inner_first_stage_data_reg[1725]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1724_ ( .D(N12923), .CP(clk), .Q(inner_first_stage_data_reg[1724]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1723_ ( .D(N12922), .CP(clk), .Q(inner_first_stage_data_reg[1723]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1722_ ( .D(N12921), .CP(clk), .Q(inner_first_stage_data_reg[1722]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1721_ ( .D(N12920), .CP(clk), .Q(inner_first_stage_data_reg[1721]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1720_ ( .D(N12919), .CP(clk), .Q(inner_first_stage_data_reg[1720]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1719_ ( .D(N12918), .CP(clk), .Q(inner_first_stage_data_reg[1719]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1718_ ( .D(N12917), .CP(clk), .Q(inner_first_stage_data_reg[1718]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1717_ ( .D(N12916), .CP(clk), .Q(inner_first_stage_data_reg[1717]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1716_ ( .D(N12915), .CP(clk), .Q(inner_first_stage_data_reg[1716]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1715_ ( .D(N12914), .CP(clk), .Q(inner_first_stage_data_reg[1715]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1714_ ( .D(N12913), .CP(clk), .Q(inner_first_stage_data_reg[1714]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1713_ ( .D(N12912), .CP(clk), .Q(inner_first_stage_data_reg[1713]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1712_ ( .D(N12911), .CP(clk), .Q(inner_first_stage_data_reg[1712]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1711_ ( .D(N12910), .CP(clk), .Q(inner_first_stage_data_reg[1711]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1710_ ( .D(N12909), .CP(clk), .Q(inner_first_stage_data_reg[1710]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1709_ ( .D(N12908), .CP(clk), .Q(inner_first_stage_data_reg[1709]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1708_ ( .D(N12907), .CP(clk), .Q(inner_first_stage_data_reg[1708]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1707_ ( .D(N12906), .CP(clk), .Q(inner_first_stage_data_reg[1707]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1706_ ( .D(N12905), .CP(clk), .Q(inner_first_stage_data_reg[1706]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1705_ ( .D(N12904), .CP(clk), .Q(inner_first_stage_data_reg[1705]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1704_ ( .D(N12903), .CP(clk), .Q(inner_first_stage_data_reg[1704]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1703_ ( .D(N12902), .CP(clk), .Q(inner_first_stage_data_reg[1703]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1702_ ( .D(N12901), .CP(clk), .Q(inner_first_stage_data_reg[1702]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1701_ ( .D(N12900), .CP(clk), .Q(inner_first_stage_data_reg[1701]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1700_ ( .D(N12899), .CP(clk), .Q(inner_first_stage_data_reg[1700]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1699_ ( .D(N12898), .CP(clk), .Q(inner_first_stage_data_reg[1699]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1698_ ( .D(N12897), .CP(clk), .Q(inner_first_stage_data_reg[1698]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1697_ ( .D(N12896), .CP(clk), .Q(inner_first_stage_data_reg[1697]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1696_ ( .D(N12895), .CP(clk), .Q(inner_first_stage_data_reg[1696]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_53_ ( .D(N12894), .CP(clk), 
        .Q(inner_first_stage_valid_reg[53]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1759_ ( .D(N13142), .CP(clk), .Q(inner_first_stage_data_reg[1759]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1758_ ( .D(N13141), .CP(clk), .Q(inner_first_stage_data_reg[1758]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1757_ ( .D(N13140), .CP(clk), .Q(inner_first_stage_data_reg[1757]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1756_ ( .D(N13139), .CP(clk), .Q(inner_first_stage_data_reg[1756]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1755_ ( .D(N13138), .CP(clk), .Q(inner_first_stage_data_reg[1755]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1754_ ( .D(N13137), .CP(clk), .Q(inner_first_stage_data_reg[1754]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1753_ ( .D(N13136), .CP(clk), .Q(inner_first_stage_data_reg[1753]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1752_ ( .D(N13135), .CP(clk), .Q(inner_first_stage_data_reg[1752]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1751_ ( .D(N13134), .CP(clk), .Q(inner_first_stage_data_reg[1751]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1750_ ( .D(N13133), .CP(clk), .Q(inner_first_stage_data_reg[1750]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1749_ ( .D(N13132), .CP(clk), .Q(inner_first_stage_data_reg[1749]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1748_ ( .D(N13131), .CP(clk), .Q(inner_first_stage_data_reg[1748]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1747_ ( .D(N13130), .CP(clk), .Q(inner_first_stage_data_reg[1747]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1746_ ( .D(N13129), .CP(clk), .Q(inner_first_stage_data_reg[1746]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1745_ ( .D(N13128), .CP(clk), .Q(inner_first_stage_data_reg[1745]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1744_ ( .D(N13127), .CP(clk), .Q(inner_first_stage_data_reg[1744]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1743_ ( .D(N13126), .CP(clk), .Q(inner_first_stage_data_reg[1743]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1742_ ( .D(N13125), .CP(clk), .Q(inner_first_stage_data_reg[1742]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1741_ ( .D(N13124), .CP(clk), .Q(inner_first_stage_data_reg[1741]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1740_ ( .D(N13123), .CP(clk), .Q(inner_first_stage_data_reg[1740]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1739_ ( .D(N13122), .CP(clk), .Q(inner_first_stage_data_reg[1739]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1738_ ( .D(N13121), .CP(clk), .Q(inner_first_stage_data_reg[1738]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1737_ ( .D(N13120), .CP(clk), .Q(inner_first_stage_data_reg[1737]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1736_ ( .D(N13119), .CP(clk), .Q(inner_first_stage_data_reg[1736]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1735_ ( .D(N13118), .CP(clk), .Q(inner_first_stage_data_reg[1735]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1734_ ( .D(N13117), .CP(clk), .Q(inner_first_stage_data_reg[1734]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1733_ ( .D(N13116), .CP(clk), .Q(inner_first_stage_data_reg[1733]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1732_ ( .D(N13115), .CP(clk), .Q(inner_first_stage_data_reg[1732]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1731_ ( .D(N13114), .CP(clk), .Q(inner_first_stage_data_reg[1731]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1730_ ( .D(N13113), .CP(clk), .Q(inner_first_stage_data_reg[1730]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1729_ ( .D(N13112), .CP(clk), .Q(inner_first_stage_data_reg[1729]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1728_ ( .D(N13111), .CP(clk), .Q(inner_first_stage_data_reg[1728]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_54_ ( .D(N13110), .CP(clk), 
        .Q(inner_first_stage_valid_reg[54]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1791_ ( .D(N13358), .CP(clk), .Q(inner_first_stage_data_reg[1791]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1790_ ( .D(N13357), .CP(clk), .Q(inner_first_stage_data_reg[1790]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1789_ ( .D(N13356), .CP(clk), .Q(inner_first_stage_data_reg[1789]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1788_ ( .D(N13355), .CP(clk), .Q(inner_first_stage_data_reg[1788]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1787_ ( .D(N13354), .CP(clk), .Q(inner_first_stage_data_reg[1787]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1786_ ( .D(N13353), .CP(clk), .Q(inner_first_stage_data_reg[1786]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1785_ ( .D(N13352), .CP(clk), .Q(inner_first_stage_data_reg[1785]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1784_ ( .D(N13351), .CP(clk), .Q(inner_first_stage_data_reg[1784]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1783_ ( .D(N13350), .CP(clk), .Q(inner_first_stage_data_reg[1783]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1782_ ( .D(N13349), .CP(clk), .Q(inner_first_stage_data_reg[1782]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1781_ ( .D(N13348), .CP(clk), .Q(inner_first_stage_data_reg[1781]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1780_ ( .D(N13347), .CP(clk), .Q(inner_first_stage_data_reg[1780]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1779_ ( .D(N13346), .CP(clk), .Q(inner_first_stage_data_reg[1779]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1778_ ( .D(N13345), .CP(clk), .Q(inner_first_stage_data_reg[1778]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1777_ ( .D(N13344), .CP(clk), .Q(inner_first_stage_data_reg[1777]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1776_ ( .D(N13343), .CP(clk), .Q(inner_first_stage_data_reg[1776]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1775_ ( .D(N13342), .CP(clk), .Q(inner_first_stage_data_reg[1775]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1774_ ( .D(N13341), .CP(clk), .Q(inner_first_stage_data_reg[1774]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1773_ ( .D(N13340), .CP(clk), .Q(inner_first_stage_data_reg[1773]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1772_ ( .D(N13339), .CP(clk), .Q(inner_first_stage_data_reg[1772]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1771_ ( .D(N13338), .CP(clk), .Q(inner_first_stage_data_reg[1771]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1770_ ( .D(N13337), .CP(clk), .Q(inner_first_stage_data_reg[1770]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1769_ ( .D(N13336), .CP(clk), .Q(inner_first_stage_data_reg[1769]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1768_ ( .D(N13335), .CP(clk), .Q(inner_first_stage_data_reg[1768]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1767_ ( .D(N13334), .CP(clk), .Q(inner_first_stage_data_reg[1767]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1766_ ( .D(N13333), .CP(clk), .Q(inner_first_stage_data_reg[1766]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1765_ ( .D(N13332), .CP(clk), .Q(inner_first_stage_data_reg[1765]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1764_ ( .D(N13331), .CP(clk), .Q(inner_first_stage_data_reg[1764]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1763_ ( .D(N13330), .CP(clk), .Q(inner_first_stage_data_reg[1763]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1762_ ( .D(N13329), .CP(clk), .Q(inner_first_stage_data_reg[1762]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1761_ ( .D(N13328), .CP(clk), .Q(inner_first_stage_data_reg[1761]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1760_ ( .D(N13327), .CP(clk), .Q(inner_first_stage_data_reg[1760]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_55_ ( .D(N13326), .CP(clk), 
        .Q(inner_first_stage_valid_reg[55]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1823_ ( .D(N13720), .CP(clk), .Q(inner_first_stage_data_reg[1823]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1822_ ( .D(N13719), .CP(clk), .Q(inner_first_stage_data_reg[1822]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1821_ ( .D(N13718), .CP(clk), .Q(inner_first_stage_data_reg[1821]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1820_ ( .D(N13717), .CP(clk), .Q(inner_first_stage_data_reg[1820]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1819_ ( .D(N13716), .CP(clk), .Q(inner_first_stage_data_reg[1819]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1818_ ( .D(N13715), .CP(clk), .Q(inner_first_stage_data_reg[1818]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1817_ ( .D(N13714), .CP(clk), .Q(inner_first_stage_data_reg[1817]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1816_ ( .D(N13713), .CP(clk), .Q(inner_first_stage_data_reg[1816]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1815_ ( .D(N13712), .CP(clk), .Q(inner_first_stage_data_reg[1815]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1814_ ( .D(N13711), .CP(clk), .Q(inner_first_stage_data_reg[1814]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1813_ ( .D(N13710), .CP(clk), .Q(inner_first_stage_data_reg[1813]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1812_ ( .D(N13709), .CP(clk), .Q(inner_first_stage_data_reg[1812]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1811_ ( .D(N13708), .CP(clk), .Q(inner_first_stage_data_reg[1811]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1810_ ( .D(N13707), .CP(clk), .Q(inner_first_stage_data_reg[1810]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1809_ ( .D(N13706), .CP(clk), .Q(inner_first_stage_data_reg[1809]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1808_ ( .D(N13705), .CP(clk), .Q(inner_first_stage_data_reg[1808]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1807_ ( .D(N13704), .CP(clk), .Q(inner_first_stage_data_reg[1807]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1806_ ( .D(N13703), .CP(clk), .Q(inner_first_stage_data_reg[1806]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1805_ ( .D(N13702), .CP(clk), .Q(inner_first_stage_data_reg[1805]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1804_ ( .D(N13701), .CP(clk), .Q(inner_first_stage_data_reg[1804]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1803_ ( .D(N13700), .CP(clk), .Q(inner_first_stage_data_reg[1803]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1802_ ( .D(N13699), .CP(clk), .Q(inner_first_stage_data_reg[1802]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1801_ ( .D(N13698), .CP(clk), .Q(inner_first_stage_data_reg[1801]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1800_ ( .D(N13697), .CP(clk), .Q(inner_first_stage_data_reg[1800]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1799_ ( .D(N13696), .CP(clk), .Q(inner_first_stage_data_reg[1799]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1798_ ( .D(N13695), .CP(clk), .Q(inner_first_stage_data_reg[1798]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1797_ ( .D(N13694), .CP(clk), .Q(inner_first_stage_data_reg[1797]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1796_ ( .D(N13693), .CP(clk), .Q(inner_first_stage_data_reg[1796]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1795_ ( .D(N13692), .CP(clk), .Q(inner_first_stage_data_reg[1795]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1794_ ( .D(N13691), .CP(clk), .Q(inner_first_stage_data_reg[1794]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1793_ ( .D(N13690), .CP(clk), .Q(inner_first_stage_data_reg[1793]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1792_ ( .D(N13689), .CP(clk), .Q(inner_first_stage_data_reg[1792]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_56_ ( .D(N13688), .CP(clk), 
        .Q(inner_first_stage_valid_reg[56]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1855_ ( .D(N13936), .CP(clk), .Q(inner_first_stage_data_reg[1855]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1854_ ( .D(N13935), .CP(clk), .Q(inner_first_stage_data_reg[1854]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1853_ ( .D(N13934), .CP(clk), .Q(inner_first_stage_data_reg[1853]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1852_ ( .D(N13933), .CP(clk), .Q(inner_first_stage_data_reg[1852]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1851_ ( .D(N13932), .CP(clk), .Q(inner_first_stage_data_reg[1851]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1850_ ( .D(N13931), .CP(clk), .Q(inner_first_stage_data_reg[1850]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1849_ ( .D(N13930), .CP(clk), .Q(inner_first_stage_data_reg[1849]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1848_ ( .D(N13929), .CP(clk), .Q(inner_first_stage_data_reg[1848]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1847_ ( .D(N13928), .CP(clk), .Q(inner_first_stage_data_reg[1847]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1846_ ( .D(N13927), .CP(clk), .Q(inner_first_stage_data_reg[1846]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1845_ ( .D(N13926), .CP(clk), .Q(inner_first_stage_data_reg[1845]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1844_ ( .D(N13925), .CP(clk), .Q(inner_first_stage_data_reg[1844]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1843_ ( .D(N13924), .CP(clk), .Q(inner_first_stage_data_reg[1843]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1842_ ( .D(N13923), .CP(clk), .Q(inner_first_stage_data_reg[1842]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1841_ ( .D(N13922), .CP(clk), .Q(inner_first_stage_data_reg[1841]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1840_ ( .D(N13921), .CP(clk), .Q(inner_first_stage_data_reg[1840]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1839_ ( .D(N13920), .CP(clk), .Q(inner_first_stage_data_reg[1839]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1838_ ( .D(N13919), .CP(clk), .Q(inner_first_stage_data_reg[1838]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1837_ ( .D(N13918), .CP(clk), .Q(inner_first_stage_data_reg[1837]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1836_ ( .D(N13917), .CP(clk), .Q(inner_first_stage_data_reg[1836]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1835_ ( .D(N13916), .CP(clk), .Q(inner_first_stage_data_reg[1835]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1834_ ( .D(N13915), .CP(clk), .Q(inner_first_stage_data_reg[1834]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1833_ ( .D(N13914), .CP(clk), .Q(inner_first_stage_data_reg[1833]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1832_ ( .D(N13913), .CP(clk), .Q(inner_first_stage_data_reg[1832]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1831_ ( .D(N13912), .CP(clk), .Q(inner_first_stage_data_reg[1831]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1830_ ( .D(N13911), .CP(clk), .Q(inner_first_stage_data_reg[1830]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1829_ ( .D(N13910), .CP(clk), .Q(inner_first_stage_data_reg[1829]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1828_ ( .D(N13909), .CP(clk), .Q(inner_first_stage_data_reg[1828]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1827_ ( .D(N13908), .CP(clk), .Q(inner_first_stage_data_reg[1827]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1826_ ( .D(N13907), .CP(clk), .Q(inner_first_stage_data_reg[1826]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1825_ ( .D(N13906), .CP(clk), .Q(inner_first_stage_data_reg[1825]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1824_ ( .D(N13905), .CP(clk), .Q(inner_first_stage_data_reg[1824]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_57_ ( .D(N13904), .CP(clk), 
        .Q(inner_first_stage_valid_reg[57]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1887_ ( .D(N14152), .CP(clk), .Q(inner_first_stage_data_reg[1887]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1886_ ( .D(N14151), .CP(clk), .Q(inner_first_stage_data_reg[1886]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1885_ ( .D(N14150), .CP(clk), .Q(inner_first_stage_data_reg[1885]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1884_ ( .D(N14149), .CP(clk), .Q(inner_first_stage_data_reg[1884]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1883_ ( .D(N14148), .CP(clk), .Q(inner_first_stage_data_reg[1883]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1882_ ( .D(N14147), .CP(clk), .Q(inner_first_stage_data_reg[1882]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1881_ ( .D(N14146), .CP(clk), .Q(inner_first_stage_data_reg[1881]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1880_ ( .D(N14145), .CP(clk), .Q(inner_first_stage_data_reg[1880]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1879_ ( .D(N14144), .CP(clk), .Q(inner_first_stage_data_reg[1879]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1878_ ( .D(N14143), .CP(clk), .Q(inner_first_stage_data_reg[1878]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1877_ ( .D(N14142), .CP(clk), .Q(inner_first_stage_data_reg[1877]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1876_ ( .D(N14141), .CP(clk), .Q(inner_first_stage_data_reg[1876]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1875_ ( .D(N14140), .CP(clk), .Q(inner_first_stage_data_reg[1875]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1874_ ( .D(N14139), .CP(clk), .Q(inner_first_stage_data_reg[1874]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1873_ ( .D(N14138), .CP(clk), .Q(inner_first_stage_data_reg[1873]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1872_ ( .D(N14137), .CP(clk), .Q(inner_first_stage_data_reg[1872]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1871_ ( .D(N14136), .CP(clk), .Q(inner_first_stage_data_reg[1871]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1870_ ( .D(N14135), .CP(clk), .Q(inner_first_stage_data_reg[1870]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1869_ ( .D(N14134), .CP(clk), .Q(inner_first_stage_data_reg[1869]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1868_ ( .D(N14133), .CP(clk), .Q(inner_first_stage_data_reg[1868]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1867_ ( .D(N14132), .CP(clk), .Q(inner_first_stage_data_reg[1867]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1866_ ( .D(N14131), .CP(clk), .Q(inner_first_stage_data_reg[1866]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1865_ ( .D(N14130), .CP(clk), .Q(inner_first_stage_data_reg[1865]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1864_ ( .D(N14129), .CP(clk), .Q(inner_first_stage_data_reg[1864]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1863_ ( .D(N14128), .CP(clk), .Q(inner_first_stage_data_reg[1863]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1862_ ( .D(N14127), .CP(clk), .Q(inner_first_stage_data_reg[1862]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1861_ ( .D(N14126), .CP(clk), .Q(inner_first_stage_data_reg[1861]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1860_ ( .D(N14125), .CP(clk), .Q(inner_first_stage_data_reg[1860]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1859_ ( .D(N14124), .CP(clk), .Q(inner_first_stage_data_reg[1859]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1858_ ( .D(N14123), .CP(clk), .Q(inner_first_stage_data_reg[1858]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1857_ ( .D(N14122), .CP(clk), .Q(inner_first_stage_data_reg[1857]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1856_ ( .D(N14121), .CP(clk), .Q(inner_first_stage_data_reg[1856]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_58_ ( .D(N14120), .CP(clk), 
        .Q(inner_first_stage_valid_reg[58]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1919_ ( .D(N14368), .CP(clk), .Q(inner_first_stage_data_reg[1919]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1918_ ( .D(N14367), .CP(clk), .Q(inner_first_stage_data_reg[1918]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1917_ ( .D(N14366), .CP(clk), .Q(inner_first_stage_data_reg[1917]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1916_ ( .D(N14365), .CP(clk), .Q(inner_first_stage_data_reg[1916]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1915_ ( .D(N14364), .CP(clk), .Q(inner_first_stage_data_reg[1915]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1914_ ( .D(N14363), .CP(clk), .Q(inner_first_stage_data_reg[1914]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1913_ ( .D(N14362), .CP(clk), .Q(inner_first_stage_data_reg[1913]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1912_ ( .D(N14361), .CP(clk), .Q(inner_first_stage_data_reg[1912]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1911_ ( .D(N14360), .CP(clk), .Q(inner_first_stage_data_reg[1911]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1910_ ( .D(N14359), .CP(clk), .Q(inner_first_stage_data_reg[1910]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1909_ ( .D(N14358), .CP(clk), .Q(inner_first_stage_data_reg[1909]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1908_ ( .D(N14357), .CP(clk), .Q(inner_first_stage_data_reg[1908]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1907_ ( .D(N14356), .CP(clk), .Q(inner_first_stage_data_reg[1907]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1906_ ( .D(N14355), .CP(clk), .Q(inner_first_stage_data_reg[1906]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1905_ ( .D(N14354), .CP(clk), .Q(inner_first_stage_data_reg[1905]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1904_ ( .D(N14353), .CP(clk), .Q(inner_first_stage_data_reg[1904]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1903_ ( .D(N14352), .CP(clk), .Q(inner_first_stage_data_reg[1903]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1902_ ( .D(N14351), .CP(clk), .Q(inner_first_stage_data_reg[1902]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1901_ ( .D(N14350), .CP(clk), .Q(inner_first_stage_data_reg[1901]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1900_ ( .D(N14349), .CP(clk), .Q(inner_first_stage_data_reg[1900]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1899_ ( .D(N14348), .CP(clk), .Q(inner_first_stage_data_reg[1899]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1898_ ( .D(N14347), .CP(clk), .Q(inner_first_stage_data_reg[1898]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1897_ ( .D(N14346), .CP(clk), .Q(inner_first_stage_data_reg[1897]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1896_ ( .D(N14345), .CP(clk), .Q(inner_first_stage_data_reg[1896]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1895_ ( .D(N14344), .CP(clk), .Q(inner_first_stage_data_reg[1895]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1894_ ( .D(N14343), .CP(clk), .Q(inner_first_stage_data_reg[1894]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1893_ ( .D(N14342), .CP(clk), .Q(inner_first_stage_data_reg[1893]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1892_ ( .D(N14341), .CP(clk), .Q(inner_first_stage_data_reg[1892]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1891_ ( .D(N14340), .CP(clk), .Q(inner_first_stage_data_reg[1891]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1890_ ( .D(N14339), .CP(clk), .Q(inner_first_stage_data_reg[1890]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1889_ ( .D(N14338), .CP(clk), .Q(inner_first_stage_data_reg[1889]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1888_ ( .D(N14337), .CP(clk), .Q(inner_first_stage_data_reg[1888]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_59_ ( .D(N14336), .CP(clk), 
        .Q(inner_first_stage_valid_reg[59]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1951_ ( .D(N14584), .CP(clk), .Q(inner_first_stage_data_reg[1951]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1950_ ( .D(N14583), .CP(clk), .Q(inner_first_stage_data_reg[1950]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1949_ ( .D(N14582), .CP(clk), .Q(inner_first_stage_data_reg[1949]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1948_ ( .D(N14581), .CP(clk), .Q(inner_first_stage_data_reg[1948]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1947_ ( .D(N14580), .CP(clk), .Q(inner_first_stage_data_reg[1947]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1946_ ( .D(N14579), .CP(clk), .Q(inner_first_stage_data_reg[1946]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1945_ ( .D(N14578), .CP(clk), .Q(inner_first_stage_data_reg[1945]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1944_ ( .D(N14577), .CP(clk), .Q(inner_first_stage_data_reg[1944]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1943_ ( .D(N14576), .CP(clk), .Q(inner_first_stage_data_reg[1943]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1942_ ( .D(N14575), .CP(clk), .Q(inner_first_stage_data_reg[1942]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1941_ ( .D(N14574), .CP(clk), .Q(inner_first_stage_data_reg[1941]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1940_ ( .D(N14573), .CP(clk), .Q(inner_first_stage_data_reg[1940]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1939_ ( .D(N14572), .CP(clk), .Q(inner_first_stage_data_reg[1939]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1938_ ( .D(N14571), .CP(clk), .Q(inner_first_stage_data_reg[1938]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1937_ ( .D(N14570), .CP(clk), .Q(inner_first_stage_data_reg[1937]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1936_ ( .D(N14569), .CP(clk), .Q(inner_first_stage_data_reg[1936]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1935_ ( .D(N14568), .CP(clk), .Q(inner_first_stage_data_reg[1935]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1934_ ( .D(N14567), .CP(clk), .Q(inner_first_stage_data_reg[1934]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1933_ ( .D(N14566), .CP(clk), .Q(inner_first_stage_data_reg[1933]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1932_ ( .D(N14565), .CP(clk), .Q(inner_first_stage_data_reg[1932]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1931_ ( .D(N14564), .CP(clk), .Q(inner_first_stage_data_reg[1931]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1930_ ( .D(N14563), .CP(clk), .Q(inner_first_stage_data_reg[1930]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1929_ ( .D(N14562), .CP(clk), .Q(inner_first_stage_data_reg[1929]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1928_ ( .D(N14561), .CP(clk), .Q(inner_first_stage_data_reg[1928]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1927_ ( .D(N14560), .CP(clk), .Q(inner_first_stage_data_reg[1927]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1926_ ( .D(N14559), .CP(clk), .Q(inner_first_stage_data_reg[1926]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1925_ ( .D(N14558), .CP(clk), .Q(inner_first_stage_data_reg[1925]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1924_ ( .D(N14557), .CP(clk), .Q(inner_first_stage_data_reg[1924]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1923_ ( .D(N14556), .CP(clk), .Q(inner_first_stage_data_reg[1923]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1922_ ( .D(N14555), .CP(clk), .Q(inner_first_stage_data_reg[1922]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1921_ ( .D(N14554), .CP(clk), .Q(inner_first_stage_data_reg[1921]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1920_ ( .D(N14553), .CP(clk), .Q(inner_first_stage_data_reg[1920]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_60_ ( .D(N14552), .CP(clk), 
        .Q(inner_first_stage_valid_reg[60]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1983_ ( .D(N14800), .CP(clk), .Q(inner_first_stage_data_reg[1983]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1982_ ( .D(N14799), .CP(clk), .Q(inner_first_stage_data_reg[1982]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1981_ ( .D(N14798), .CP(clk), .Q(inner_first_stage_data_reg[1981]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1980_ ( .D(N14797), .CP(clk), .Q(inner_first_stage_data_reg[1980]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1979_ ( .D(N14796), .CP(clk), .Q(inner_first_stage_data_reg[1979]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1978_ ( .D(N14795), .CP(clk), .Q(inner_first_stage_data_reg[1978]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1977_ ( .D(N14794), .CP(clk), .Q(inner_first_stage_data_reg[1977]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1976_ ( .D(N14793), .CP(clk), .Q(inner_first_stage_data_reg[1976]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1975_ ( .D(N14792), .CP(clk), .Q(inner_first_stage_data_reg[1975]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1974_ ( .D(N14791), .CP(clk), .Q(inner_first_stage_data_reg[1974]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1973_ ( .D(N14790), .CP(clk), .Q(inner_first_stage_data_reg[1973]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1972_ ( .D(N14789), .CP(clk), .Q(inner_first_stage_data_reg[1972]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1971_ ( .D(N14788), .CP(clk), .Q(inner_first_stage_data_reg[1971]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1970_ ( .D(N14787), .CP(clk), .Q(inner_first_stage_data_reg[1970]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1969_ ( .D(N14786), .CP(clk), .Q(inner_first_stage_data_reg[1969]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1968_ ( .D(N14785), .CP(clk), .Q(inner_first_stage_data_reg[1968]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1967_ ( .D(N14784), .CP(clk), .Q(inner_first_stage_data_reg[1967]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1966_ ( .D(N14783), .CP(clk), .Q(inner_first_stage_data_reg[1966]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1965_ ( .D(N14782), .CP(clk), .Q(inner_first_stage_data_reg[1965]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1964_ ( .D(N14781), .CP(clk), .Q(inner_first_stage_data_reg[1964]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1963_ ( .D(N14780), .CP(clk), .Q(inner_first_stage_data_reg[1963]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1962_ ( .D(N14779), .CP(clk), .Q(inner_first_stage_data_reg[1962]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1961_ ( .D(N14778), .CP(clk), .Q(inner_first_stage_data_reg[1961]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1960_ ( .D(N14777), .CP(clk), .Q(inner_first_stage_data_reg[1960]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1959_ ( .D(N14776), .CP(clk), .Q(inner_first_stage_data_reg[1959]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1958_ ( .D(N14775), .CP(clk), .Q(inner_first_stage_data_reg[1958]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1957_ ( .D(N14774), .CP(clk), .Q(inner_first_stage_data_reg[1957]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1956_ ( .D(N14773), .CP(clk), .Q(inner_first_stage_data_reg[1956]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1955_ ( .D(N14772), .CP(clk), .Q(inner_first_stage_data_reg[1955]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1954_ ( .D(N14771), .CP(clk), .Q(inner_first_stage_data_reg[1954]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1953_ ( .D(N14770), .CP(clk), .Q(inner_first_stage_data_reg[1953]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1952_ ( .D(N14769), .CP(clk), .Q(inner_first_stage_data_reg[1952]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_61_ ( .D(N14768), .CP(clk), 
        .Q(inner_first_stage_valid_reg[61]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2015_ ( .D(N15016), .CP(clk), .Q(inner_first_stage_data_reg[2015]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2014_ ( .D(N15015), .CP(clk), .Q(inner_first_stage_data_reg[2014]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2013_ ( .D(N15014), .CP(clk), .Q(inner_first_stage_data_reg[2013]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2012_ ( .D(N15013), .CP(clk), .Q(inner_first_stage_data_reg[2012]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2011_ ( .D(N15012), .CP(clk), .Q(inner_first_stage_data_reg[2011]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2010_ ( .D(N15011), .CP(clk), .Q(inner_first_stage_data_reg[2010]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2009_ ( .D(N15010), .CP(clk), .Q(inner_first_stage_data_reg[2009]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2008_ ( .D(N15009), .CP(clk), .Q(inner_first_stage_data_reg[2008]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2007_ ( .D(N15008), .CP(clk), .Q(inner_first_stage_data_reg[2007]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2006_ ( .D(N15007), .CP(clk), .Q(inner_first_stage_data_reg[2006]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2005_ ( .D(N15006), .CP(clk), .Q(inner_first_stage_data_reg[2005]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2004_ ( .D(N15005), .CP(clk), .Q(inner_first_stage_data_reg[2004]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2003_ ( .D(N15004), .CP(clk), .Q(inner_first_stage_data_reg[2003]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2002_ ( .D(N15003), .CP(clk), .Q(inner_first_stage_data_reg[2002]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2001_ ( .D(N15002), .CP(clk), .Q(inner_first_stage_data_reg[2001]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2000_ ( .D(N15001), .CP(clk), .Q(inner_first_stage_data_reg[2000]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1999_ ( .D(N15000), .CP(clk), .Q(inner_first_stage_data_reg[1999]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1998_ ( .D(N14999), .CP(clk), .Q(inner_first_stage_data_reg[1998]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1997_ ( .D(N14998), .CP(clk), .Q(inner_first_stage_data_reg[1997]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1996_ ( .D(N14997), .CP(clk), .Q(inner_first_stage_data_reg[1996]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1995_ ( .D(N14996), .CP(clk), .Q(inner_first_stage_data_reg[1995]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1994_ ( .D(N14995), .CP(clk), .Q(inner_first_stage_data_reg[1994]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1993_ ( .D(N14994), .CP(clk), .Q(inner_first_stage_data_reg[1993]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1992_ ( .D(N14993), .CP(clk), .Q(inner_first_stage_data_reg[1992]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1991_ ( .D(N14992), .CP(clk), .Q(inner_first_stage_data_reg[1991]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1990_ ( .D(N14991), .CP(clk), .Q(inner_first_stage_data_reg[1990]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1989_ ( .D(N14990), .CP(clk), .Q(inner_first_stage_data_reg[1989]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1988_ ( .D(N14989), .CP(clk), .Q(inner_first_stage_data_reg[1988]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1987_ ( .D(N14988), .CP(clk), .Q(inner_first_stage_data_reg[1987]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1986_ ( .D(N14987), .CP(clk), .Q(inner_first_stage_data_reg[1986]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1985_ ( .D(N14986), .CP(clk), .Q(inner_first_stage_data_reg[1985]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1984_ ( .D(N14985), .CP(clk), .Q(inner_first_stage_data_reg[1984]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_62_ ( .D(N14984), .CP(clk), 
        .Q(inner_first_stage_valid_reg[62]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2047_ ( .D(N15232), .CP(clk), .Q(inner_first_stage_data_reg[2047]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2046_ ( .D(N15231), .CP(clk), .Q(inner_first_stage_data_reg[2046]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2045_ ( .D(N15230), .CP(clk), .Q(inner_first_stage_data_reg[2045]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2044_ ( .D(N15229), .CP(clk), .Q(inner_first_stage_data_reg[2044]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2043_ ( .D(N15228), .CP(clk), .Q(inner_first_stage_data_reg[2043]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2042_ ( .D(N15227), .CP(clk), .Q(inner_first_stage_data_reg[2042]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2041_ ( .D(N15226), .CP(clk), .Q(inner_first_stage_data_reg[2041]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2040_ ( .D(N15225), .CP(clk), .Q(inner_first_stage_data_reg[2040]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2039_ ( .D(N15224), .CP(clk), .Q(inner_first_stage_data_reg[2039]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2038_ ( .D(N15223), .CP(clk), .Q(inner_first_stage_data_reg[2038]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2037_ ( .D(N15222), .CP(clk), .Q(inner_first_stage_data_reg[2037]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2036_ ( .D(N15221), .CP(clk), .Q(inner_first_stage_data_reg[2036]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2035_ ( .D(N15220), .CP(clk), .Q(inner_first_stage_data_reg[2035]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2034_ ( .D(N15219), .CP(clk), .Q(inner_first_stage_data_reg[2034]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2033_ ( .D(N15218), .CP(clk), .Q(inner_first_stage_data_reg[2033]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2032_ ( .D(N15217), .CP(clk), .Q(inner_first_stage_data_reg[2032]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2031_ ( .D(N15216), .CP(clk), .Q(inner_first_stage_data_reg[2031]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2030_ ( .D(N15215), .CP(clk), .Q(inner_first_stage_data_reg[2030]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2029_ ( .D(N15214), .CP(clk), .Q(inner_first_stage_data_reg[2029]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2028_ ( .D(N15213), .CP(clk), .Q(inner_first_stage_data_reg[2028]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2027_ ( .D(N15212), .CP(clk), .Q(inner_first_stage_data_reg[2027]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2026_ ( .D(N15211), .CP(clk), .Q(inner_first_stage_data_reg[2026]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2025_ ( .D(N15210), .CP(clk), .Q(inner_first_stage_data_reg[2025]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2024_ ( .D(N15209), .CP(clk), .Q(inner_first_stage_data_reg[2024]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2023_ ( .D(N15208), .CP(clk), .Q(inner_first_stage_data_reg[2023]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2022_ ( .D(N15207), .CP(clk), .Q(inner_first_stage_data_reg[2022]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2021_ ( .D(N15206), .CP(clk), .Q(inner_first_stage_data_reg[2021]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2020_ ( .D(N15205), .CP(clk), .Q(inner_first_stage_data_reg[2020]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2019_ ( .D(N15204), .CP(clk), .Q(inner_first_stage_data_reg[2019]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2018_ ( .D(N15203), .CP(clk), .Q(inner_first_stage_data_reg[2018]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2017_ ( .D(N15202), .CP(clk), .Q(inner_first_stage_data_reg[2017]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2016_ ( .D(N15201), .CP(clk), .Q(inner_first_stage_data_reg[2016]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_63_ ( .D(N15200), .CP(clk), 
        .Q(inner_first_stage_valid_reg[63]) );
  DFQD2BWP30P140LVT o_valid_reg_reg_7_ ( .D(N15346), .CP(clk), .Q(o_valid[7])
         );
  DFQD2BWP30P140LVT o_valid_reg_reg_6_ ( .D(N13472), .CP(clk), .Q(o_valid[6])
         );
  DFQD2BWP30P140LVT o_valid_reg_reg_5_ ( .D(N11598), .CP(clk), .Q(o_valid[5])
         );
  DFQD2BWP30P140LVT o_valid_reg_reg_4_ ( .D(N9724), .CP(clk), .Q(o_valid[4])
         );
  DFQD2BWP30P140LVT o_valid_reg_reg_3_ ( .D(N7850), .CP(clk), .Q(o_valid[3])
         );
  DFQD2BWP30P140LVT o_valid_reg_reg_2_ ( .D(N5976), .CP(clk), .Q(o_valid[2])
         );
  DFQD2BWP30P140LVT o_valid_reg_reg_1_ ( .D(N4102), .CP(clk), .Q(o_valid[1])
         );
  DFQD2BWP30P140LVT o_valid_reg_reg_0_ ( .D(N2228), .CP(clk), .Q(o_valid[0])
         );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N15378), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N15377), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N15376), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N15375), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N15374), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N15373), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N15372), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N15371), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N15370), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N15369), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N15368), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N15367), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N15366), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N15365), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N15364), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N15363), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N15362), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N15361), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N15360), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N15359), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N15358), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N15357), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N15356), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N15355), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N15354), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N15353), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N15352), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N15351), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N15350), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N15349), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N15348), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N15347), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N13504), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N13503), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N13502), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N13501), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N13500), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N13499), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N13498), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N13497), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N13496), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N13495), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N13494), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N13493), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N13492), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N13491), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N13490), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N13489), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N13488), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N13487), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N13486), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N13485), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N13484), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N13483), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N13482), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N13481), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N13480), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N13479), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N13478), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N13477), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N13476), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N13475), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N13474), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N13473), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N11630), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N11629), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N11628), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N11627), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N11626), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N11625), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N11624), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N11623), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N11622), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N11621), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N11620), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N11619), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N11618), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N11617), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N11616), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N11615), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N11614), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N11613), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N11612), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N11611), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N11610), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N11609), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N11608), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N11607), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N11606), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N11605), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N11604), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N11603), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N11602), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N11601), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N11600), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N11599), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N9756), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N9755), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N9754), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N9753), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N9752), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N9751), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N9750), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N9749), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N9748), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N9747), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N9746), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N9745), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N9744), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N9743), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N9742), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N9741), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N9740), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N9739), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N9738), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N9737), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N9736), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N9735), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N9734), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N9733), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N9732), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N9731), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N9730), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N9729), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N9728), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N9727), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N9726), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N9725), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N7882), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N7881), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N7880), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N7879), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N7878), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N7877), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N7876), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N7875), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N7874), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N7873), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N7872), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N7871), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N7870), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N7869), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N7868), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N7867), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N7866), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N7865), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N7864), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N7863), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N7862), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N7861), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N7860), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N7859), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N7858), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N7857), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N7856), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N7855), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N7854), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N7853), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N7852), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N7851), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N6008), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N6007), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N6006), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N6005), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N6004), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N6003), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N6002), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N6001), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N6000), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N5999), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N5998), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N5997), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N5996), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N5995), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N5994), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N5993), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N5992), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N5991), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N5990), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N5989), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N5988), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N5987), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N5986), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N5985), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N5984), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N5983), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N5982), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N5981), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N5980), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N5979), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N5978), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N5977), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N4134), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N4133), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N4132), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N4131), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N4130), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N4129), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N4128), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N4127), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N4126), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N4125), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N4124), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N4123), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N4122), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N4121), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N4120), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N4119), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N4118), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N4117), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N4116), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N4115), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N4114), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N4113), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N4112), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N4111), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N4110), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N4109), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N4108), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N4107), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N4106), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N4105), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N4104), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N4103), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N2260), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N2259), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N2258), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N2257), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N2256), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N2255), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N2254), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N2253), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N2252), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N2251), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N2250), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N2249), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N2248), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N2247), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N2246), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N2245), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N2244), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N2243), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N2242), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N2241), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N2240), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N2239), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N2238), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N2237), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N2236), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N2235), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N2234), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N2233), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N2232), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N2231), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N2230), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N2229), .CP(clk), .Q(
        o_data_bus[0]) );
  DFD1BWP30P140LVT inner_first_stage_valid_reg_reg_18_ ( .D(N4750), .CP(clk), 
        .Q(inner_first_stage_valid_reg[18]), .QN(n11767) );
  NR3D1P5BWP30P140LVT U8269 ( .A1(inner_first_stage_valid_reg[20]), .A2(n10373), .A3(n10371), .ZN(n11076) );
  INVD1BWP30P140LVT U8270 ( .I(n5891), .ZN(n11075) );
  IND2D6BWP30P140LVT U8271 ( .A1(rst), .B1(i_en), .ZN(n10380) );
  NR2D1BWP30P140LVT U8272 ( .A1(n10380), .A2(inner_first_stage_valid_reg[60]), 
        .ZN(n10295) );
  NR3D1P5BWP30P140LVT U8273 ( .A1(inner_first_stage_valid_reg[41]), .A2(n10355), .A3(n10354), .ZN(n11486) );
  OR3D1BWP30P140LVT U8274 ( .A1(inner_first_stage_valid_reg[17]), .A2(n10372), 
        .A3(n10371), .Z(n5891) );
  INR3D1BWP30P140LVT U8275 ( .A1(inner_first_stage_valid_reg[43]), .B1(
        inner_first_stage_valid_reg[42]), .B2(n10353), .ZN(n11490) );
  ND2D1BWP30P140LVT U8276 ( .A1(n6124), .A2(n6121), .ZN(n6122) );
  ND2D1BWP30P140LVT U8277 ( .A1(n5913), .A2(n5912), .ZN(n5917) );
  NR3D1P5BWP30P140LVT U8278 ( .A1(inner_first_stage_valid_reg[18]), .A2(n10368), .A3(n10367), .ZN(n11081) );
  NR3D1P5BWP30P140LVT U8279 ( .A1(inner_first_stage_valid_reg[19]), .A2(n11767), .A3(n10367), .ZN(n11082) );
  ND2D1BWP30P140LVT U8280 ( .A1(n6120), .A2(n6129), .ZN(n6127) );
  ND2D1BWP30P140LVT U8281 ( .A1(n5907), .A2(n5911), .ZN(n5915) );
  ND2D1BWP30P140LVT U8282 ( .A1(n5940), .A2(n5938), .ZN(n5941) );
  ND2D1BWP30P140LVT U8283 ( .A1(n9855), .A2(n9856), .ZN(n9859) );
  ND2D1BWP30P140LVT U8284 ( .A1(n5980), .A2(n5982), .ZN(n5983) );
  ND2D1BWP30P140LVT U8285 ( .A1(n9835), .A2(n9840), .ZN(n9836) );
  ND2D1BWP30P140LVT U8286 ( .A1(n5990), .A2(n5988), .ZN(n5991) );
  ND2D1BWP30P140LVT U8287 ( .A1(n5928), .A2(n5930), .ZN(n5931) );
  ND2D1BWP30P140LVT U8288 ( .A1(n9846), .A2(n9845), .ZN(n9849) );
  ND2D1BWP30P140LVT U8289 ( .A1(n10025), .A2(n10027), .ZN(n10029) );
  ND2D1BWP30P140LVT U8290 ( .A1(n10017), .A2(n10016), .ZN(n10020) );
  ND2D1BWP30P140LVT U8291 ( .A1(n5946), .A2(n5948), .ZN(n5949) );
  ND2D1BWP30P140LVT U8292 ( .A1(n5920), .A2(n5922), .ZN(n5923) );
  ND2D1BWP30P140LVT U8293 ( .A1(n6010), .A2(n6012), .ZN(n6013) );
  ND2D1BWP30P140LVT U8294 ( .A1(n5960), .A2(n5958), .ZN(n5961) );
  ND2D1BWP30P140LVT U8295 ( .A1(n5998), .A2(n5996), .ZN(n5999) );
  ND2D1BWP30P140LVT U8296 ( .A1(n5954), .A2(n5952), .ZN(n5955) );
  ND2D1BWP30P140LVT U8297 ( .A1(n9811), .A2(n9810), .ZN(n9814) );
  INR3D1BWP30P140LVT U8298 ( .A1(n10355), .B1(n10349), .B2(n10354), .ZN(n11487) );
  NR3D0P7BWP30P140LVT U8299 ( .A1(n10360), .A2(n10359), .A3(n10358), .ZN(n5892) );
  NR3D0P7BWP30P140LVT U8300 ( .A1(n10360), .A2(n10359), .A3(n10358), .ZN(n5893) );
  ND2OPTIBD1BWP30P140LVT U8301 ( .A1(n5900), .A2(n10347), .ZN(n10359) );
  NR2D1BWP30P140LVT U8302 ( .A1(inner_first_stage_valid_reg[12]), .A2(n10380), 
        .ZN(n10335) );
  NR2D1BWP30P140LVT U8303 ( .A1(inner_first_stage_valid_reg[36]), .A2(n10380), 
        .ZN(n6120) );
  NR2D1BWP30P140LVT U8304 ( .A1(inner_first_stage_valid_reg[42]), .A2(
        inner_first_stage_valid_reg[43]), .ZN(n10347) );
  NR2D1BWP30P140LVT U8305 ( .A1(inner_first_stage_valid_reg[0]), .A2(n5915), 
        .ZN(n5912) );
  ND2D1BWP30P140LVT U8306 ( .A1(n10338), .A2(n10335), .ZN(n10343) );
  NR2D1BWP30P140LVT U8307 ( .A1(inner_first_stage_valid_reg[32]), .A2(n6127), 
        .ZN(n6124) );
  NR2D1BWP30P140LVT U8308 ( .A1(inner_first_stage_valid_reg[2]), .A2(
        inner_first_stage_valid_reg[3]), .ZN(n5914) );
  NR2D1BWP30P140LVT U8309 ( .A1(inner_first_stage_valid_reg[4]), .A2(n10380), 
        .ZN(n5907) );
  ND2D1BWP30P140LVT U8310 ( .A1(n10390), .A2(n10379), .ZN(n10382) );
  NR2D1BWP30P140LVT U8311 ( .A1(inner_first_stage_valid_reg[28]), .A2(n10380), 
        .ZN(n10383) );
  NR2D1BWP30P140LVT U8312 ( .A1(n10380), .A2(inner_first_stage_valid_reg[40]), 
        .ZN(n10352) );
  IND2D1BWP30P140LVT U8313 ( .A1(n5915), .B1(n5914), .ZN(n5916) );
  NR2D1BWP30P140LVT U8314 ( .A1(inner_first_stage_valid_reg[6]), .A2(
        inner_first_stage_valid_reg[7]), .ZN(n5911) );
  ND2D1BWP30P140LVT U8315 ( .A1(n5907), .A2(n5910), .ZN(n5909) );
  IND2D1BWP30P140LVT U8316 ( .A1(n10343), .B1(n10333), .ZN(n10337) );
  ND2D1BWP30P140LVT U8317 ( .A1(n10370), .A2(n10374), .ZN(n10371) );
  IND2D1BWP30P140LVT U8318 ( .A1(n10369), .B1(n10365), .ZN(n10363) );
  INVD1BWP30P140LVT U8319 ( .I(inner_first_stage_valid_reg[19]), .ZN(n10368)
         );
  ND2D1BWP30P140LVT U8320 ( .A1(n10383), .A2(n10387), .ZN(n10384) );
  IND2D1BWP30P140LVT U8321 ( .A1(n6127), .B1(n6126), .ZN(n6130) );
  NR2D1BWP30P140LVT U8322 ( .A1(inner_first_stage_valid_reg[39]), .A2(
        inner_first_stage_valid_reg[38]), .ZN(n6129) );
  ND2D1BWP30P140LVT U8323 ( .A1(n6120), .A2(n6128), .ZN(n6123) );
  IND2D1BWP30P140LVT U8324 ( .A1(n10358), .B1(n10352), .ZN(n10353) );
  ND2OPTIBD1BWP30P140LVT U8325 ( .A1(n10348), .A2(n10360), .ZN(n10354) );
  INVD1BWP30P140LVT U8326 ( .I(inner_first_stage_valid_reg[40]), .ZN(n10360)
         );
  OR2D1BWP30P140LVT U8327 ( .A1(n10357), .A2(inner_first_stage_valid_reg[44]), 
        .Z(n10356) );
  INVD1BWP30P140LVT U8328 ( .I(n10380), .ZN(n5900) );
  ND2D1BWP30P140LVT U8329 ( .A1(n5898), .A2(n5901), .ZN(n5899) );
  NR2D1BWP30P140LVT U8330 ( .A1(inner_first_stage_valid_reg[52]), .A2(n10380), 
        .ZN(n5898) );
  ND2D1BWP30P140LVT U8331 ( .A1(n5896), .A2(n5895), .ZN(n5897) );
  ND2D1BWP30P140LVT U8332 ( .A1(n5894), .A2(n5895), .ZN(n5903) );
  OR2D1BWP30P140LVT U8333 ( .A1(n5899), .A2(inner_first_stage_valid_reg[51]), 
        .Z(n5904) );
  ND2D1BWP30P140LVT U8334 ( .A1(n10296), .A2(n10298), .ZN(n10293) );
  ND2D1BWP30P140LVT U8335 ( .A1(n10304), .A2(n10303), .ZN(n10299) );
  ND2D1BWP30P140LVT U8336 ( .A1(n10295), .A2(n10301), .ZN(n10297) );
  INVD1BWP30P140LVT U8337 ( .I(i_cmd[247]), .ZN(n6654) );
  ND2D1BWP30P140LVT U8338 ( .A1(n6654), .A2(n6656), .ZN(n6653) );
  INVD1BWP30P140LVT U8339 ( .I(i_cmd[231]), .ZN(n6656) );
  OR2D1BWP30P140LVT U8340 ( .A1(i_cmd[255]), .A2(i_cmd[239]), .Z(n6655) );
  INVD1BWP30P140LVT U8341 ( .I(i_cmd[215]), .ZN(n6237) );
  ND2D1BWP30P140LVT U8342 ( .A1(n6237), .A2(n6236), .ZN(n6238) );
  INVD1BWP30P140LVT U8343 ( .I(i_cmd[199]), .ZN(n6236) );
  OR2D1BWP30P140LVT U8344 ( .A1(i_cmd[223]), .A2(i_cmd[207]), .Z(n6235) );
  INVD1BWP30P140LVT U8345 ( .I(i_cmd[183]), .ZN(n5998) );
  INVD1BWP30P140LVT U8346 ( .I(i_cmd[167]), .ZN(n5996) );
  OR2D1BWP30P140LVT U8347 ( .A1(i_cmd[191]), .A2(i_cmd[175]), .Z(n5997) );
  INVD1BWP30P140LVT U8348 ( .I(i_cmd[159]), .ZN(n5946) );
  INVD1BWP30P140LVT U8349 ( .I(i_cmd[143]), .ZN(n5948) );
  OR2D1BWP30P140LVT U8350 ( .A1(i_cmd[135]), .A2(i_cmd[151]), .Z(n5947) );
  INVD1BWP30P140LVT U8351 ( .I(i_cmd[119]), .ZN(n6294) );
  ND2D1BWP30P140LVT U8352 ( .A1(n6294), .A2(n6296), .ZN(n6293) );
  INVD1BWP30P140LVT U8353 ( .I(i_cmd[103]), .ZN(n6296) );
  OR2D1BWP30P140LVT U8354 ( .A1(i_cmd[127]), .A2(i_cmd[111]), .Z(n6295) );
  INVD1BWP30P140LVT U8355 ( .I(i_cmd[95]), .ZN(n6276) );
  ND2D1BWP30P140LVT U8356 ( .A1(n6276), .A2(n6278), .ZN(n6275) );
  INVD1BWP30P140LVT U8357 ( .I(i_cmd[79]), .ZN(n6278) );
  OR2D1BWP30P140LVT U8358 ( .A1(i_cmd[71]), .A2(i_cmd[87]), .Z(n6277) );
  INVD1BWP30P140LVT U8359 ( .I(i_cmd[39]), .ZN(n6367) );
  ND2D1BWP30P140LVT U8360 ( .A1(n6367), .A2(n6370), .ZN(n6368) );
  INVD1BWP30P140LVT U8361 ( .I(i_cmd[55]), .ZN(n6370) );
  OR2D1BWP30P140LVT U8362 ( .A1(i_cmd[63]), .A2(i_cmd[47]), .Z(n6369) );
  INVD1BWP30P140LVT U8363 ( .I(i_cmd[23]), .ZN(n7831) );
  ND2D1BWP30P140LVT U8364 ( .A1(n7831), .A2(n7833), .ZN(n7834) );
  INVD1BWP30P140LVT U8365 ( .I(i_cmd[7]), .ZN(n7833) );
  OR2D1BWP30P140LVT U8366 ( .A1(i_cmd[31]), .A2(i_cmd[15]), .Z(n7832) );
  INVD1BWP30P140LVT U8367 ( .I(i_cmd[246]), .ZN(n5928) );
  INVD1BWP30P140LVT U8368 ( .I(i_cmd[230]), .ZN(n5930) );
  OR2D1BWP30P140LVT U8369 ( .A1(i_cmd[254]), .A2(i_cmd[238]), .Z(n5929) );
  INVD1BWP30P140LVT U8370 ( .I(i_cmd[214]), .ZN(n6227) );
  ND2D1BWP30P140LVT U8371 ( .A1(n6227), .A2(n6225), .ZN(n6228) );
  INVD1BWP30P140LVT U8372 ( .I(i_cmd[198]), .ZN(n6225) );
  OR2D1BWP30P140LVT U8373 ( .A1(i_cmd[222]), .A2(i_cmd[206]), .Z(n6226) );
  INVD1BWP30P140LVT U8374 ( .I(i_cmd[166]), .ZN(n6496) );
  ND2D1BWP30P140LVT U8375 ( .A1(n6496), .A2(n6498), .ZN(n6495) );
  INVD1BWP30P140LVT U8376 ( .I(i_cmd[182]), .ZN(n6498) );
  OR2D1BWP30P140LVT U8377 ( .A1(i_cmd[190]), .A2(i_cmd[174]), .Z(n6497) );
  INVD1BWP30P140LVT U8378 ( .I(i_cmd[158]), .ZN(n7037) );
  INVD1BWP30P140LVT U8379 ( .I(i_cmd[142]), .ZN(n7038) );
  OR2D1BWP30P140LVT U8380 ( .A1(i_cmd[134]), .A2(i_cmd[150]), .Z(n7039) );
  ND2D1BWP30P140LVT U8381 ( .A1(n7037), .A2(n7038), .ZN(n7040) );
  INVD1BWP30P140LVT U8382 ( .I(i_cmd[102]), .ZN(n6249) );
  ND2D1BWP30P140LVT U8383 ( .A1(n6249), .A2(n6248), .ZN(n6250) );
  INVD1BWP30P140LVT U8384 ( .I(i_cmd[118]), .ZN(n6248) );
  OR2D1BWP30P140LVT U8385 ( .A1(i_cmd[126]), .A2(i_cmd[110]), .Z(n6247) );
  INVD1BWP30P140LVT U8386 ( .I(i_cmd[94]), .ZN(n6382) );
  ND2D1BWP30P140LVT U8387 ( .A1(n6382), .A2(n6384), .ZN(n6381) );
  INVD1BWP30P140LVT U8388 ( .I(i_cmd[78]), .ZN(n6384) );
  OR2D1BWP30P140LVT U8389 ( .A1(i_cmd[70]), .A2(i_cmd[86]), .Z(n6383) );
  INVD1BWP30P140LVT U8390 ( .I(i_cmd[46]), .ZN(n6878) );
  ND2D1BWP30P140LVT U8391 ( .A1(n6878), .A2(n6880), .ZN(n6877) );
  INVD1BWP30P140LVT U8392 ( .I(i_cmd[62]), .ZN(n6880) );
  OR2D1BWP30P140LVT U8393 ( .A1(i_cmd[54]), .A2(i_cmd[38]), .Z(n6879) );
  ND2D1BWP30P140LVT U8394 ( .A1(n6647), .A2(n6650), .ZN(n6648) );
  INVD1BWP30P140LVT U8395 ( .I(i_cmd[14]), .ZN(n6647) );
  INVD1BWP30P140LVT U8396 ( .I(i_cmd[30]), .ZN(n6650) );
  OR2D1BWP30P140LVT U8397 ( .A1(i_cmd[22]), .A2(i_cmd[6]), .Z(n6649) );
  INVD1BWP30P140LVT U8398 ( .I(i_cmd[245]), .ZN(n5920) );
  INVD1BWP30P140LVT U8399 ( .I(i_cmd[229]), .ZN(n5922) );
  OR2D1BWP30P140LVT U8400 ( .A1(i_cmd[253]), .A2(i_cmd[237]), .Z(n5921) );
  INVD1BWP30P140LVT U8401 ( .I(i_cmd[221]), .ZN(n6328) );
  ND2D1BWP30P140LVT U8402 ( .A1(n6328), .A2(n6325), .ZN(n6326) );
  INVD1BWP30P140LVT U8403 ( .I(i_cmd[205]), .ZN(n6325) );
  OR2D1BWP30P140LVT U8404 ( .A1(i_cmd[213]), .A2(i_cmd[197]), .Z(n6327) );
  INVD1BWP30P140LVT U8405 ( .I(i_cmd[181]), .ZN(n6010) );
  INVD1BWP30P140LVT U8406 ( .I(i_cmd[165]), .ZN(n6012) );
  OR2D1BWP30P140LVT U8407 ( .A1(i_cmd[189]), .A2(i_cmd[173]), .Z(n6011) );
  INVD1BWP30P140LVT U8408 ( .I(i_cmd[157]), .ZN(n7163) );
  INVD1BWP30P140LVT U8409 ( .I(i_cmd[141]), .ZN(n7162) );
  OR2D1BWP30P140LVT U8410 ( .A1(i_cmd[133]), .A2(i_cmd[149]), .Z(n7161) );
  ND2D1BWP30P140LVT U8411 ( .A1(n7163), .A2(n7162), .ZN(n7164) );
  INVD1BWP30P140LVT U8412 ( .I(i_cmd[109]), .ZN(n6283) );
  ND2D1BWP30P140LVT U8413 ( .A1(n6283), .A2(n6286), .ZN(n6284) );
  INVD1BWP30P140LVT U8414 ( .I(i_cmd[125]), .ZN(n6286) );
  OR2D1BWP30P140LVT U8415 ( .A1(i_cmd[101]), .A2(i_cmd[117]), .Z(n6285) );
  INVD1BWP30P140LVT U8416 ( .I(i_cmd[93]), .ZN(n6409) );
  ND2D1BWP30P140LVT U8417 ( .A1(n6409), .A2(n6412), .ZN(n6410) );
  INVD1BWP30P140LVT U8418 ( .I(i_cmd[77]), .ZN(n6412) );
  OR2D1BWP30P140LVT U8419 ( .A1(i_cmd[85]), .A2(i_cmd[69]), .Z(n6411) );
  INVD1BWP30P140LVT U8420 ( .I(i_cmd[61]), .ZN(n6318) );
  ND2D1BWP30P140LVT U8421 ( .A1(n6318), .A2(n6320), .ZN(n6317) );
  INVD1BWP30P140LVT U8422 ( .I(i_cmd[45]), .ZN(n6320) );
  OR2D1BWP30P140LVT U8423 ( .A1(i_cmd[37]), .A2(i_cmd[53]), .Z(n6319) );
  INVD1BWP30P140LVT U8424 ( .I(i_cmd[21]), .ZN(n7270) );
  ND2D1BWP30P140LVT U8425 ( .A1(n7270), .A2(n7272), .ZN(n7269) );
  INVD1BWP30P140LVT U8426 ( .I(i_cmd[5]), .ZN(n7272) );
  OR2D1BWP30P140LVT U8427 ( .A1(i_cmd[29]), .A2(i_cmd[13]), .Z(n7271) );
  ND2D1BWP30P140LVT U8428 ( .A1(n6537), .A2(n6540), .ZN(n6538) );
  INVD1BWP30P140LVT U8429 ( .I(i_cmd[252]), .ZN(n6537) );
  INVD1BWP30P140LVT U8430 ( .I(i_cmd[236]), .ZN(n6540) );
  OR2D1BWP30P140LVT U8431 ( .A1(i_cmd[244]), .A2(i_cmd[228]), .Z(n6539) );
  INVD1BWP30P140LVT U8432 ( .I(i_cmd[196]), .ZN(n6219) );
  ND2D1BWP30P140LVT U8433 ( .A1(n6219), .A2(n6218), .ZN(n6220) );
  INVD1BWP30P140LVT U8434 ( .I(i_cmd[212]), .ZN(n6218) );
  OR2D1BWP30P140LVT U8435 ( .A1(i_cmd[220]), .A2(i_cmd[204]), .Z(n6217) );
  INVD1BWP30P140LVT U8436 ( .I(i_cmd[188]), .ZN(n7289) );
  INVD1BWP30P140LVT U8437 ( .I(i_cmd[172]), .ZN(n7290) );
  OR2D1BWP30P140LVT U8438 ( .A1(i_cmd[180]), .A2(i_cmd[164]), .Z(n7291) );
  ND2D1BWP30P140LVT U8439 ( .A1(n7290), .A2(n7289), .ZN(n7292) );
  INVD1BWP30P140LVT U8440 ( .I(i_cmd[156]), .ZN(n7253) );
  INVD1BWP30P140LVT U8441 ( .I(i_cmd[140]), .ZN(n7254) );
  OR2D1BWP30P140LVT U8442 ( .A1(i_cmd[148]), .A2(i_cmd[132]), .Z(n7255) );
  ND2D1BWP30P140LVT U8443 ( .A1(n7253), .A2(n7254), .ZN(n7256) );
  INVD1BWP30P140LVT U8444 ( .I(i_cmd[124]), .ZN(n6244) );
  ND2D1BWP30P140LVT U8445 ( .A1(n6244), .A2(n6241), .ZN(n6242) );
  INVD1BWP30P140LVT U8446 ( .I(i_cmd[108]), .ZN(n6241) );
  OR2D1BWP30P140LVT U8447 ( .A1(i_cmd[116]), .A2(i_cmd[100]), .Z(n6243) );
  INVD1BWP30P140LVT U8448 ( .I(i_cmd[92]), .ZN(n6466) );
  ND2D1BWP30P140LVT U8449 ( .A1(n6466), .A2(n6468), .ZN(n6465) );
  INVD1BWP30P140LVT U8450 ( .I(i_cmd[76]), .ZN(n6468) );
  OR2D1BWP30P140LVT U8451 ( .A1(i_cmd[84]), .A2(i_cmd[68]), .Z(n6467) );
  INVD1BWP30P140LVT U8452 ( .I(i_cmd[36]), .ZN(n6376) );
  ND2D1BWP30P140LVT U8453 ( .A1(n6376), .A2(n6378), .ZN(n6375) );
  INVD1BWP30P140LVT U8454 ( .I(i_cmd[52]), .ZN(n6378) );
  OR2D1BWP30P140LVT U8455 ( .A1(i_cmd[60]), .A2(i_cmd[44]), .Z(n6377) );
  INVD1BWP30P140LVT U8456 ( .I(i_cmd[28]), .ZN(n6431) );
  ND2D1BWP30P140LVT U8457 ( .A1(n6431), .A2(n6434), .ZN(n6432) );
  INVD1BWP30P140LVT U8458 ( .I(i_cmd[12]), .ZN(n6434) );
  OR2D1BWP30P140LVT U8459 ( .A1(i_cmd[20]), .A2(i_cmd[4]), .Z(n6433) );
  INVD1BWP30P140LVT U8460 ( .I(i_cmd[243]), .ZN(n6701) );
  INVD1BWP30P140LVT U8461 ( .I(i_cmd[227]), .ZN(n6702) );
  OR2D1BWP30P140LVT U8462 ( .A1(i_cmd[251]), .A2(i_cmd[235]), .Z(n6703) );
  ND2D1BWP30P140LVT U8463 ( .A1(n6701), .A2(n6702), .ZN(n6704) );
  INVD1BWP30P140LVT U8464 ( .I(i_cmd[203]), .ZN(n7191) );
  ND2D1BWP30P140LVT U8465 ( .A1(n7191), .A2(n7194), .ZN(n7192) );
  INVD1BWP30P140LVT U8466 ( .I(i_cmd[219]), .ZN(n7194) );
  OR2D1BWP30P140LVT U8467 ( .A1(i_cmd[211]), .A2(i_cmd[195]), .Z(n7193) );
  INVD1BWP30P140LVT U8468 ( .I(i_cmd[163]), .ZN(n6740) );
  ND2D1BWP30P140LVT U8469 ( .A1(n6740), .A2(n6742), .ZN(n6739) );
  INVD1BWP30P140LVT U8470 ( .I(i_cmd[179]), .ZN(n6742) );
  OR2D1BWP30P140LVT U8471 ( .A1(i_cmd[171]), .A2(i_cmd[187]), .Z(n6741) );
  INVD1BWP30P140LVT U8472 ( .I(i_cmd[155]), .ZN(n5954) );
  INVD1BWP30P140LVT U8473 ( .I(i_cmd[139]), .ZN(n5952) );
  OR2D1BWP30P140LVT U8474 ( .A1(i_cmd[131]), .A2(i_cmd[147]), .Z(n5953) );
  INVD1BWP30P140LVT U8475 ( .I(i_cmd[99]), .ZN(n6169) );
  ND2D1BWP30P140LVT U8476 ( .A1(n6169), .A2(n6168), .ZN(n6170) );
  INVD1BWP30P140LVT U8477 ( .I(i_cmd[115]), .ZN(n6168) );
  OR2D1BWP30P140LVT U8478 ( .A1(i_cmd[123]), .A2(i_cmd[107]), .Z(n6167) );
  INVD1BWP30P140LVT U8479 ( .I(i_cmd[91]), .ZN(n5940) );
  INVD1BWP30P140LVT U8480 ( .I(i_cmd[75]), .ZN(n5938) );
  OR2D1BWP30P140LVT U8481 ( .A1(i_cmd[67]), .A2(i_cmd[83]), .Z(n5939) );
  INVD1BWP30P140LVT U8482 ( .I(i_cmd[35]), .ZN(n6784) );
  INVD1BWP30P140LVT U8483 ( .I(i_cmd[51]), .ZN(n6783) );
  OR2D1BWP30P140LVT U8484 ( .A1(i_cmd[59]), .A2(i_cmd[43]), .Z(n6785) );
  ND2D1BWP30P140LVT U8485 ( .A1(n6783), .A2(n6784), .ZN(n6786) );
  INVD1BWP30P140LVT U8486 ( .I(i_cmd[3]), .ZN(n7312) );
  INVD1BWP30P140LVT U8487 ( .I(i_cmd[19]), .ZN(n7311) );
  OR2D1BWP30P140LVT U8488 ( .A1(i_cmd[27]), .A2(i_cmd[11]), .Z(n7313) );
  ND2D1BWP30P140LVT U8489 ( .A1(n7311), .A2(n7312), .ZN(n7314) );
  INVD1BWP30P140LVT U8490 ( .I(i_cmd[250]), .ZN(n7125) );
  INVD1BWP30P140LVT U8491 ( .I(i_cmd[234]), .ZN(n7127) );
  OR2D1BWP30P140LVT U8492 ( .A1(i_cmd[242]), .A2(i_cmd[226]), .Z(n7128) );
  ND2D1BWP30P140LVT U8493 ( .A1(n7127), .A2(n7125), .ZN(n7126) );
  INVD1BWP30P140LVT U8494 ( .I(i_cmd[202]), .ZN(n6358) );
  INVD1BWP30P140LVT U8495 ( .I(i_cmd[218]), .ZN(n6359) );
  OR2D1BWP30P140LVT U8496 ( .A1(i_cmd[210]), .A2(i_cmd[194]), .Z(n6360) );
  ND2D1BWP30P140LVT U8497 ( .A1(n6359), .A2(n6358), .ZN(n6357) );
  INVD1BWP30P140LVT U8498 ( .I(i_cmd[178]), .ZN(n6716) );
  ND2D1BWP30P140LVT U8499 ( .A1(n6716), .A2(n6718), .ZN(n6715) );
  INVD1BWP30P140LVT U8500 ( .I(i_cmd[162]), .ZN(n6718) );
  OR2D1BWP30P140LVT U8501 ( .A1(i_cmd[186]), .A2(i_cmd[170]), .Z(n6717) );
  INVD1BWP30P140LVT U8502 ( .I(i_cmd[154]), .ZN(n7156) );
  INVD1BWP30P140LVT U8503 ( .I(i_cmd[138]), .ZN(n7155) );
  OR2D1BWP30P140LVT U8504 ( .A1(i_cmd[146]), .A2(i_cmd[130]), .Z(n7157) );
  ND2D1BWP30P140LVT U8505 ( .A1(n7156), .A2(n7155), .ZN(n7158) );
  INVD1BWP30P140LVT U8506 ( .I(i_cmd[122]), .ZN(n5990) );
  INVD1BWP30P140LVT U8507 ( .I(i_cmd[106]), .ZN(n5988) );
  OR2D1BWP30P140LVT U8508 ( .A1(i_cmd[98]), .A2(i_cmd[114]), .Z(n5989) );
  INVD1BWP30P140LVT U8509 ( .I(i_cmd[90]), .ZN(n5980) );
  INVD1BWP30P140LVT U8510 ( .I(i_cmd[74]), .ZN(n5982) );
  OR2D1BWP30P140LVT U8511 ( .A1(i_cmd[66]), .A2(i_cmd[82]), .Z(n5981) );
  INVD1BWP30P140LVT U8512 ( .I(i_cmd[34]), .ZN(n6838) );
  ND2D1BWP30P140LVT U8513 ( .A1(n6838), .A2(n6840), .ZN(n6837) );
  INVD1BWP30P140LVT U8514 ( .I(i_cmd[50]), .ZN(n6840) );
  OR2D1BWP30P140LVT U8515 ( .A1(i_cmd[58]), .A2(i_cmd[42]), .Z(n6839) );
  INVD1BWP30P140LVT U8516 ( .I(i_cmd[2]), .ZN(n6582) );
  ND2D1BWP30P140LVT U8517 ( .A1(n6582), .A2(n6584), .ZN(n6581) );
  INVD1BWP30P140LVT U8518 ( .I(i_cmd[18]), .ZN(n6584) );
  OR2D1BWP30P140LVT U8519 ( .A1(i_cmd[26]), .A2(i_cmd[10]), .Z(n6583) );
  INVD1BWP30P140LVT U8520 ( .I(i_cmd[225]), .ZN(n6815) );
  INVD1BWP30P140LVT U8521 ( .I(i_cmd[241]), .ZN(n6817) );
  OR2D1BWP30P140LVT U8522 ( .A1(i_cmd[249]), .A2(i_cmd[233]), .Z(n6816) );
  ND2D1BWP30P140LVT U8523 ( .A1(n6815), .A2(n6817), .ZN(n6818) );
  INVD1BWP30P140LVT U8524 ( .I(i_cmd[201]), .ZN(n6442) );
  INVD1BWP30P140LVT U8525 ( .I(i_cmd[217]), .ZN(n6443) );
  OR2D1BWP30P140LVT U8526 ( .A1(i_cmd[209]), .A2(i_cmd[193]), .Z(n6444) );
  ND2D1BWP30P140LVT U8527 ( .A1(n6442), .A2(n6443), .ZN(n6441) );
  INVD1BWP30P140LVT U8528 ( .I(i_cmd[161]), .ZN(n7197) );
  INVD1BWP30P140LVT U8529 ( .I(i_cmd[177]), .ZN(n7198) );
  OR2D1BWP30P140LVT U8530 ( .A1(i_cmd[185]), .A2(i_cmd[169]), .Z(n7199) );
  ND2D1BWP30P140LVT U8531 ( .A1(n7197), .A2(n7198), .ZN(n7200) );
  INVD1BWP30P140LVT U8532 ( .I(i_cmd[153]), .ZN(n6509) );
  ND2D1BWP30P140LVT U8533 ( .A1(n6509), .A2(n6512), .ZN(n6510) );
  INVD1BWP30P140LVT U8534 ( .I(i_cmd[137]), .ZN(n6512) );
  OR2D1BWP30P140LVT U8535 ( .A1(i_cmd[145]), .A2(i_cmd[129]), .Z(n6511) );
  INVD1BWP30P140LVT U8536 ( .I(i_cmd[105]), .ZN(n6299) );
  ND2D1BWP30P140LVT U8537 ( .A1(n6299), .A2(n6302), .ZN(n6300) );
  INVD1BWP30P140LVT U8538 ( .I(i_cmd[121]), .ZN(n6302) );
  OR2D1BWP30P140LVT U8539 ( .A1(i_cmd[113]), .A2(i_cmd[97]), .Z(n6301) );
  INVD1BWP30P140LVT U8540 ( .I(i_cmd[81]), .ZN(n6399) );
  ND2D1BWP30P140LVT U8541 ( .A1(n6399), .A2(n6402), .ZN(n6400) );
  INVD1BWP30P140LVT U8542 ( .I(i_cmd[65]), .ZN(n6402) );
  OR2D1BWP30P140LVT U8543 ( .A1(i_cmd[89]), .A2(i_cmd[73]), .Z(n6401) );
  INVD1BWP30P140LVT U8544 ( .I(i_cmd[57]), .ZN(n5960) );
  INVD1BWP30P140LVT U8545 ( .I(i_cmd[41]), .ZN(n5958) );
  OR2D1BWP30P140LVT U8546 ( .A1(i_cmd[33]), .A2(i_cmd[49]), .Z(n5959) );
  INVD1BWP30P140LVT U8547 ( .I(i_cmd[25]), .ZN(n6619) );
  ND2D1BWP30P140LVT U8548 ( .A1(n6619), .A2(n6622), .ZN(n6620) );
  INVD1BWP30P140LVT U8549 ( .I(i_cmd[9]), .ZN(n6622) );
  OR2D1BWP30P140LVT U8550 ( .A1(i_cmd[17]), .A2(i_cmd[1]), .Z(n6621) );
  INVD1BWP30P140LVT U8551 ( .I(i_cmd[240]), .ZN(n10025) );
  ND2OPTIBD1BWP30P140LVT U8552 ( .A1(n5900), .A2(i_valid[30]), .ZN(n10024) );
  ND2OPTIBD1BWP30P140LVT U8553 ( .A1(n5900), .A2(i_valid[31]), .ZN(n10030) );
  ND2OPTIBD1BWP30P140LVT U8554 ( .A1(n5900), .A2(i_valid[29]), .ZN(n10023) );
  INVD1BWP30P140LVT U8555 ( .I(i_cmd[224]), .ZN(n10027) );
  ND2OPTIBD1BWP30P140LVT U8556 ( .A1(n5900), .A2(i_valid[28]), .ZN(n10028) );
  OR2D1BWP30P140LVT U8557 ( .A1(i_cmd[232]), .A2(i_cmd[248]), .Z(n10026) );
  INVD1BWP30P140LVT U8558 ( .I(i_cmd[192]), .ZN(n9745) );
  ND2OPTIBD1BWP30P140LVT U8559 ( .A1(n5900), .A2(i_valid[24]), .ZN(n9744) );
  ND2OPTIBD1BWP30P140LVT U8560 ( .A1(n5900), .A2(i_valid[25]), .ZN(n9743) );
  ND2OPTIBD1BWP30P140LVT U8561 ( .A1(n5900), .A2(i_valid[27]), .ZN(n9747) );
  ND2D1BWP30P140LVT U8562 ( .A1(n9742), .A2(n9745), .ZN(n9748) );
  INVD1BWP30P140LVT U8563 ( .I(i_cmd[208]), .ZN(n9742) );
  ND2OPTIBD1BWP30P140LVT U8564 ( .A1(n5900), .A2(i_valid[26]), .ZN(n9741) );
  OR2D1BWP30P140LVT U8565 ( .A1(i_cmd[200]), .A2(i_cmd[216]), .Z(n9746) );
  INVD1BWP30P140LVT U8566 ( .I(i_cmd[184]), .ZN(n9845) );
  ND2OPTIBD1BWP30P140LVT U8567 ( .A1(n5900), .A2(i_valid[23]), .ZN(n9844) );
  ND2OPTIBD1BWP30P140LVT U8568 ( .A1(n5900), .A2(i_valid[22]), .ZN(n9850) );
  ND2OPTIBD1BWP30P140LVT U8569 ( .A1(n5900), .A2(i_valid[20]), .ZN(n9843) );
  INVD1BWP30P140LVT U8570 ( .I(i_cmd[168]), .ZN(n9846) );
  ND2OPTIBD1BWP30P140LVT U8571 ( .A1(n5900), .A2(i_valid[21]), .ZN(n9847) );
  OR2D1BWP30P140LVT U8572 ( .A1(i_cmd[160]), .A2(i_cmd[176]), .Z(n9848) );
  INVD1BWP30P140LVT U8573 ( .I(i_cmd[144]), .ZN(n9835) );
  ND2OPTIBD1BWP30P140LVT U8574 ( .A1(n5900), .A2(i_valid[18]), .ZN(n9834) );
  INVD1BWP30P140LVT U8575 ( .I(i_cmd[128]), .ZN(n9840) );
  ND2OPTIBD1BWP30P140LVT U8576 ( .A1(n5900), .A2(i_valid[16]), .ZN(n9839) );
  OR2D1BWP30P140LVT U8577 ( .A1(i_cmd[152]), .A2(i_cmd[136]), .Z(n9838) );
  ND2OPTIBD1BWP30P140LVT U8578 ( .A1(n5900), .A2(i_valid[17]), .ZN(n9833) );
  ND2OPTIBD1BWP30P140LVT U8579 ( .A1(n5900), .A2(i_valid[19]), .ZN(n9837) );
  INVD1BWP30P140LVT U8580 ( .I(i_cmd[112]), .ZN(n9763) );
  ND2OPTIBD1BWP30P140LVT U8581 ( .A1(n5900), .A2(i_valid[14]), .ZN(n9761) );
  ND2OPTIBD1BWP30P140LVT U8582 ( .A1(n5900), .A2(i_valid[13]), .ZN(n9760) );
  ND2OPTIBD1BWP30P140LVT U8583 ( .A1(n5900), .A2(i_valid[15]), .ZN(n9764) );
  ND2D1BWP30P140LVT U8584 ( .A1(n9763), .A2(n9759), .ZN(n9765) );
  INVD1BWP30P140LVT U8585 ( .I(i_cmd[96]), .ZN(n9759) );
  ND2OPTIBD1BWP30P140LVT U8586 ( .A1(n5900), .A2(i_valid[12]), .ZN(n9758) );
  OR2D1BWP30P140LVT U8587 ( .A1(i_cmd[120]), .A2(i_cmd[104]), .Z(n9762) );
  INVD1BWP30P140LVT U8588 ( .I(i_cmd[64]), .ZN(n9810) );
  ND2OPTIBD1BWP30P140LVT U8589 ( .A1(n5900), .A2(i_valid[8]), .ZN(n9808) );
  INVD1BWP30P140LVT U8590 ( .I(i_cmd[80]), .ZN(n9811) );
  ND2OPTIBD1BWP30P140LVT U8591 ( .A1(n5900), .A2(i_valid[10]), .ZN(n9807) );
  OR2D1BWP30P140LVT U8592 ( .A1(i_cmd[88]), .A2(i_cmd[72]), .Z(n9809) );
  ND2OPTIBD1BWP30P140LVT U8593 ( .A1(n5900), .A2(i_valid[9]), .ZN(n9813) );
  ND2OPTIBD1BWP30P140LVT U8594 ( .A1(n5900), .A2(i_valid[11]), .ZN(n9812) );
  INVD1BWP30P140LVT U8595 ( .I(i_cmd[48]), .ZN(n9855) );
  ND2OPTIBD1BWP30P140LVT U8596 ( .A1(n5900), .A2(i_valid[6]), .ZN(n9854) );
  ND2OPTIBD1BWP30P140LVT U8597 ( .A1(n5900), .A2(i_valid[7]), .ZN(n9860) );
  ND2OPTIBD1BWP30P140LVT U8598 ( .A1(n5900), .A2(i_valid[5]), .ZN(n9853) );
  INVD1BWP30P140LVT U8599 ( .I(i_cmd[32]), .ZN(n9856) );
  ND2OPTIBD1BWP30P140LVT U8600 ( .A1(n5900), .A2(i_valid[4]), .ZN(n9857) );
  OR2D1BWP30P140LVT U8601 ( .A1(i_cmd[56]), .A2(i_cmd[40]), .Z(n9858) );
  INVD1BWP30P140LVT U8602 ( .I(i_cmd[16]), .ZN(n10017) );
  ND2OPTIBD1BWP30P140LVT U8603 ( .A1(n5900), .A2(i_valid[2]), .ZN(n10014) );
  INVD1BWP30P140LVT U8604 ( .I(i_cmd[0]), .ZN(n10016) );
  ND2OPTIBD1BWP30P140LVT U8605 ( .A1(n5900), .A2(i_valid[0]), .ZN(n10013) );
  OR2D1BWP30P140LVT U8606 ( .A1(i_cmd[8]), .A2(i_cmd[24]), .Z(n10015) );
  ND2OPTIBD1BWP30P140LVT U8607 ( .A1(n5900), .A2(i_valid[3]), .ZN(n10019) );
  ND2OPTIBD1BWP30P140LVT U8608 ( .A1(n5900), .A2(i_valid[1]), .ZN(n10018) );
  AN4D1BWP30P140LVT U8609 ( .A1(n5900), .A2(inner_first_stage_valid_reg[4]), 
        .A3(n5911), .A4(n5910), .Z(n10804) );
  AN3D1BWP30P140LVT U8610 ( .A1(inner_first_stage_valid_reg[5]), .A2(n5912), 
        .A3(n5908), .Z(n10803) );
  AN4D1BWP30P140LVT U8611 ( .A1(n5900), .A2(inner_first_stage_valid_reg[12]), 
        .A3(n10338), .A4(n10341), .Z(n10940) );
  AN4D1BWP30P140LVT U8612 ( .A1(n10342), .A2(inner_first_stage_valid_reg[9]), 
        .A3(n10339), .A4(n10340), .Z(n10939) );
  AN3D1BWP30P140LVT U8613 ( .A1(inner_first_stage_valid_reg[8]), .A2(n10341), 
        .A3(n10340), .Z(n10942) );
  NR3D0P7BWP30P140LVT U8614 ( .A1(inner_first_stage_valid_reg[27]), .A2(n10390), .A3(n10389), .ZN(n11211) );
  NR4D0BWP30P140LVT U8615 ( .A1(inner_first_stage_valid_reg[29]), .A2(
        inner_first_stage_valid_reg[25]), .A3(n10385), .A4(n10386), .ZN(n11214) );
  AN3D1BWP30P140LVT U8616 ( .A1(inner_first_stage_valid_reg[28]), .A2(n10388), 
        .A3(n10387), .Z(n11212) );
  NR3D0P7BWP30P140LVT U8617 ( .A1(inner_first_stage_valid_reg[26]), .A2(n10379), .A3(n10389), .ZN(n11216) );
  AN4D1BWP30P140LVT U8618 ( .A1(n5900), .A2(inner_first_stage_valid_reg[36]), 
        .A3(n6129), .A4(n6128), .Z(n11349) );
  AN3D1BWP30P140LVT U8619 ( .A1(n6125), .A2(inner_first_stage_valid_reg[37]), 
        .A3(n6124), .Z(n11348) );
  NR3D0P7BWP30P140LVT U8620 ( .A1(n10360), .A2(n10359), .A3(n10358), .ZN(
        n11483) );
  AN4D1BWP30P140LVT U8621 ( .A1(n5902), .A2(n5900), .A3(
        inner_first_stage_valid_reg[52]), .A4(n5901), .Z(n11619) );
  AN3D1BWP30P140LVT U8622 ( .A1(inner_first_stage_valid_reg[60]), .A2(n10302), 
        .A3(n10301), .Z(n11757) );
  NR3D0P7BWP30P140LVT U8623 ( .A1(inner_first_stage_valid_reg[63]), .A2(n10296), .A3(n10297), .ZN(n11762) );
  NR3D0P7BWP30P140LVT U8624 ( .A1(inner_first_stage_valid_reg[62]), .A2(n10298), .A3(n10297), .ZN(n11761) );
  ND2D1BWP30P140LVT U8625 ( .A1(n10377), .A2(n10376), .ZN(N5976) );
  ND2D1BWP30P140LVT U8626 ( .A1(n10362), .A2(n10361), .ZN(N11598) );
  ND2D1BWP30P140LVT U8627 ( .A1(n10306), .A2(n10305), .ZN(N15346) );
  ND2D1BWP30P140LVT U8628 ( .A1(n10332), .A2(n10331), .ZN(N2085) );
  ND2D1BWP30P140LVT U8629 ( .A1(n10310), .A2(n10309), .ZN(N2088) );
  ND2D1BWP30P140LVT U8630 ( .A1(n10308), .A2(n10307), .ZN(N2091) );
  ND2D1BWP30P140LVT U8631 ( .A1(n10328), .A2(n10327), .ZN(N2092) );
  ND2D1BWP30P140LVT U8632 ( .A1(n10314), .A2(n10313), .ZN(N2093) );
  ND2D1BWP30P140LVT U8633 ( .A1(n10312), .A2(n10311), .ZN(N2096) );
  ND2D1BWP30P140LVT U8634 ( .A1(n10318), .A2(n10317), .ZN(N2101) );
  ND2D1BWP30P140LVT U8635 ( .A1(n10316), .A2(n10315), .ZN(N2103) );
  ND2D1BWP30P140LVT U8636 ( .A1(n10330), .A2(n10329), .ZN(N2104) );
  ND2D1BWP30P140LVT U8637 ( .A1(n10326), .A2(n10325), .ZN(N2108) );
  ND2D1BWP30P140LVT U8638 ( .A1(n10324), .A2(n10323), .ZN(N2109) );
  ND2D1BWP30P140LVT U8639 ( .A1(n10320), .A2(n10319), .ZN(N2111) );
  ND2D1BWP30P140LVT U8640 ( .A1(n10322), .A2(n10321), .ZN(N2112) );
  ND2D1BWP30P140LVT U8641 ( .A1(n10222), .A2(n10221), .ZN(N1647) );
  ND2D1BWP30P140LVT U8642 ( .A1(n10228), .A2(n10227), .ZN(N1651) );
  ND2D1BWP30P140LVT U8643 ( .A1(n10224), .A2(n10223), .ZN(N1653) );
  ND2D1BWP30P140LVT U8644 ( .A1(n10226), .A2(n10225), .ZN(N1656) );
  ND2D1BWP30P140LVT U8645 ( .A1(n10204), .A2(n10203), .ZN(N1659) );
  ND2D1BWP30P140LVT U8646 ( .A1(n10220), .A2(n10219), .ZN(N1660) );
  ND2D1BWP30P140LVT U8647 ( .A1(n10212), .A2(n10211), .ZN(N1662) );
  ND2D1BWP30P140LVT U8648 ( .A1(n10214), .A2(n10213), .ZN(N1664) );
  ND2D1BWP30P140LVT U8649 ( .A1(n10208), .A2(n10207), .ZN(N1665) );
  ND2D1BWP30P140LVT U8650 ( .A1(n10206), .A2(n10205), .ZN(N1668) );
  ND2D1BWP30P140LVT U8651 ( .A1(n10210), .A2(n10209), .ZN(N1670) );
  ND2D1BWP30P140LVT U8652 ( .A1(n10216), .A2(n10215), .ZN(N1671) );
  ND2D1BWP30P140LVT U8653 ( .A1(n10218), .A2(n10217), .ZN(N1673) );
  ND2D1BWP30P140LVT U8654 ( .A1(n10196), .A2(n10195), .ZN(N1424) );
  ND2D1BWP30P140LVT U8655 ( .A1(n10194), .A2(n10193), .ZN(N1425) );
  ND2D1BWP30P140LVT U8656 ( .A1(n10192), .A2(n10191), .ZN(N1426) );
  ND2D1BWP30P140LVT U8657 ( .A1(n10202), .A2(n10201), .ZN(N1434) );
  ND2D1BWP30P140LVT U8658 ( .A1(n10178), .A2(n10177), .ZN(N1441) );
  ND2D1BWP30P140LVT U8659 ( .A1(n10200), .A2(n10199), .ZN(N1444) );
  ND2D1BWP30P140LVT U8660 ( .A1(n10176), .A2(n10175), .ZN(N1446) );
  ND2D1BWP30P140LVT U8661 ( .A1(n10172), .A2(n10171), .ZN(N1447) );
  ND2D1BWP30P140LVT U8662 ( .A1(n10180), .A2(n10179), .ZN(N1452) );
  ND2D1BWP30P140LVT U8663 ( .A1(n10182), .A2(n10181), .ZN(N1454) );
  ND2D1BWP30P140LVT U8664 ( .A1(n10234), .A2(n10233), .ZN(N765) );
  ND2D1BWP30P140LVT U8665 ( .A1(n10248), .A2(n10247), .ZN(N769) );
  ND2D1BWP30P140LVT U8666 ( .A1(n10236), .A2(n10235), .ZN(N771) );
  ND2D1BWP30P140LVT U8667 ( .A1(n10230), .A2(n10229), .ZN(N772) );
  ND2D1BWP30P140LVT U8668 ( .A1(n10254), .A2(n10253), .ZN(N774) );
  ND2D1BWP30P140LVT U8669 ( .A1(n10232), .A2(n10231), .ZN(N775) );
  ND2D1BWP30P140LVT U8670 ( .A1(n10244), .A2(n10243), .ZN(N776) );
  ND2D1BWP30P140LVT U8671 ( .A1(n10238), .A2(n10237), .ZN(N778) );
  ND2D1BWP30P140LVT U8672 ( .A1(n10258), .A2(n10257), .ZN(N779) );
  ND2D1BWP30P140LVT U8673 ( .A1(n10240), .A2(n10239), .ZN(N780) );
  ND2D1BWP30P140LVT U8674 ( .A1(n10242), .A2(n10241), .ZN(N785) );
  ND2D1BWP30P140LVT U8675 ( .A1(n10246), .A2(n10245), .ZN(N787) );
  ND2D1BWP30P140LVT U8676 ( .A1(n10250), .A2(n10249), .ZN(N792) );
  ND2D1BWP30P140LVT U8677 ( .A1(n10252), .A2(n10251), .ZN(N793) );
  ND2D1BWP30P140LVT U8678 ( .A1(n10256), .A2(n10255), .ZN(N794) );
  ND2D1BWP30P140LVT U8679 ( .A1(n10292), .A2(n10291), .ZN(N545) );
  ND2D1BWP30P140LVT U8680 ( .A1(n10286), .A2(n10285), .ZN(N546) );
  ND2D1BWP30P140LVT U8681 ( .A1(n10270), .A2(n10269), .ZN(N548) );
  ND2D1BWP30P140LVT U8682 ( .A1(n10274), .A2(n10273), .ZN(N550) );
  ND2D1BWP30P140LVT U8683 ( .A1(n10272), .A2(n10271), .ZN(N552) );
  ND2D1BWP30P140LVT U8684 ( .A1(n10266), .A2(n10265), .ZN(N553) );
  ND2D1BWP30P140LVT U8685 ( .A1(n10264), .A2(n10263), .ZN(N554) );
  ND2D1BWP30P140LVT U8686 ( .A1(n10262), .A2(n10261), .ZN(N555) );
  ND2D1BWP30P140LVT U8687 ( .A1(n10260), .A2(n10259), .ZN(N556) );
  ND2D1BWP30P140LVT U8688 ( .A1(n10290), .A2(n10289), .ZN(N561) );
  ND2D1BWP30P140LVT U8689 ( .A1(n10284), .A2(n10283), .ZN(N562) );
  ND2D1BWP30P140LVT U8690 ( .A1(n10268), .A2(n10267), .ZN(N565) );
  ND2D1BWP30P140LVT U8691 ( .A1(n10280), .A2(n10279), .ZN(N568) );
  ND2D1BWP30P140LVT U8692 ( .A1(n10278), .A2(n10277), .ZN(N569) );
  ND2D1BWP30P140LVT U8693 ( .A1(n10276), .A2(n10275), .ZN(N572) );
  ND2D1BWP30P140LVT U8694 ( .A1(n10288), .A2(n10287), .ZN(N573) );
  ND2D1BWP30P140LVT U8695 ( .A1(n10282), .A2(n10281), .ZN(N574) );
  INR4D1BWP30P140LVT U8696 ( .A1(inner_first_stage_valid_reg[33]), .B1(
        inner_first_stage_valid_reg[37]), .B2(inner_first_stage_valid_reg[32]), 
        .B3(n6130), .ZN(n11339) );
  INR4D1BWP30P140LVT U8697 ( .A1(i_cmd[216]), .B1(i_cmd[200]), .B2(n9748), 
        .B3(n9747), .ZN(n9749) );
  INR4D1BWP30P140LVT U8698 ( .A1(i_cmd[120]), .B1(i_cmd[104]), .B2(n9765), 
        .B3(n9764), .ZN(n9766) );
  NR2D1BWP30P140LVT U8699 ( .A1(inner_first_stage_valid_reg[54]), .A2(
        inner_first_stage_valid_reg[55]), .ZN(n5894) );
  NR3D0P7BWP30P140LVT U8700 ( .A1(inner_first_stage_valid_reg[51]), .A2(
        inner_first_stage_valid_reg[49]), .A3(inner_first_stage_valid_reg[53]), 
        .ZN(n5902) );
  INR3D0BWP30P140LVT U8701 ( .A1(n5902), .B1(inner_first_stage_valid_reg[52]), 
        .B2(n10380), .ZN(n5895) );
  INR3D2BWP30P140LVT U8702 ( .A1(inner_first_stage_valid_reg[50]), .B1(
        inner_first_stage_valid_reg[48]), .B2(n5903), .ZN(n11624) );
  NR2D1BWP30P140LVT U8703 ( .A1(inner_first_stage_valid_reg[50]), .A2(
        inner_first_stage_valid_reg[48]), .ZN(n5896) );
  INR3D2BWP30P140LVT U8704 ( .A1(inner_first_stage_valid_reg[54]), .B1(
        inner_first_stage_valid_reg[55]), .B2(n5897), .ZN(n11626) );
  INR3D2BWP30P140LVT U8705 ( .A1(inner_first_stage_valid_reg[55]), .B1(
        inner_first_stage_valid_reg[54]), .B2(n5897), .ZN(n11625) );
  NR4D0BWP30P140LVT U8706 ( .A1(inner_first_stage_valid_reg[54]), .A2(
        inner_first_stage_valid_reg[55]), .A3(inner_first_stage_valid_reg[50]), 
        .A4(inner_first_stage_valid_reg[48]), .ZN(n5901) );
  INR3D2BWP30P140LVT U8707 ( .A1(inner_first_stage_valid_reg[49]), .B1(
        inner_first_stage_valid_reg[53]), .B2(n5904), .ZN(n11623) );
  NR4D0BWP30P140LVT U8708 ( .A1(n11624), .A2(n11626), .A3(n11625), .A4(n11623), 
        .ZN(n5906) );
  INR4D1BWP30P140LVT U8709 ( .A1(inner_first_stage_valid_reg[51]), .B1(
        inner_first_stage_valid_reg[53]), .B2(inner_first_stage_valid_reg[49]), 
        .B3(n5899), .ZN(n11620) );
  INR3D2BWP30P140LVT U8710 ( .A1(inner_first_stage_valid_reg[48]), .B1(
        inner_first_stage_valid_reg[50]), .B2(n5903), .ZN(n11622) );
  INR3D2BWP30P140LVT U8711 ( .A1(inner_first_stage_valid_reg[53]), .B1(
        inner_first_stage_valid_reg[49]), .B2(n5904), .ZN(n11621) );
  NR4D0BWP30P140LVT U8712 ( .A1(n11620), .A2(n11619), .A3(n11622), .A4(n11621), 
        .ZN(n5905) );
  ND2D1BWP30P140LVT U8713 ( .A1(n5906), .A2(n5905), .ZN(N13472) );
  INR4D0BWP30P140LVT U8714 ( .A1(n5914), .B1(inner_first_stage_valid_reg[1]), 
        .B2(inner_first_stage_valid_reg[5]), .B3(
        inner_first_stage_valid_reg[0]), .ZN(n5910) );
  INR3D2BWP30P140LVT U8715 ( .A1(inner_first_stage_valid_reg[7]), .B1(
        inner_first_stage_valid_reg[6]), .B2(n5909), .ZN(n10805) );
  NR3D0P7BWP30P140LVT U8716 ( .A1(inner_first_stage_valid_reg[2]), .A2(
        inner_first_stage_valid_reg[3]), .A3(inner_first_stage_valid_reg[1]), 
        .ZN(n5908) );
  INR3D2BWP30P140LVT U8717 ( .A1(inner_first_stage_valid_reg[6]), .B1(
        inner_first_stage_valid_reg[7]), .B2(n5909), .ZN(n10802) );
  NR4D0BWP30P140LVT U8718 ( .A1(n10805), .A2(n10803), .A3(n10802), .A4(n10804), 
        .ZN(n5919) );
  NR2D1BWP30P140LVT U8719 ( .A1(inner_first_stage_valid_reg[1]), .A2(
        inner_first_stage_valid_reg[5]), .ZN(n5913) );
  INR3D2BWP30P140LVT U8720 ( .A1(inner_first_stage_valid_reg[2]), .B1(
        inner_first_stage_valid_reg[3]), .B2(n5917), .ZN(n10814) );
  INR4D1BWP30P140LVT U8721 ( .A1(inner_first_stage_valid_reg[0]), .B1(
        inner_first_stage_valid_reg[1]), .B2(inner_first_stage_valid_reg[5]), 
        .B3(n5916), .ZN(n10808) );
  INR4D1BWP30P140LVT U8722 ( .A1(inner_first_stage_valid_reg[1]), .B1(
        inner_first_stage_valid_reg[0]), .B2(inner_first_stage_valid_reg[5]), 
        .B3(n5916), .ZN(n10807) );
  INR3D2BWP30P140LVT U8723 ( .A1(inner_first_stage_valid_reg[3]), .B1(
        inner_first_stage_valid_reg[2]), .B2(n5917), .ZN(n10806) );
  NR4D0BWP30P140LVT U8724 ( .A1(n10814), .A2(n10808), .A3(n10807), .A4(n10806), 
        .ZN(n5918) );
  ND2D1BWP30P140LVT U8725 ( .A1(n5919), .A2(n5918), .ZN(N2228) );
  NR4D1BWP30P140LVT U8726 ( .A1(i_cmd[229]), .A2(n5920), .A3(n10024), .A4(
        n5921), .ZN(n10459) );
  INR4D1BWP30P140LVT U8727 ( .A1(i_cmd[253]), .B1(i_cmd[237]), .B2(n5923), 
        .B3(n10030), .ZN(n10457) );
  AOI22D1BWP30P140LVT U8728 ( .A1(i_data_bus[985]), .A2(n10459), .B1(
        i_data_bus[1017]), .B2(n10457), .ZN(n5925) );
  NR4D1BWP30P140LVT U8729 ( .A1(i_cmd[245]), .A2(n10028), .A3(n5922), .A4(
        n5921), .ZN(n10458) );
  INR4D1BWP30P140LVT U8730 ( .A1(i_cmd[237]), .B1(i_cmd[253]), .B2(n5923), 
        .B3(n10023), .ZN(n10460) );
  AOI22D1BWP30P140LVT U8731 ( .A1(i_data_bus[921]), .A2(n10458), .B1(
        i_data_bus[953]), .B2(n10460), .ZN(n5924) );
  ND2D1BWP30P140LVT U8732 ( .A1(n5925), .A2(n5924), .ZN(N11478) );
  AOI22D1BWP30P140LVT U8733 ( .A1(i_data_bus[970]), .A2(n10459), .B1(
        i_data_bus[1002]), .B2(n10457), .ZN(n5927) );
  AOI22D1BWP30P140LVT U8734 ( .A1(i_data_bus[906]), .A2(n10458), .B1(
        i_data_bus[938]), .B2(n10460), .ZN(n5926) );
  ND2D1BWP30P140LVT U8735 ( .A1(n5927), .A2(n5926), .ZN(N11463) );
  NR4D1BWP30P140LVT U8736 ( .A1(i_cmd[230]), .A2(n5928), .A3(n10024), .A4(
        n5929), .ZN(n10426) );
  INR4D1BWP30P140LVT U8737 ( .A1(i_cmd[254]), .B1(i_cmd[238]), .B2(n5931), 
        .B3(n10030), .ZN(n10427) );
  AOI22D1BWP30P140LVT U8738 ( .A1(i_data_bus[985]), .A2(n10426), .B1(
        i_data_bus[1017]), .B2(n10427), .ZN(n5933) );
  NR4D1BWP30P140LVT U8739 ( .A1(i_cmd[246]), .A2(n10028), .A3(n5930), .A4(
        n5929), .ZN(n10425) );
  INR4D1BWP30P140LVT U8740 ( .A1(i_cmd[238]), .B1(i_cmd[254]), .B2(n5931), 
        .B3(n10023), .ZN(n10428) );
  AOI22D1BWP30P140LVT U8741 ( .A1(i_data_bus[921]), .A2(n10425), .B1(
        i_data_bus[953]), .B2(n10428), .ZN(n5932) );
  ND2D1BWP30P140LVT U8742 ( .A1(n5933), .A2(n5932), .ZN(N13352) );
  AOI22D1BWP30P140LVT U8743 ( .A1(i_data_bus[969]), .A2(n10426), .B1(
        i_data_bus[1001]), .B2(n10427), .ZN(n5935) );
  AOI22D1BWP30P140LVT U8744 ( .A1(i_data_bus[905]), .A2(n10425), .B1(
        i_data_bus[937]), .B2(n10428), .ZN(n5934) );
  ND2D1BWP30P140LVT U8745 ( .A1(n5935), .A2(n5934), .ZN(N13336) );
  AOI22D1BWP30P140LVT U8746 ( .A1(i_data_bus[917]), .A2(n10425), .B1(
        i_data_bus[1013]), .B2(n10427), .ZN(n5937) );
  AOI22D1BWP30P140LVT U8747 ( .A1(i_data_bus[981]), .A2(n10426), .B1(
        i_data_bus[949]), .B2(n10428), .ZN(n5936) );
  ND2D1BWP30P140LVT U8748 ( .A1(n5937), .A2(n5936), .ZN(N13348) );
  NR4D1BWP30P140LVT U8749 ( .A1(i_cmd[91]), .A2(n9813), .A3(n5938), .A4(n5939), 
        .ZN(n10541) );
  INR4D1BWP30P140LVT U8750 ( .A1(i_cmd[83]), .B1(i_cmd[67]), .B2(n5941), .B3(
        n9807), .ZN(n10544) );
  AOI22D1BWP30P140LVT U8751 ( .A1(i_data_bus[295]), .A2(n10541), .B1(
        i_data_bus[327]), .B2(n10544), .ZN(n5943) );
  NR4D1BWP30P140LVT U8752 ( .A1(i_cmd[75]), .A2(n5940), .A3(n9812), .A4(n5939), 
        .ZN(n10542) );
  INR4D1BWP30P140LVT U8753 ( .A1(i_cmd[67]), .B1(i_cmd[83]), .B2(n5941), .B3(
        n9808), .ZN(n10543) );
  AOI22D1BWP30P140LVT U8754 ( .A1(i_data_bus[359]), .A2(n10542), .B1(
        i_data_bus[263]), .B2(n10543), .ZN(n5942) );
  ND2D1BWP30P140LVT U8755 ( .A1(n5943), .A2(n5942), .ZN(N6632) );
  AOI22D1BWP30P140LVT U8756 ( .A1(i_data_bus[355]), .A2(n10542), .B1(
        i_data_bus[323]), .B2(n10544), .ZN(n5945) );
  AOI22D1BWP30P140LVT U8757 ( .A1(i_data_bus[291]), .A2(n10541), .B1(
        i_data_bus[259]), .B2(n10543), .ZN(n5944) );
  ND2D1BWP30P140LVT U8758 ( .A1(n5945), .A2(n5944), .ZN(N6628) );
  NR4D1BWP30P140LVT U8759 ( .A1(i_cmd[143]), .A2(n5946), .A3(n9837), .A4(n5947), .ZN(n10407) );
  INR4D1BWP30P140LVT U8760 ( .A1(i_cmd[151]), .B1(i_cmd[135]), .B2(n5949), 
        .B3(n9834), .ZN(n10408) );
  AOI22D1BWP30P140LVT U8761 ( .A1(i_data_bus[616]), .A2(n10407), .B1(
        i_data_bus[584]), .B2(n10408), .ZN(n5951) );
  NR4D1BWP30P140LVT U8762 ( .A1(i_cmd[159]), .A2(n9833), .A3(n5948), .A4(n5947), .ZN(n10406) );
  INR4D1BWP30P140LVT U8763 ( .A1(i_cmd[135]), .B1(i_cmd[151]), .B2(n5949), 
        .B3(n9839), .ZN(n10405) );
  AOI22D1BWP30P140LVT U8764 ( .A1(i_data_bus[552]), .A2(n10406), .B1(
        i_data_bus[520]), .B2(n10405), .ZN(n5950) );
  ND2D1BWP30P140LVT U8765 ( .A1(n5951), .A2(n5950), .ZN(N14561) );
  NR4D1BWP30P140LVT U8766 ( .A1(i_cmd[155]), .A2(n9833), .A3(n5952), .A4(n5953), .ZN(n10535) );
  INR4D1BWP30P140LVT U8767 ( .A1(i_cmd[147]), .B1(i_cmd[131]), .B2(n5955), 
        .B3(n9834), .ZN(n10536) );
  AOI22D1BWP30P140LVT U8768 ( .A1(i_data_bus[571]), .A2(n10535), .B1(
        i_data_bus[603]), .B2(n10536), .ZN(n5957) );
  NR4D1BWP30P140LVT U8769 ( .A1(i_cmd[139]), .A2(n5954), .A3(n9837), .A4(n5953), .ZN(n10534) );
  INR4D1BWP30P140LVT U8770 ( .A1(i_cmd[131]), .B1(i_cmd[147]), .B2(n5955), 
        .B3(n9839), .ZN(n10533) );
  AOI22D1BWP30P140LVT U8771 ( .A1(i_data_bus[635]), .A2(n10534), .B1(
        i_data_bus[539]), .B2(n10533), .ZN(n5956) );
  ND2D1BWP30P140LVT U8772 ( .A1(n5957), .A2(n5956), .ZN(N7084) );
  NR4D1BWP30P140LVT U8773 ( .A1(i_cmd[57]), .A2(n9853), .A3(n5958), .A4(n5959), 
        .ZN(n10609) );
  INR4D1BWP30P140LVT U8774 ( .A1(i_cmd[33]), .B1(i_cmd[49]), .B2(n5961), .B3(
        n9857), .ZN(n10612) );
  AOI22D1BWP30P140LVT U8775 ( .A1(i_data_bus[170]), .A2(n10609), .B1(
        i_data_bus[138]), .B2(n10612), .ZN(n5963) );
  NR4D1BWP30P140LVT U8776 ( .A1(i_cmd[41]), .A2(n5960), .A3(n9860), .A4(n5959), 
        .ZN(n10611) );
  INR4D1BWP30P140LVT U8777 ( .A1(i_cmd[49]), .B1(i_cmd[33]), .B2(n5961), .B3(
        n9854), .ZN(n10610) );
  AOI22D1BWP30P140LVT U8778 ( .A1(i_data_bus[234]), .A2(n10611), .B1(
        i_data_bus[202]), .B2(n10610), .ZN(n5962) );
  ND2D1BWP30P140LVT U8779 ( .A1(n5963), .A2(n5962), .ZN(N2671) );
  AOI22D1BWP30P140LVT U8780 ( .A1(i_data_bus[172]), .A2(n10609), .B1(
        i_data_bus[140]), .B2(n10612), .ZN(n5965) );
  AOI22D1BWP30P140LVT U8781 ( .A1(i_data_bus[236]), .A2(n10611), .B1(
        i_data_bus[204]), .B2(n10610), .ZN(n5964) );
  ND2D1BWP30P140LVT U8782 ( .A1(n5965), .A2(n5964), .ZN(N2673) );
  AOI22D1BWP30P140LVT U8783 ( .A1(i_data_bus[231]), .A2(n10611), .B1(
        i_data_bus[135]), .B2(n10612), .ZN(n5967) );
  AOI22D1BWP30P140LVT U8784 ( .A1(i_data_bus[167]), .A2(n10609), .B1(
        i_data_bus[199]), .B2(n10610), .ZN(n5966) );
  ND2D1BWP30P140LVT U8785 ( .A1(n5967), .A2(n5966), .ZN(N2668) );
  AOI22D1BWP30P140LVT U8786 ( .A1(i_data_bus[227]), .A2(n10611), .B1(
        i_data_bus[131]), .B2(n10612), .ZN(n5969) );
  AOI22D1BWP30P140LVT U8787 ( .A1(i_data_bus[163]), .A2(n10609), .B1(
        i_data_bus[195]), .B2(n10610), .ZN(n5968) );
  ND2D1BWP30P140LVT U8788 ( .A1(n5969), .A2(n5968), .ZN(N2664) );
  AOI22D1BWP30P140LVT U8789 ( .A1(i_data_bus[186]), .A2(n10609), .B1(
        i_data_bus[154]), .B2(n10612), .ZN(n5971) );
  AOI22D1BWP30P140LVT U8790 ( .A1(i_data_bus[250]), .A2(n10611), .B1(
        i_data_bus[218]), .B2(n10610), .ZN(n5970) );
  ND2D1BWP30P140LVT U8791 ( .A1(n5971), .A2(n5970), .ZN(N2687) );
  AOI22D1BWP30P140LVT U8792 ( .A1(i_data_bus[916]), .A2(n10425), .B1(
        i_data_bus[948]), .B2(n10428), .ZN(n5973) );
  AOI22D1BWP30P140LVT U8793 ( .A1(i_data_bus[980]), .A2(n10426), .B1(
        i_data_bus[1012]), .B2(n10427), .ZN(n5972) );
  ND2D1BWP30P140LVT U8794 ( .A1(n5973), .A2(n5972), .ZN(N13347) );
  AOI22D1BWP30P140LVT U8795 ( .A1(i_data_bus[924]), .A2(n10425), .B1(
        i_data_bus[956]), .B2(n10428), .ZN(n5975) );
  AOI22D1BWP30P140LVT U8796 ( .A1(i_data_bus[988]), .A2(n10426), .B1(
        i_data_bus[1020]), .B2(n10427), .ZN(n5974) );
  ND2D1BWP30P140LVT U8797 ( .A1(n5975), .A2(n5974), .ZN(N13355) );
  AOI22D1BWP30P140LVT U8798 ( .A1(i_data_bus[989]), .A2(n10426), .B1(
        i_data_bus[957]), .B2(n10428), .ZN(n5977) );
  AOI22D1BWP30P140LVT U8799 ( .A1(i_data_bus[925]), .A2(n10425), .B1(
        i_data_bus[1021]), .B2(n10427), .ZN(n5976) );
  ND2D1BWP30P140LVT U8800 ( .A1(n5977), .A2(n5976), .ZN(N13356) );
  AOI22D1BWP30P140LVT U8801 ( .A1(i_data_bus[906]), .A2(n10425), .B1(
        i_data_bus[938]), .B2(n10428), .ZN(n5979) );
  AOI22D1BWP30P140LVT U8802 ( .A1(i_data_bus[970]), .A2(n10426), .B1(
        i_data_bus[1002]), .B2(n10427), .ZN(n5978) );
  ND2D1BWP30P140LVT U8803 ( .A1(n5979), .A2(n5978), .ZN(N13337) );
  NR4D1BWP30P140LVT U8804 ( .A1(i_cmd[74]), .A2(n5980), .A3(n9812), .A4(n5981), 
        .ZN(n10574) );
  INR4D1BWP30P140LVT U8805 ( .A1(i_cmd[82]), .B1(i_cmd[66]), .B2(n5983), .B3(
        n9807), .ZN(n10576) );
  AOI22D1BWP30P140LVT U8806 ( .A1(i_data_bus[372]), .A2(n10574), .B1(
        i_data_bus[340]), .B2(n10576), .ZN(n5985) );
  NR4D1BWP30P140LVT U8807 ( .A1(i_cmd[90]), .A2(n9813), .A3(n5982), .A4(n5981), 
        .ZN(n10573) );
  INR4D1BWP30P140LVT U8808 ( .A1(i_cmd[66]), .B1(i_cmd[82]), .B2(n5983), .B3(
        n9808), .ZN(n10575) );
  AOI22D1BWP30P140LVT U8809 ( .A1(i_data_bus[308]), .A2(n10573), .B1(
        i_data_bus[276]), .B2(n10575), .ZN(n5984) );
  ND2D1BWP30P140LVT U8810 ( .A1(n5985), .A2(n5984), .ZN(N4771) );
  AOI22D1BWP30P140LVT U8811 ( .A1(i_data_bus[369]), .A2(n10574), .B1(
        i_data_bus[337]), .B2(n10576), .ZN(n5987) );
  AOI22D1BWP30P140LVT U8812 ( .A1(i_data_bus[305]), .A2(n10573), .B1(
        i_data_bus[273]), .B2(n10575), .ZN(n5986) );
  ND2D1BWP30P140LVT U8813 ( .A1(n5987), .A2(n5986), .ZN(N4768) );
  NR4D1BWP30P140LVT U8814 ( .A1(i_cmd[122]), .A2(n9760), .A3(n5988), .A4(n5989), .ZN(n10569) );
  INR4D1BWP30P140LVT U8815 ( .A1(i_cmd[98]), .B1(i_cmd[114]), .B2(n5991), .B3(
        n9758), .ZN(n10572) );
  AOI22D1BWP30P140LVT U8816 ( .A1(i_data_bus[431]), .A2(n10569), .B1(
        i_data_bus[399]), .B2(n10572), .ZN(n5993) );
  NR4D1BWP30P140LVT U8817 ( .A1(i_cmd[106]), .A2(n5990), .A3(n9764), .A4(n5989), .ZN(n10571) );
  INR4D1BWP30P140LVT U8818 ( .A1(i_cmd[114]), .B1(i_cmd[98]), .B2(n5991), .B3(
        n9761), .ZN(n10570) );
  AOI22D1BWP30P140LVT U8819 ( .A1(i_data_bus[495]), .A2(n10571), .B1(
        i_data_bus[463]), .B2(n10570), .ZN(n5992) );
  ND2D1BWP30P140LVT U8820 ( .A1(n5993), .A2(n5992), .ZN(N4982) );
  AOI22D1BWP30P140LVT U8821 ( .A1(i_data_bus[498]), .A2(n10571), .B1(
        i_data_bus[402]), .B2(n10572), .ZN(n5995) );
  AOI22D1BWP30P140LVT U8822 ( .A1(i_data_bus[434]), .A2(n10569), .B1(
        i_data_bus[466]), .B2(n10570), .ZN(n5994) );
  ND2D1BWP30P140LVT U8823 ( .A1(n5995), .A2(n5994), .ZN(N4985) );
  NR4D1BWP30P140LVT U8824 ( .A1(i_cmd[183]), .A2(n9843), .A3(n5996), .A4(n5997), .ZN(n10401) );
  INR4D1BWP30P140LVT U8825 ( .A1(i_cmd[191]), .B1(i_cmd[175]), .B2(n5999), 
        .B3(n9844), .ZN(n10403) );
  AOI22D1BWP30P140LVT U8826 ( .A1(i_data_bus[658]), .A2(n10401), .B1(
        i_data_bus[754]), .B2(n10403), .ZN(n6001) );
  NR4D1BWP30P140LVT U8827 ( .A1(i_cmd[167]), .A2(n5998), .A3(n9850), .A4(n5997), .ZN(n10402) );
  INR4D1BWP30P140LVT U8828 ( .A1(i_cmd[175]), .B1(i_cmd[191]), .B2(n5999), 
        .B3(n9847), .ZN(n10404) );
  AOI22D1BWP30P140LVT U8829 ( .A1(i_data_bus[722]), .A2(n10402), .B1(
        i_data_bus[690]), .B2(n10404), .ZN(n6000) );
  ND2D1BWP30P140LVT U8830 ( .A1(n6001), .A2(n6000), .ZN(N14787) );
  AOI22D1BWP30P140LVT U8831 ( .A1(i_data_bus[379]), .A2(n10574), .B1(
        i_data_bus[283]), .B2(n10575), .ZN(n6003) );
  AOI22D1BWP30P140LVT U8832 ( .A1(i_data_bus[315]), .A2(n10573), .B1(
        i_data_bus[347]), .B2(n10576), .ZN(n6002) );
  ND2D1BWP30P140LVT U8833 ( .A1(n6003), .A2(n6002), .ZN(N4778) );
  AOI22D1BWP30P140LVT U8834 ( .A1(i_data_bus[355]), .A2(n10574), .B1(
        i_data_bus[259]), .B2(n10575), .ZN(n6005) );
  AOI22D1BWP30P140LVT U8835 ( .A1(i_data_bus[291]), .A2(n10573), .B1(
        i_data_bus[323]), .B2(n10576), .ZN(n6004) );
  ND2D1BWP30P140LVT U8836 ( .A1(n6005), .A2(n6004), .ZN(N4754) );
  AOI22D1BWP30P140LVT U8837 ( .A1(i_data_bus[733]), .A2(n10402), .B1(
        i_data_bus[765]), .B2(n10403), .ZN(n6007) );
  AOI22D1BWP30P140LVT U8838 ( .A1(i_data_bus[669]), .A2(n10401), .B1(
        i_data_bus[701]), .B2(n10404), .ZN(n6006) );
  ND2D1BWP30P140LVT U8839 ( .A1(n6007), .A2(n6006), .ZN(N14798) );
  AOI22D1BWP30P140LVT U8840 ( .A1(i_data_bus[358]), .A2(n10574), .B1(
        i_data_bus[262]), .B2(n10575), .ZN(n6009) );
  AOI22D1BWP30P140LVT U8841 ( .A1(i_data_bus[294]), .A2(n10573), .B1(
        i_data_bus[326]), .B2(n10576), .ZN(n6008) );
  ND2D1BWP30P140LVT U8842 ( .A1(n6009), .A2(n6008), .ZN(N4757) );
  NR4D1BWP30P140LVT U8843 ( .A1(i_cmd[165]), .A2(n6010), .A3(n9850), .A4(n6011), .ZN(n10465) );
  INR4D1BWP30P140LVT U8844 ( .A1(i_cmd[173]), .B1(i_cmd[189]), .B2(n6013), 
        .B3(n9847), .ZN(n10468) );
  AOI22D1BWP30P140LVT U8845 ( .A1(i_data_bus[733]), .A2(n10465), .B1(
        i_data_bus[701]), .B2(n10468), .ZN(n6015) );
  NR4D1BWP30P140LVT U8846 ( .A1(i_cmd[181]), .A2(n9843), .A3(n6012), .A4(n6011), .ZN(n10467) );
  INR4D1BWP30P140LVT U8847 ( .A1(i_cmd[189]), .B1(i_cmd[173]), .B2(n6013), 
        .B3(n9844), .ZN(n10466) );
  AOI22D1BWP30P140LVT U8848 ( .A1(i_data_bus[669]), .A2(n10467), .B1(
        i_data_bus[765]), .B2(n10466), .ZN(n6014) );
  ND2D1BWP30P140LVT U8849 ( .A1(n6015), .A2(n6014), .ZN(N11050) );
  AOI22D1BWP30P140LVT U8850 ( .A1(i_data_bus[372]), .A2(n10542), .B1(
        i_data_bus[308]), .B2(n10541), .ZN(n6017) );
  AOI22D1BWP30P140LVT U8851 ( .A1(i_data_bus[340]), .A2(n10544), .B1(
        i_data_bus[276]), .B2(n10543), .ZN(n6016) );
  ND2D1BWP30P140LVT U8852 ( .A1(n6017), .A2(n6016), .ZN(N6645) );
  AOI22D1BWP30P140LVT U8853 ( .A1(i_data_bus[728]), .A2(n10465), .B1(
        i_data_bus[696]), .B2(n10468), .ZN(n6019) );
  AOI22D1BWP30P140LVT U8854 ( .A1(i_data_bus[664]), .A2(n10467), .B1(
        i_data_bus[760]), .B2(n10466), .ZN(n6018) );
  ND2D1BWP30P140LVT U8855 ( .A1(n6019), .A2(n6018), .ZN(N11045) );
  AOI22D1BWP30P140LVT U8856 ( .A1(i_data_bus[348]), .A2(n10544), .B1(
        i_data_bus[316]), .B2(n10541), .ZN(n6021) );
  AOI22D1BWP30P140LVT U8857 ( .A1(i_data_bus[380]), .A2(n10542), .B1(
        i_data_bus[284]), .B2(n10543), .ZN(n6020) );
  ND2D1BWP30P140LVT U8858 ( .A1(n6021), .A2(n6020), .ZN(N6653) );
  AOI22D1BWP30P140LVT U8859 ( .A1(i_data_bus[713]), .A2(n10465), .B1(
        i_data_bus[681]), .B2(n10468), .ZN(n6023) );
  AOI22D1BWP30P140LVT U8860 ( .A1(i_data_bus[649]), .A2(n10467), .B1(
        i_data_bus[745]), .B2(n10466), .ZN(n6022) );
  ND2D1BWP30P140LVT U8861 ( .A1(n6023), .A2(n6022), .ZN(N11030) );
  AOI22D1BWP30P140LVT U8862 ( .A1(i_data_bus[352]), .A2(n10542), .B1(
        i_data_bus[288]), .B2(n10541), .ZN(n6025) );
  AOI22D1BWP30P140LVT U8863 ( .A1(i_data_bus[320]), .A2(n10544), .B1(
        i_data_bus[256]), .B2(n10543), .ZN(n6024) );
  ND2D1BWP30P140LVT U8864 ( .A1(n6025), .A2(n6024), .ZN(N6625) );
  AOI22D1BWP30P140LVT U8865 ( .A1(i_data_bus[642]), .A2(n10467), .B1(
        i_data_bus[674]), .B2(n10468), .ZN(n6027) );
  AOI22D1BWP30P140LVT U8866 ( .A1(i_data_bus[706]), .A2(n10465), .B1(
        i_data_bus[738]), .B2(n10466), .ZN(n6026) );
  ND2D1BWP30P140LVT U8867 ( .A1(n6027), .A2(n6026), .ZN(N11023) );
  AOI22D1BWP30P140LVT U8868 ( .A1(i_data_bus[279]), .A2(n10543), .B1(
        i_data_bus[311]), .B2(n10541), .ZN(n6029) );
  AOI22D1BWP30P140LVT U8869 ( .A1(i_data_bus[375]), .A2(n10542), .B1(
        i_data_bus[343]), .B2(n10544), .ZN(n6028) );
  ND2D1BWP30P140LVT U8870 ( .A1(n6029), .A2(n6028), .ZN(N6648) );
  AOI22D1BWP30P140LVT U8871 ( .A1(i_data_bus[269]), .A2(n10543), .B1(
        i_data_bus[301]), .B2(n10541), .ZN(n6031) );
  AOI22D1BWP30P140LVT U8872 ( .A1(i_data_bus[365]), .A2(n10542), .B1(
        i_data_bus[333]), .B2(n10544), .ZN(n6030) );
  ND2D1BWP30P140LVT U8873 ( .A1(n6031), .A2(n6030), .ZN(N6638) );
  AOI22D1BWP30P140LVT U8874 ( .A1(i_data_bus[716]), .A2(n10402), .B1(
        i_data_bus[684]), .B2(n10404), .ZN(n6033) );
  AOI22D1BWP30P140LVT U8875 ( .A1(i_data_bus[652]), .A2(n10401), .B1(
        i_data_bus[748]), .B2(n10403), .ZN(n6032) );
  ND2D1BWP30P140LVT U8876 ( .A1(n6033), .A2(n6032), .ZN(N14781) );
  AOI22D1BWP30P140LVT U8877 ( .A1(i_data_bus[710]), .A2(n10402), .B1(
        i_data_bus[678]), .B2(n10404), .ZN(n6035) );
  AOI22D1BWP30P140LVT U8878 ( .A1(i_data_bus[646]), .A2(n10401), .B1(
        i_data_bus[742]), .B2(n10403), .ZN(n6034) );
  ND2D1BWP30P140LVT U8879 ( .A1(n6035), .A2(n6034), .ZN(N14775) );
  AOI22D1BWP30P140LVT U8880 ( .A1(i_data_bus[493]), .A2(n10571), .B1(
        i_data_bus[461]), .B2(n10570), .ZN(n6037) );
  AOI22D1BWP30P140LVT U8881 ( .A1(i_data_bus[429]), .A2(n10569), .B1(
        i_data_bus[397]), .B2(n10572), .ZN(n6036) );
  ND2D1BWP30P140LVT U8882 ( .A1(n6037), .A2(n6036), .ZN(N4980) );
  AOI22D1BWP30P140LVT U8883 ( .A1(i_data_bus[444]), .A2(n10569), .B1(
        i_data_bus[476]), .B2(n10570), .ZN(n6039) );
  AOI22D1BWP30P140LVT U8884 ( .A1(i_data_bus[508]), .A2(n10571), .B1(
        i_data_bus[412]), .B2(n10572), .ZN(n6038) );
  ND2D1BWP30P140LVT U8885 ( .A1(n6039), .A2(n6038), .ZN(N4995) );
  AOI22D1BWP30P140LVT U8886 ( .A1(i_data_bus[645]), .A2(n10467), .B1(
        i_data_bus[741]), .B2(n10466), .ZN(n6041) );
  AOI22D1BWP30P140LVT U8887 ( .A1(i_data_bus[709]), .A2(n10465), .B1(
        i_data_bus[677]), .B2(n10468), .ZN(n6040) );
  ND2D1BWP30P140LVT U8888 ( .A1(n6041), .A2(n6040), .ZN(N11026) );
  AOI22D1BWP30P140LVT U8889 ( .A1(i_data_bus[722]), .A2(n10465), .B1(
        i_data_bus[754]), .B2(n10466), .ZN(n6043) );
  AOI22D1BWP30P140LVT U8890 ( .A1(i_data_bus[658]), .A2(n10467), .B1(
        i_data_bus[690]), .B2(n10468), .ZN(n6042) );
  ND2D1BWP30P140LVT U8891 ( .A1(n6043), .A2(n6042), .ZN(N11039) );
  AOI22D1BWP30P140LVT U8892 ( .A1(i_data_bus[710]), .A2(n10465), .B1(
        i_data_bus[742]), .B2(n10466), .ZN(n6045) );
  AOI22D1BWP30P140LVT U8893 ( .A1(i_data_bus[646]), .A2(n10467), .B1(
        i_data_bus[678]), .B2(n10468), .ZN(n6044) );
  ND2D1BWP30P140LVT U8894 ( .A1(n6045), .A2(n6044), .ZN(N11027) );
  AOI22D1BWP30P140LVT U8895 ( .A1(i_data_bus[566]), .A2(n10535), .B1(
        i_data_bus[534]), .B2(n10533), .ZN(n6047) );
  AOI22D1BWP30P140LVT U8896 ( .A1(i_data_bus[630]), .A2(n10534), .B1(
        i_data_bus[598]), .B2(n10536), .ZN(n6046) );
  ND2D1BWP30P140LVT U8897 ( .A1(n6047), .A2(n6046), .ZN(N7079) );
  AOI22D1BWP30P140LVT U8898 ( .A1(i_data_bus[628]), .A2(n10407), .B1(
        i_data_bus[532]), .B2(n10405), .ZN(n6049) );
  AOI22D1BWP30P140LVT U8899 ( .A1(i_data_bus[564]), .A2(n10406), .B1(
        i_data_bus[596]), .B2(n10408), .ZN(n6048) );
  ND2D1BWP30P140LVT U8900 ( .A1(n6049), .A2(n6048), .ZN(N14573) );
  AOI22D1BWP30P140LVT U8901 ( .A1(i_data_bus[618]), .A2(n10407), .B1(
        i_data_bus[522]), .B2(n10405), .ZN(n6051) );
  AOI22D1BWP30P140LVT U8902 ( .A1(i_data_bus[554]), .A2(n10406), .B1(
        i_data_bus[586]), .B2(n10408), .ZN(n6050) );
  ND2D1BWP30P140LVT U8903 ( .A1(n6051), .A2(n6050), .ZN(N14563) );
  AOI22D1BWP30P140LVT U8904 ( .A1(i_data_bus[550]), .A2(n10406), .B1(
        i_data_bus[518]), .B2(n10405), .ZN(n6053) );
  AOI22D1BWP30P140LVT U8905 ( .A1(i_data_bus[614]), .A2(n10407), .B1(
        i_data_bus[582]), .B2(n10408), .ZN(n6052) );
  ND2D1BWP30P140LVT U8906 ( .A1(n6053), .A2(n6052), .ZN(N14559) );
  AOI22D1BWP30P140LVT U8907 ( .A1(i_data_bus[608]), .A2(n10534), .B1(
        i_data_bus[512]), .B2(n10533), .ZN(n6055) );
  AOI22D1BWP30P140LVT U8908 ( .A1(i_data_bus[544]), .A2(n10535), .B1(
        i_data_bus[576]), .B2(n10536), .ZN(n6054) );
  ND2D1BWP30P140LVT U8909 ( .A1(n6055), .A2(n6054), .ZN(N7057) );
  AOI22D1BWP30P140LVT U8910 ( .A1(i_data_bus[560]), .A2(n10406), .B1(
        i_data_bus[528]), .B2(n10405), .ZN(n6057) );
  AOI22D1BWP30P140LVT U8911 ( .A1(i_data_bus[624]), .A2(n10407), .B1(
        i_data_bus[592]), .B2(n10408), .ZN(n6056) );
  ND2D1BWP30P140LVT U8912 ( .A1(n6057), .A2(n6056), .ZN(N14569) );
  AOI22D1BWP30P140LVT U8913 ( .A1(i_data_bus[557]), .A2(n10406), .B1(
        i_data_bus[525]), .B2(n10405), .ZN(n6059) );
  AOI22D1BWP30P140LVT U8914 ( .A1(i_data_bus[621]), .A2(n10407), .B1(
        i_data_bus[589]), .B2(n10408), .ZN(n6058) );
  ND2D1BWP30P140LVT U8915 ( .A1(n6059), .A2(n6058), .ZN(N14566) );
  AOI22D1BWP30P140LVT U8916 ( .A1(i_data_bus[638]), .A2(n10407), .B1(
        i_data_bus[542]), .B2(n10405), .ZN(n6061) );
  AOI22D1BWP30P140LVT U8917 ( .A1(i_data_bus[574]), .A2(n10406), .B1(
        i_data_bus[606]), .B2(n10408), .ZN(n6060) );
  ND2D1BWP30P140LVT U8918 ( .A1(n6061), .A2(n6060), .ZN(N14583) );
  AOI22D1BWP30P140LVT U8919 ( .A1(i_data_bus[638]), .A2(n10534), .B1(
        i_data_bus[542]), .B2(n10533), .ZN(n6063) );
  AOI22D1BWP30P140LVT U8920 ( .A1(i_data_bus[574]), .A2(n10535), .B1(
        i_data_bus[606]), .B2(n10536), .ZN(n6062) );
  ND2D1BWP30P140LVT U8921 ( .A1(n6063), .A2(n6062), .ZN(N7087) );
  AOI22D1BWP30P140LVT U8922 ( .A1(i_data_bus[625]), .A2(n10534), .B1(
        i_data_bus[529]), .B2(n10533), .ZN(n6065) );
  AOI22D1BWP30P140LVT U8923 ( .A1(i_data_bus[561]), .A2(n10535), .B1(
        i_data_bus[593]), .B2(n10536), .ZN(n6064) );
  ND2D1BWP30P140LVT U8924 ( .A1(n6065), .A2(n6064), .ZN(N7074) );
  AOI22D1BWP30P140LVT U8925 ( .A1(i_data_bus[628]), .A2(n10534), .B1(
        i_data_bus[532]), .B2(n10533), .ZN(n6067) );
  AOI22D1BWP30P140LVT U8926 ( .A1(i_data_bus[564]), .A2(n10535), .B1(
        i_data_bus[596]), .B2(n10536), .ZN(n6066) );
  ND2D1BWP30P140LVT U8927 ( .A1(n6067), .A2(n6066), .ZN(N7077) );
  AOI22D1BWP30P140LVT U8928 ( .A1(i_data_bus[614]), .A2(n10534), .B1(
        i_data_bus[518]), .B2(n10533), .ZN(n6069) );
  AOI22D1BWP30P140LVT U8929 ( .A1(i_data_bus[550]), .A2(n10535), .B1(
        i_data_bus[582]), .B2(n10536), .ZN(n6068) );
  ND2D1BWP30P140LVT U8930 ( .A1(n6069), .A2(n6068), .ZN(N7063) );
  AOI22D1BWP30P140LVT U8931 ( .A1(i_data_bus[621]), .A2(n10534), .B1(
        i_data_bus[525]), .B2(n10533), .ZN(n6071) );
  AOI22D1BWP30P140LVT U8932 ( .A1(i_data_bus[557]), .A2(n10535), .B1(
        i_data_bus[589]), .B2(n10536), .ZN(n6070) );
  ND2D1BWP30P140LVT U8933 ( .A1(n6071), .A2(n6070), .ZN(N7070) );
  AOI22D1BWP30P140LVT U8934 ( .A1(i_data_bus[353]), .A2(n10574), .B1(
        i_data_bus[289]), .B2(n10573), .ZN(n6073) );
  AOI22D1BWP30P140LVT U8935 ( .A1(i_data_bus[257]), .A2(n10575), .B1(
        i_data_bus[321]), .B2(n10576), .ZN(n6072) );
  ND2D1BWP30P140LVT U8936 ( .A1(n6073), .A2(n6072), .ZN(N4752) );
  AOI22D1BWP30P140LVT U8937 ( .A1(i_data_bus[352]), .A2(n10574), .B1(
        i_data_bus[288]), .B2(n10573), .ZN(n6075) );
  AOI22D1BWP30P140LVT U8938 ( .A1(i_data_bus[320]), .A2(n10576), .B1(
        i_data_bus[256]), .B2(n10575), .ZN(n6074) );
  ND2D1BWP30P140LVT U8939 ( .A1(n6075), .A2(n6074), .ZN(N4751) );
  AOI22D1BWP30P140LVT U8940 ( .A1(i_data_bus[357]), .A2(n10574), .B1(
        i_data_bus[293]), .B2(n10573), .ZN(n6077) );
  AOI22D1BWP30P140LVT U8941 ( .A1(i_data_bus[325]), .A2(n10576), .B1(
        i_data_bus[261]), .B2(n10575), .ZN(n6076) );
  ND2D1BWP30P140LVT U8942 ( .A1(n6077), .A2(n6076), .ZN(N4756) );
  AOI22D1BWP30P140LVT U8943 ( .A1(i_data_bus[269]), .A2(n10575), .B1(
        i_data_bus[301]), .B2(n10573), .ZN(n6079) );
  AOI22D1BWP30P140LVT U8944 ( .A1(i_data_bus[365]), .A2(n10574), .B1(
        i_data_bus[333]), .B2(n10576), .ZN(n6078) );
  ND2D1BWP30P140LVT U8945 ( .A1(n6079), .A2(n6078), .ZN(N4764) );
  AOI22D1BWP30P140LVT U8946 ( .A1(i_data_bus[284]), .A2(n10575), .B1(
        i_data_bus[316]), .B2(n10573), .ZN(n6081) );
  AOI22D1BWP30P140LVT U8947 ( .A1(i_data_bus[380]), .A2(n10574), .B1(
        i_data_bus[348]), .B2(n10576), .ZN(n6080) );
  ND2D1BWP30P140LVT U8948 ( .A1(n6081), .A2(n6080), .ZN(N4779) );
  AOI22D1BWP30P140LVT U8949 ( .A1(i_data_bus[363]), .A2(n10574), .B1(
        i_data_bus[299]), .B2(n10573), .ZN(n6083) );
  AOI22D1BWP30P140LVT U8950 ( .A1(i_data_bus[267]), .A2(n10575), .B1(
        i_data_bus[331]), .B2(n10576), .ZN(n6082) );
  ND2D1BWP30P140LVT U8951 ( .A1(n6083), .A2(n6082), .ZN(N4762) );
  AOI22D1BWP30P140LVT U8952 ( .A1(i_data_bus[132]), .A2(n10612), .B1(
        i_data_bus[164]), .B2(n10609), .ZN(n6085) );
  AOI22D1BWP30P140LVT U8953 ( .A1(i_data_bus[228]), .A2(n10611), .B1(
        i_data_bus[196]), .B2(n10610), .ZN(n6084) );
  ND2D1BWP30P140LVT U8954 ( .A1(n6085), .A2(n6084), .ZN(N2665) );
  AOI22D1BWP30P140LVT U8955 ( .A1(i_data_bus[436]), .A2(n10569), .B1(
        i_data_bus[500]), .B2(n10571), .ZN(n6087) );
  AOI22D1BWP30P140LVT U8956 ( .A1(i_data_bus[404]), .A2(n10572), .B1(
        i_data_bus[468]), .B2(n10570), .ZN(n6086) );
  ND2D1BWP30P140LVT U8957 ( .A1(n6087), .A2(n6086), .ZN(N4987) );
  AOI22D1BWP30P140LVT U8958 ( .A1(i_data_bus[233]), .A2(n10611), .B1(
        i_data_bus[169]), .B2(n10609), .ZN(n6089) );
  AOI22D1BWP30P140LVT U8959 ( .A1(i_data_bus[201]), .A2(n10610), .B1(
        i_data_bus[137]), .B2(n10612), .ZN(n6088) );
  ND2D1BWP30P140LVT U8960 ( .A1(n6089), .A2(n6088), .ZN(N2670) );
  AOI22D1BWP30P140LVT U8961 ( .A1(i_data_bus[230]), .A2(n10611), .B1(
        i_data_bus[166]), .B2(n10609), .ZN(n6091) );
  AOI22D1BWP30P140LVT U8962 ( .A1(i_data_bus[198]), .A2(n10610), .B1(
        i_data_bus[134]), .B2(n10612), .ZN(n6090) );
  ND2D1BWP30P140LVT U8963 ( .A1(n6091), .A2(n6090), .ZN(N2667) );
  AOI22D1BWP30P140LVT U8964 ( .A1(i_data_bus[174]), .A2(n10609), .B1(
        i_data_bus[206]), .B2(n10610), .ZN(n6093) );
  AOI22D1BWP30P140LVT U8965 ( .A1(i_data_bus[238]), .A2(n10611), .B1(
        i_data_bus[142]), .B2(n10612), .ZN(n6092) );
  ND2D1BWP30P140LVT U8966 ( .A1(n6093), .A2(n6092), .ZN(N2675) );
  AOI22D1BWP30P140LVT U8967 ( .A1(i_data_bus[249]), .A2(n10611), .B1(
        i_data_bus[185]), .B2(n10609), .ZN(n6095) );
  AOI22D1BWP30P140LVT U8968 ( .A1(i_data_bus[217]), .A2(n10610), .B1(
        i_data_bus[153]), .B2(n10612), .ZN(n6094) );
  ND2D1BWP30P140LVT U8969 ( .A1(n6095), .A2(n6094), .ZN(N2686) );
  AOI22D1BWP30P140LVT U8970 ( .A1(i_data_bus[253]), .A2(n10611), .B1(
        i_data_bus[221]), .B2(n10610), .ZN(n6097) );
  AOI22D1BWP30P140LVT U8971 ( .A1(i_data_bus[189]), .A2(n10609), .B1(
        i_data_bus[157]), .B2(n10612), .ZN(n6096) );
  ND2D1BWP30P140LVT U8972 ( .A1(n6097), .A2(n6096), .ZN(N2690) );
  AOI22D1BWP30P140LVT U8973 ( .A1(i_data_bus[954]), .A2(n10428), .B1(
        i_data_bus[922]), .B2(n10425), .ZN(n6099) );
  AOI22D1BWP30P140LVT U8974 ( .A1(i_data_bus[986]), .A2(n10426), .B1(
        i_data_bus[1018]), .B2(n10427), .ZN(n6098) );
  ND2D1BWP30P140LVT U8975 ( .A1(n6099), .A2(n6098), .ZN(N13353) );
  AOI22D1BWP30P140LVT U8976 ( .A1(i_data_bus[1008]), .A2(n10427), .B1(
        i_data_bus[912]), .B2(n10425), .ZN(n6101) );
  AOI22D1BWP30P140LVT U8977 ( .A1(i_data_bus[976]), .A2(n10426), .B1(
        i_data_bus[944]), .B2(n10428), .ZN(n6100) );
  ND2D1BWP30P140LVT U8978 ( .A1(n6101), .A2(n6100), .ZN(N13343) );
  AOI22D1BWP30P140LVT U8979 ( .A1(i_data_bus[997]), .A2(n10427), .B1(
        i_data_bus[901]), .B2(n10425), .ZN(n6103) );
  AOI22D1BWP30P140LVT U8980 ( .A1(i_data_bus[965]), .A2(n10426), .B1(
        i_data_bus[933]), .B2(n10428), .ZN(n6102) );
  ND2D1BWP30P140LVT U8981 ( .A1(n6103), .A2(n6102), .ZN(N13332) );
  AOI22D1BWP30P140LVT U8982 ( .A1(i_data_bus[973]), .A2(n10426), .B1(
        i_data_bus[909]), .B2(n10425), .ZN(n6105) );
  AOI22D1BWP30P140LVT U8983 ( .A1(i_data_bus[1005]), .A2(n10427), .B1(
        i_data_bus[941]), .B2(n10428), .ZN(n6104) );
  ND2D1BWP30P140LVT U8984 ( .A1(n6105), .A2(n6104), .ZN(N13340) );
  AOI22D1BWP30P140LVT U8985 ( .A1(i_data_bus[966]), .A2(n10426), .B1(
        i_data_bus[902]), .B2(n10425), .ZN(n6107) );
  AOI22D1BWP30P140LVT U8986 ( .A1(i_data_bus[934]), .A2(n10428), .B1(
        i_data_bus[998]), .B2(n10427), .ZN(n6106) );
  ND2D1BWP30P140LVT U8987 ( .A1(n6107), .A2(n6106), .ZN(N13333) );
  AOI22D1BWP30P140LVT U8988 ( .A1(i_data_bus[610]), .A2(n10534), .B1(
        i_data_bus[546]), .B2(n10535), .ZN(n6109) );
  AOI22D1BWP30P140LVT U8989 ( .A1(i_data_bus[578]), .A2(n10536), .B1(
        i_data_bus[514]), .B2(n10533), .ZN(n6108) );
  ND2D1BWP30P140LVT U8990 ( .A1(n6109), .A2(n6108), .ZN(N7059) );
  AOI22D1BWP30P140LVT U8991 ( .A1(i_data_bus[619]), .A2(n10534), .B1(
        i_data_bus[555]), .B2(n10535), .ZN(n6111) );
  AOI22D1BWP30P140LVT U8992 ( .A1(i_data_bus[587]), .A2(n10536), .B1(
        i_data_bus[523]), .B2(n10533), .ZN(n6110) );
  ND2D1BWP30P140LVT U8993 ( .A1(n6111), .A2(n6110), .ZN(N7068) );
  AOI22D1BWP30P140LVT U8994 ( .A1(i_data_bus[626]), .A2(n10534), .B1(
        i_data_bus[562]), .B2(n10535), .ZN(n6113) );
  AOI22D1BWP30P140LVT U8995 ( .A1(i_data_bus[594]), .A2(n10536), .B1(
        i_data_bus[530]), .B2(n10533), .ZN(n6112) );
  ND2D1BWP30P140LVT U8996 ( .A1(n6113), .A2(n6112), .ZN(N7075) );
  AOI22D1BWP30P140LVT U8997 ( .A1(i_data_bus[541]), .A2(n10533), .B1(
        i_data_bus[573]), .B2(n10535), .ZN(n6115) );
  AOI22D1BWP30P140LVT U8998 ( .A1(i_data_bus[637]), .A2(n10534), .B1(
        i_data_bus[605]), .B2(n10536), .ZN(n6114) );
  ND2D1BWP30P140LVT U8999 ( .A1(n6115), .A2(n6114), .ZN(N7086) );
  AOI22D1BWP30P140LVT U9000 ( .A1(i_data_bus[609]), .A2(n10534), .B1(
        i_data_bus[545]), .B2(n10535), .ZN(n6117) );
  AOI22D1BWP30P140LVT U9001 ( .A1(i_data_bus[513]), .A2(n10533), .B1(
        i_data_bus[577]), .B2(n10536), .ZN(n6116) );
  ND2D1BWP30P140LVT U9002 ( .A1(n6117), .A2(n6116), .ZN(N7058) );
  AOI22D1BWP30P140LVT U9003 ( .A1(i_data_bus[515]), .A2(n10533), .B1(
        i_data_bus[547]), .B2(n10535), .ZN(n6119) );
  AOI22D1BWP30P140LVT U9004 ( .A1(i_data_bus[611]), .A2(n10534), .B1(
        i_data_bus[579]), .B2(n10536), .ZN(n6118) );
  ND2D1BWP30P140LVT U9005 ( .A1(n6119), .A2(n6118), .ZN(N7060) );
  NR3D0P7BWP30P140LVT U9006 ( .A1(inner_first_stage_valid_reg[33]), .A2(
        inner_first_stage_valid_reg[34]), .A3(inner_first_stage_valid_reg[35]), 
        .ZN(n6125) );
  INR3D0BWP30P140LVT U9007 ( .A1(n6125), .B1(inner_first_stage_valid_reg[37]), 
        .B2(inner_first_stage_valid_reg[32]), .ZN(n6128) );
  INR3D2BWP30P140LVT U9008 ( .A1(inner_first_stage_valid_reg[39]), .B1(
        inner_first_stage_valid_reg[38]), .B2(n6123), .ZN(n11354) );
  NR2D1BWP30P140LVT U9009 ( .A1(inner_first_stage_valid_reg[37]), .A2(
        inner_first_stage_valid_reg[33]), .ZN(n6121) );
  INR3D2BWP30P140LVT U9010 ( .A1(inner_first_stage_valid_reg[34]), .B1(
        inner_first_stage_valid_reg[35]), .B2(n6122), .ZN(n11353) );
  INR3D2BWP30P140LVT U9011 ( .A1(inner_first_stage_valid_reg[35]), .B1(
        inner_first_stage_valid_reg[34]), .B2(n6122), .ZN(n11352) );
  INR3D2BWP30P140LVT U9012 ( .A1(inner_first_stage_valid_reg[38]), .B1(
        inner_first_stage_valid_reg[39]), .B2(n6123), .ZN(n11351) );
  NR4D0BWP30P140LVT U9013 ( .A1(n11354), .A2(n11353), .A3(n11352), .A4(n11351), 
        .ZN(n6132) );
  NR2D1BWP30P140LVT U9014 ( .A1(inner_first_stage_valid_reg[34]), .A2(
        inner_first_stage_valid_reg[35]), .ZN(n6126) );
  INR4D1BWP30P140LVT U9015 ( .A1(inner_first_stage_valid_reg[32]), .B1(
        inner_first_stage_valid_reg[37]), .B2(inner_first_stage_valid_reg[33]), 
        .B3(n6130), .ZN(n11350) );
  NR4D0BWP30P140LVT U9016 ( .A1(n11348), .A2(n11350), .A3(n11349), .A4(n11339), 
        .ZN(n6131) );
  ND2D1BWP30P140LVT U9017 ( .A1(n6132), .A2(n6131), .ZN(N9724) );
  AOI22D1BWP30P140LVT U9018 ( .A1(i_data_bus[732]), .A2(n10465), .B1(
        i_data_bus[668]), .B2(n10467), .ZN(n6134) );
  AOI22D1BWP30P140LVT U9019 ( .A1(i_data_bus[764]), .A2(n10466), .B1(
        i_data_bus[700]), .B2(n10468), .ZN(n6133) );
  ND2D1BWP30P140LVT U9020 ( .A1(n6134), .A2(n6133), .ZN(N11049) );
  AOI22D1BWP30P140LVT U9021 ( .A1(i_data_bus[702]), .A2(n10468), .B1(
        i_data_bus[670]), .B2(n10467), .ZN(n6136) );
  AOI22D1BWP30P140LVT U9022 ( .A1(i_data_bus[734]), .A2(n10465), .B1(
        i_data_bus[766]), .B2(n10466), .ZN(n6135) );
  ND2D1BWP30P140LVT U9023 ( .A1(n6136), .A2(n6135), .ZN(N11051) );
  AOI22D1BWP30P140LVT U9024 ( .A1(i_data_bus[715]), .A2(n10465), .B1(
        i_data_bus[651]), .B2(n10467), .ZN(n6138) );
  AOI22D1BWP30P140LVT U9025 ( .A1(i_data_bus[747]), .A2(n10466), .B1(
        i_data_bus[683]), .B2(n10468), .ZN(n6137) );
  ND2D1BWP30P140LVT U9026 ( .A1(n6138), .A2(n6137), .ZN(N11032) );
  AOI22D1BWP30P140LVT U9027 ( .A1(i_data_bus[686]), .A2(n10468), .B1(
        i_data_bus[654]), .B2(n10467), .ZN(n6140) );
  AOI22D1BWP30P140LVT U9028 ( .A1(i_data_bus[718]), .A2(n10465), .B1(
        i_data_bus[750]), .B2(n10466), .ZN(n6139) );
  ND2D1BWP30P140LVT U9029 ( .A1(n6140), .A2(n6139), .ZN(N11035) );
  AOI22D1BWP30P140LVT U9030 ( .A1(i_data_bus[725]), .A2(n10465), .B1(
        i_data_bus[661]), .B2(n10467), .ZN(n6142) );
  AOI22D1BWP30P140LVT U9031 ( .A1(i_data_bus[757]), .A2(n10466), .B1(
        i_data_bus[693]), .B2(n10468), .ZN(n6141) );
  ND2D1BWP30P140LVT U9032 ( .A1(n6142), .A2(n6141), .ZN(N11042) );
  AOI22D1BWP30P140LVT U9033 ( .A1(i_data_bus[716]), .A2(n10465), .B1(
        i_data_bus[652]), .B2(n10467), .ZN(n6144) );
  AOI22D1BWP30P140LVT U9034 ( .A1(i_data_bus[684]), .A2(n10468), .B1(
        i_data_bus[748]), .B2(n10466), .ZN(n6143) );
  ND2D1BWP30P140LVT U9035 ( .A1(n6144), .A2(n6143), .ZN(N11033) );
  AOI22D1BWP30P140LVT U9036 ( .A1(i_data_bus[626]), .A2(n10407), .B1(
        i_data_bus[562]), .B2(n10406), .ZN(n6146) );
  AOI22D1BWP30P140LVT U9037 ( .A1(i_data_bus[594]), .A2(n10408), .B1(
        i_data_bus[530]), .B2(n10405), .ZN(n6145) );
  ND2D1BWP30P140LVT U9038 ( .A1(n6146), .A2(n6145), .ZN(N14571) );
  AOI22D1BWP30P140LVT U9039 ( .A1(i_data_bus[629]), .A2(n10407), .B1(
        i_data_bus[565]), .B2(n10406), .ZN(n6148) );
  AOI22D1BWP30P140LVT U9040 ( .A1(i_data_bus[597]), .A2(n10408), .B1(
        i_data_bus[533]), .B2(n10405), .ZN(n6147) );
  ND2D1BWP30P140LVT U9041 ( .A1(n6148), .A2(n6147), .ZN(N14574) );
  AOI22D1BWP30P140LVT U9042 ( .A1(i_data_bus[578]), .A2(n10408), .B1(
        i_data_bus[546]), .B2(n10406), .ZN(n6150) );
  AOI22D1BWP30P140LVT U9043 ( .A1(i_data_bus[610]), .A2(n10407), .B1(
        i_data_bus[514]), .B2(n10405), .ZN(n6149) );
  ND2D1BWP30P140LVT U9044 ( .A1(n6150), .A2(n6149), .ZN(N14555) );
  AOI22D1BWP30P140LVT U9045 ( .A1(i_data_bus[602]), .A2(n10408), .B1(
        i_data_bus[570]), .B2(n10406), .ZN(n6152) );
  AOI22D1BWP30P140LVT U9046 ( .A1(i_data_bus[634]), .A2(n10407), .B1(
        i_data_bus[538]), .B2(n10405), .ZN(n6151) );
  ND2D1BWP30P140LVT U9047 ( .A1(n6152), .A2(n6151), .ZN(N14579) );
  AOI22D1BWP30P140LVT U9048 ( .A1(i_data_bus[515]), .A2(n10405), .B1(
        i_data_bus[547]), .B2(n10406), .ZN(n6154) );
  AOI22D1BWP30P140LVT U9049 ( .A1(i_data_bus[611]), .A2(n10407), .B1(
        i_data_bus[579]), .B2(n10408), .ZN(n6153) );
  ND2D1BWP30P140LVT U9050 ( .A1(n6154), .A2(n6153), .ZN(N14556) );
  AOI22D1BWP30P140LVT U9051 ( .A1(i_data_bus[627]), .A2(n10407), .B1(
        i_data_bus[563]), .B2(n10406), .ZN(n6156) );
  AOI22D1BWP30P140LVT U9052 ( .A1(i_data_bus[531]), .A2(n10405), .B1(
        i_data_bus[595]), .B2(n10408), .ZN(n6155) );
  ND2D1BWP30P140LVT U9053 ( .A1(n6156), .A2(n6155), .ZN(N14572) );
  AOI22D1BWP30P140LVT U9054 ( .A1(i_data_bus[512]), .A2(n10405), .B1(
        i_data_bus[544]), .B2(n10406), .ZN(n6158) );
  AOI22D1BWP30P140LVT U9055 ( .A1(i_data_bus[608]), .A2(n10407), .B1(
        i_data_bus[576]), .B2(n10408), .ZN(n6157) );
  ND2D1BWP30P140LVT U9056 ( .A1(n6158), .A2(n6157), .ZN(N14553) );
  AOI22D1BWP30P140LVT U9057 ( .A1(i_data_bus[979]), .A2(n10459), .B1(
        i_data_bus[915]), .B2(n10458), .ZN(n6160) );
  AOI22D1BWP30P140LVT U9058 ( .A1(i_data_bus[947]), .A2(n10460), .B1(
        i_data_bus[1011]), .B2(n10457), .ZN(n6159) );
  ND2D1BWP30P140LVT U9059 ( .A1(n6160), .A2(n6159), .ZN(N11472) );
  AOI22D1BWP30P140LVT U9060 ( .A1(i_data_bus[933]), .A2(n10460), .B1(
        i_data_bus[901]), .B2(n10458), .ZN(n6162) );
  AOI22D1BWP30P140LVT U9061 ( .A1(i_data_bus[965]), .A2(n10459), .B1(
        i_data_bus[997]), .B2(n10457), .ZN(n6161) );
  ND2D1BWP30P140LVT U9062 ( .A1(n6162), .A2(n6161), .ZN(N11458) );
  AOI22D1BWP30P140LVT U9063 ( .A1(i_data_bus[988]), .A2(n10459), .B1(
        i_data_bus[924]), .B2(n10458), .ZN(n6164) );
  AOI22D1BWP30P140LVT U9064 ( .A1(i_data_bus[1020]), .A2(n10457), .B1(
        i_data_bus[956]), .B2(n10460), .ZN(n6163) );
  ND2D1BWP30P140LVT U9065 ( .A1(n6164), .A2(n6163), .ZN(N11481) );
  AOI22D1BWP30P140LVT U9066 ( .A1(i_data_bus[1001]), .A2(n10457), .B1(
        i_data_bus[905]), .B2(n10458), .ZN(n6166) );
  AOI22D1BWP30P140LVT U9067 ( .A1(i_data_bus[969]), .A2(n10459), .B1(
        i_data_bus[937]), .B2(n10460), .ZN(n6165) );
  ND2D1BWP30P140LVT U9068 ( .A1(n6166), .A2(n6165), .ZN(N11462) );
  NR4D1BWP30P140LVT U9069 ( .A1(i_cmd[115]), .A2(n6169), .A3(n9758), .A4(n6167), .ZN(n10537) );
  NR4D1BWP30P140LVT U9070 ( .A1(i_cmd[99]), .A2(n9761), .A3(n6168), .A4(n6167), 
        .ZN(n10538) );
  AOI22D1BWP30P140LVT U9071 ( .A1(i_data_bus[384]), .A2(n10537), .B1(
        i_data_bus[448]), .B2(n10538), .ZN(n6172) );
  INR4D1BWP30P140LVT U9072 ( .A1(i_cmd[107]), .B1(i_cmd[123]), .B2(n9760), 
        .B3(n6170), .ZN(n10540) );
  INR4D1BWP30P140LVT U9073 ( .A1(i_cmd[123]), .B1(i_cmd[107]), .B2(n9764), 
        .B3(n6170), .ZN(n10539) );
  AOI22D1BWP30P140LVT U9074 ( .A1(i_data_bus[416]), .A2(n10540), .B1(
        i_data_bus[480]), .B2(n10539), .ZN(n6171) );
  ND2D1BWP30P140LVT U9075 ( .A1(n6172), .A2(n6171), .ZN(N6841) );
  AOI22D1BWP30P140LVT U9076 ( .A1(i_data_bus[408]), .A2(n10537), .B1(
        i_data_bus[472]), .B2(n10538), .ZN(n6174) );
  AOI22D1BWP30P140LVT U9077 ( .A1(i_data_bus[440]), .A2(n10540), .B1(
        i_data_bus[504]), .B2(n10539), .ZN(n6173) );
  ND2D1BWP30P140LVT U9078 ( .A1(n6174), .A2(n6173), .ZN(N6865) );
  AOI22D1BWP30P140LVT U9079 ( .A1(i_data_bus[397]), .A2(n10537), .B1(
        i_data_bus[461]), .B2(n10538), .ZN(n6176) );
  AOI22D1BWP30P140LVT U9080 ( .A1(i_data_bus[429]), .A2(n10540), .B1(
        i_data_bus[493]), .B2(n10539), .ZN(n6175) );
  ND2D1BWP30P140LVT U9081 ( .A1(n6176), .A2(n6175), .ZN(N6854) );
  AOI22D1BWP30P140LVT U9082 ( .A1(i_data_bus[404]), .A2(n10537), .B1(
        i_data_bus[468]), .B2(n10538), .ZN(n6178) );
  AOI22D1BWP30P140LVT U9083 ( .A1(i_data_bus[436]), .A2(n10540), .B1(
        i_data_bus[500]), .B2(n10539), .ZN(n6177) );
  ND2D1BWP30P140LVT U9084 ( .A1(n6178), .A2(n6177), .ZN(N6861) );
  AOI22D1BWP30P140LVT U9085 ( .A1(i_data_bus[455]), .A2(n10570), .B1(
        i_data_bus[423]), .B2(n10569), .ZN(n6180) );
  AOI22D1BWP30P140LVT U9086 ( .A1(i_data_bus[487]), .A2(n10571), .B1(
        i_data_bus[391]), .B2(n10572), .ZN(n6179) );
  ND2D1BWP30P140LVT U9087 ( .A1(n6180), .A2(n6179), .ZN(N4974) );
  AOI22D1BWP30P140LVT U9088 ( .A1(i_data_bus[482]), .A2(n10571), .B1(
        i_data_bus[418]), .B2(n10569), .ZN(n6182) );
  AOI22D1BWP30P140LVT U9089 ( .A1(i_data_bus[450]), .A2(n10570), .B1(
        i_data_bus[386]), .B2(n10572), .ZN(n6181) );
  ND2D1BWP30P140LVT U9090 ( .A1(n6182), .A2(n6181), .ZN(N4969) );
  AOI22D1BWP30P140LVT U9091 ( .A1(i_data_bus[410]), .A2(n10572), .B1(
        i_data_bus[442]), .B2(n10569), .ZN(n6184) );
  AOI22D1BWP30P140LVT U9092 ( .A1(i_data_bus[506]), .A2(n10571), .B1(
        i_data_bus[474]), .B2(n10570), .ZN(n6183) );
  ND2D1BWP30P140LVT U9093 ( .A1(n6184), .A2(n6183), .ZN(N4993) );
  AOI22D1BWP30P140LVT U9094 ( .A1(i_data_bus[704]), .A2(n10402), .B1(
        i_data_bus[640]), .B2(n10401), .ZN(n6186) );
  AOI22D1BWP30P140LVT U9095 ( .A1(i_data_bus[672]), .A2(n10404), .B1(
        i_data_bus[736]), .B2(n10403), .ZN(n6185) );
  ND2D1BWP30P140LVT U9096 ( .A1(n6186), .A2(n6185), .ZN(N14769) );
  AOI22D1BWP30P140LVT U9097 ( .A1(i_data_bus[740]), .A2(n10403), .B1(
        i_data_bus[644]), .B2(n10401), .ZN(n6188) );
  AOI22D1BWP30P140LVT U9098 ( .A1(i_data_bus[708]), .A2(n10402), .B1(
        i_data_bus[676]), .B2(n10404), .ZN(n6187) );
  ND2D1BWP30P140LVT U9099 ( .A1(n6188), .A2(n6187), .ZN(N14773) );
  AOI22D1BWP30P140LVT U9100 ( .A1(i_data_bus[711]), .A2(n10402), .B1(
        i_data_bus[647]), .B2(n10401), .ZN(n6190) );
  AOI22D1BWP30P140LVT U9101 ( .A1(i_data_bus[679]), .A2(n10404), .B1(
        i_data_bus[743]), .B2(n10403), .ZN(n6189) );
  ND2D1BWP30P140LVT U9102 ( .A1(n6190), .A2(n6189), .ZN(N14776) );
  AOI22D1BWP30P140LVT U9103 ( .A1(i_data_bus[702]), .A2(n10404), .B1(
        i_data_bus[670]), .B2(n10401), .ZN(n6192) );
  AOI22D1BWP30P140LVT U9104 ( .A1(i_data_bus[734]), .A2(n10402), .B1(
        i_data_bus[766]), .B2(n10403), .ZN(n6191) );
  ND2D1BWP30P140LVT U9105 ( .A1(n6192), .A2(n6191), .ZN(N14799) );
  AOI22D1BWP30P140LVT U9106 ( .A1(i_data_bus[696]), .A2(n10404), .B1(
        i_data_bus[664]), .B2(n10401), .ZN(n6194) );
  AOI22D1BWP30P140LVT U9107 ( .A1(i_data_bus[728]), .A2(n10402), .B1(
        i_data_bus[760]), .B2(n10403), .ZN(n6193) );
  ND2D1BWP30P140LVT U9108 ( .A1(n6194), .A2(n6193), .ZN(N14793) );
  AOI22D1BWP30P140LVT U9109 ( .A1(i_data_bus[751]), .A2(n10403), .B1(
        i_data_bus[655]), .B2(n10401), .ZN(n6196) );
  AOI22D1BWP30P140LVT U9110 ( .A1(i_data_bus[719]), .A2(n10402), .B1(
        i_data_bus[687]), .B2(n10404), .ZN(n6195) );
  ND2D1BWP30P140LVT U9111 ( .A1(n6196), .A2(n6195), .ZN(N14784) );
  AOI22D1BWP30P140LVT U9112 ( .A1(i_data_bus[713]), .A2(n10402), .B1(
        i_data_bus[649]), .B2(n10401), .ZN(n6198) );
  AOI22D1BWP30P140LVT U9113 ( .A1(i_data_bus[681]), .A2(n10404), .B1(
        i_data_bus[745]), .B2(n10403), .ZN(n6197) );
  ND2D1BWP30P140LVT U9114 ( .A1(n6198), .A2(n6197), .ZN(N14778) );
  AOI22D1BWP30P140LVT U9115 ( .A1(i_data_bus[709]), .A2(n10402), .B1(
        i_data_bus[645]), .B2(n10401), .ZN(n6200) );
  AOI22D1BWP30P140LVT U9116 ( .A1(i_data_bus[677]), .A2(n10404), .B1(
        i_data_bus[741]), .B2(n10403), .ZN(n6199) );
  ND2D1BWP30P140LVT U9117 ( .A1(n6200), .A2(n6199), .ZN(N14774) );
  AOI22D1BWP30P140LVT U9118 ( .A1(i_data_bus[752]), .A2(n10403), .B1(
        i_data_bus[656]), .B2(n10401), .ZN(n6202) );
  AOI22D1BWP30P140LVT U9119 ( .A1(i_data_bus[720]), .A2(n10402), .B1(
        i_data_bus[688]), .B2(n10404), .ZN(n6201) );
  ND2D1BWP30P140LVT U9120 ( .A1(n6202), .A2(n6201), .ZN(N14785) );
  AOI22D1BWP30P140LVT U9121 ( .A1(i_data_bus[700]), .A2(n10404), .B1(
        i_data_bus[668]), .B2(n10401), .ZN(n6204) );
  AOI22D1BWP30P140LVT U9122 ( .A1(i_data_bus[732]), .A2(n10402), .B1(
        i_data_bus[764]), .B2(n10403), .ZN(n6203) );
  ND2D1BWP30P140LVT U9123 ( .A1(n6204), .A2(n6203), .ZN(N14797) );
  AOI22D1BWP30P140LVT U9124 ( .A1(i_data_bus[370]), .A2(n10542), .B1(
        i_data_bus[274]), .B2(n10543), .ZN(n6206) );
  AOI22D1BWP30P140LVT U9125 ( .A1(i_data_bus[338]), .A2(n10544), .B1(
        i_data_bus[306]), .B2(n10541), .ZN(n6205) );
  ND2D1BWP30P140LVT U9126 ( .A1(n6206), .A2(n6205), .ZN(N6643) );
  AOI22D1BWP30P140LVT U9127 ( .A1(i_data_bus[262]), .A2(n10543), .B1(
        i_data_bus[326]), .B2(n10544), .ZN(n6208) );
  AOI22D1BWP30P140LVT U9128 ( .A1(i_data_bus[358]), .A2(n10542), .B1(
        i_data_bus[294]), .B2(n10541), .ZN(n6207) );
  ND2D1BWP30P140LVT U9129 ( .A1(n6208), .A2(n6207), .ZN(N6631) );
  AOI22D1BWP30P140LVT U9130 ( .A1(i_data_bus[382]), .A2(n10542), .B1(
        i_data_bus[350]), .B2(n10544), .ZN(n6210) );
  AOI22D1BWP30P140LVT U9131 ( .A1(i_data_bus[286]), .A2(n10543), .B1(
        i_data_bus[318]), .B2(n10541), .ZN(n6209) );
  ND2D1BWP30P140LVT U9132 ( .A1(n6210), .A2(n6209), .ZN(N6655) );
  AOI22D1BWP30P140LVT U9133 ( .A1(i_data_bus[364]), .A2(n10542), .B1(
        i_data_bus[268]), .B2(n10543), .ZN(n6212) );
  AOI22D1BWP30P140LVT U9134 ( .A1(i_data_bus[332]), .A2(n10544), .B1(
        i_data_bus[300]), .B2(n10541), .ZN(n6211) );
  ND2D1BWP30P140LVT U9135 ( .A1(n6212), .A2(n6211), .ZN(N6637) );
  AOI22D1BWP30P140LVT U9136 ( .A1(i_data_bus[336]), .A2(n10544), .B1(
        i_data_bus[272]), .B2(n10543), .ZN(n6214) );
  AOI22D1BWP30P140LVT U9137 ( .A1(i_data_bus[368]), .A2(n10542), .B1(
        i_data_bus[304]), .B2(n10541), .ZN(n6213) );
  ND2D1BWP30P140LVT U9138 ( .A1(n6214), .A2(n6213), .ZN(N6641) );
  AOI22D1BWP30P140LVT U9139 ( .A1(i_data_bus[280]), .A2(n10543), .B1(
        i_data_bus[344]), .B2(n10544), .ZN(n6216) );
  AOI22D1BWP30P140LVT U9140 ( .A1(i_data_bus[376]), .A2(n10542), .B1(
        i_data_bus[312]), .B2(n10541), .ZN(n6215) );
  ND2D1BWP30P140LVT U9141 ( .A1(n6216), .A2(n6215), .ZN(N6649) );
  NR4D1BWP30P140LVT U9142 ( .A1(i_cmd[212]), .A2(n6219), .A3(n9744), .A4(n6217), .ZN(n10493) );
  NR4D1BWP30P140LVT U9143 ( .A1(i_cmd[196]), .A2(n9741), .A3(n6218), .A4(n6217), .ZN(n10495) );
  AOI22D1BWP30P140LVT U9144 ( .A1(i_data_bus[780]), .A2(n10493), .B1(
        i_data_bus[844]), .B2(n10495), .ZN(n6222) );
  INR4D1BWP30P140LVT U9145 ( .A1(i_cmd[204]), .B1(i_cmd[220]), .B2(n9743), 
        .B3(n6220), .ZN(n10496) );
  INR4D1BWP30P140LVT U9146 ( .A1(i_cmd[220]), .B1(i_cmd[204]), .B2(n9747), 
        .B3(n6220), .ZN(n10494) );
  AOI22D1BWP30P140LVT U9147 ( .A1(i_data_bus[812]), .A2(n10496), .B1(
        i_data_bus[876]), .B2(n10494), .ZN(n6221) );
  ND2D1BWP30P140LVT U9148 ( .A1(n6222), .A2(n6221), .ZN(N9375) );
  AOI22D1BWP30P140LVT U9149 ( .A1(i_data_bus[813]), .A2(n10496), .B1(
        i_data_bus[845]), .B2(n10495), .ZN(n6224) );
  AOI22D1BWP30P140LVT U9150 ( .A1(i_data_bus[781]), .A2(n10493), .B1(
        i_data_bus[877]), .B2(n10494), .ZN(n6223) );
  ND2D1BWP30P140LVT U9151 ( .A1(n6224), .A2(n6223), .ZN(N9376) );
  INR4D1BWP30P140LVT U9152 ( .A1(i_cmd[206]), .B1(i_cmd[222]), .B2(n9743), 
        .B3(n6228), .ZN(n10430) );
  NR4D1BWP30P140LVT U9153 ( .A1(i_cmd[214]), .A2(n9744), .A3(n6225), .A4(n6226), .ZN(n10429) );
  AOI22D1BWP30P140LVT U9154 ( .A1(i_data_bus[825]), .A2(n10430), .B1(
        i_data_bus[793]), .B2(n10429), .ZN(n6230) );
  NR4D1BWP30P140LVT U9155 ( .A1(i_cmd[198]), .A2(n6227), .A3(n9741), .A4(n6226), .ZN(n10432) );
  INR4D1BWP30P140LVT U9156 ( .A1(i_cmd[222]), .B1(i_cmd[206]), .B2(n9747), 
        .B3(n6228), .ZN(n10431) );
  AOI22D1BWP30P140LVT U9157 ( .A1(i_data_bus[857]), .A2(n10432), .B1(
        i_data_bus[889]), .B2(n10431), .ZN(n6229) );
  ND2D1BWP30P140LVT U9158 ( .A1(n6230), .A2(n6229), .ZN(N13136) );
  AOI22D1BWP30P140LVT U9159 ( .A1(i_data_bus[813]), .A2(n10430), .B1(
        i_data_bus[781]), .B2(n10429), .ZN(n6232) );
  AOI22D1BWP30P140LVT U9160 ( .A1(i_data_bus[845]), .A2(n10432), .B1(
        i_data_bus[877]), .B2(n10431), .ZN(n6231) );
  ND2D1BWP30P140LVT U9161 ( .A1(n6232), .A2(n6231), .ZN(N13124) );
  AOI22D1BWP30P140LVT U9162 ( .A1(i_data_bus[800]), .A2(n10430), .B1(
        i_data_bus[768]), .B2(n10429), .ZN(n6234) );
  AOI22D1BWP30P140LVT U9163 ( .A1(i_data_bus[832]), .A2(n10432), .B1(
        i_data_bus[864]), .B2(n10431), .ZN(n6233) );
  ND2D1BWP30P140LVT U9164 ( .A1(n6234), .A2(n6233), .ZN(N13111) );
  NR4D1BWP30P140LVT U9165 ( .A1(i_cmd[199]), .A2(n6237), .A3(n9741), .A4(n6235), .ZN(n10399) );
  NR4D1BWP30P140LVT U9166 ( .A1(i_cmd[215]), .A2(n9744), .A3(n6236), .A4(n6235), .ZN(n10397) );
  AOI22D1BWP30P140LVT U9167 ( .A1(i_data_bus[843]), .A2(n10399), .B1(
        i_data_bus[779]), .B2(n10397), .ZN(n6240) );
  INR4D1BWP30P140LVT U9168 ( .A1(i_cmd[207]), .B1(i_cmd[223]), .B2(n9743), 
        .B3(n6238), .ZN(n10400) );
  INR4D1BWP30P140LVT U9169 ( .A1(i_cmd[223]), .B1(i_cmd[207]), .B2(n9747), 
        .B3(n6238), .ZN(n10398) );
  AOI22D1BWP30P140LVT U9170 ( .A1(i_data_bus[811]), .A2(n10400), .B1(
        i_data_bus[875]), .B2(n10398), .ZN(n6239) );
  ND2D1BWP30P140LVT U9171 ( .A1(n6240), .A2(n6239), .ZN(N14996) );
  INR4D1BWP30P140LVT U9172 ( .A1(i_cmd[116]), .B1(i_cmd[100]), .B2(n9761), 
        .B3(n6242), .ZN(n10508) );
  NR4D1BWP30P140LVT U9173 ( .A1(i_cmd[124]), .A2(n9760), .A3(n6241), .A4(n6243), .ZN(n10507) );
  AOI22D1BWP30P140LVT U9174 ( .A1(i_data_bus[473]), .A2(n10508), .B1(
        i_data_bus[441]), .B2(n10507), .ZN(n6246) );
  INR4D1BWP30P140LVT U9175 ( .A1(i_cmd[100]), .B1(i_cmd[116]), .B2(n9758), 
        .B3(n6242), .ZN(n10505) );
  NR4D1BWP30P140LVT U9176 ( .A1(i_cmd[108]), .A2(n6244), .A3(n9764), .A4(n6243), .ZN(n10506) );
  AOI22D1BWP30P140LVT U9177 ( .A1(i_data_bus[409]), .A2(n10505), .B1(
        i_data_bus[505]), .B2(n10506), .ZN(n6245) );
  ND2D1BWP30P140LVT U9178 ( .A1(n6246), .A2(n6245), .ZN(N8740) );
  NR4D1BWP30P140LVT U9179 ( .A1(i_cmd[118]), .A2(n6249), .A3(n9758), .A4(n6247), .ZN(n10441) );
  NR4D1BWP30P140LVT U9180 ( .A1(i_cmd[102]), .A2(n9761), .A3(n6248), .A4(n6247), .ZN(n10442) );
  AOI22D1BWP30P140LVT U9181 ( .A1(i_data_bus[398]), .A2(n10441), .B1(
        i_data_bus[462]), .B2(n10442), .ZN(n6252) );
  INR4D1BWP30P140LVT U9182 ( .A1(i_cmd[110]), .B1(i_cmd[126]), .B2(n9760), 
        .B3(n6250), .ZN(n10443) );
  INR4D1BWP30P140LVT U9183 ( .A1(i_cmd[126]), .B1(i_cmd[110]), .B2(n9764), 
        .B3(n6250), .ZN(n10444) );
  AOI22D1BWP30P140LVT U9184 ( .A1(i_data_bus[430]), .A2(n10443), .B1(
        i_data_bus[494]), .B2(n10444), .ZN(n6251) );
  ND2D1BWP30P140LVT U9185 ( .A1(n6252), .A2(n6251), .ZN(N12477) );
  AOI22D1BWP30P140LVT U9186 ( .A1(i_data_bus[360]), .A2(n10574), .B1(
        i_data_bus[264]), .B2(n10575), .ZN(n6254) );
  AOI22D1BWP30P140LVT U9187 ( .A1(i_data_bus[328]), .A2(n10576), .B1(
        i_data_bus[296]), .B2(n10573), .ZN(n6253) );
  ND2D1BWP30P140LVT U9188 ( .A1(n6254), .A2(n6253), .ZN(N4759) );
  AOI22D1BWP30P140LVT U9189 ( .A1(i_data_bus[385]), .A2(n10441), .B1(
        i_data_bus[449]), .B2(n10442), .ZN(n6256) );
  AOI22D1BWP30P140LVT U9190 ( .A1(i_data_bus[417]), .A2(n10443), .B1(
        i_data_bus[481]), .B2(n10444), .ZN(n6255) );
  ND2D1BWP30P140LVT U9191 ( .A1(n6256), .A2(n6255), .ZN(N12464) );
  AOI22D1BWP30P140LVT U9192 ( .A1(i_data_bus[270]), .A2(n10575), .B1(
        i_data_bus[334]), .B2(n10576), .ZN(n6258) );
  AOI22D1BWP30P140LVT U9193 ( .A1(i_data_bus[366]), .A2(n10574), .B1(
        i_data_bus[302]), .B2(n10573), .ZN(n6257) );
  ND2D1BWP30P140LVT U9194 ( .A1(n6258), .A2(n6257), .ZN(N4765) );
  AOI22D1BWP30P140LVT U9195 ( .A1(i_data_bus[371]), .A2(n10574), .B1(
        i_data_bus[339]), .B2(n10576), .ZN(n6260) );
  AOI22D1BWP30P140LVT U9196 ( .A1(i_data_bus[275]), .A2(n10575), .B1(
        i_data_bus[307]), .B2(n10573), .ZN(n6259) );
  ND2D1BWP30P140LVT U9197 ( .A1(n6260), .A2(n6259), .ZN(N4770) );
  AOI22D1BWP30P140LVT U9198 ( .A1(i_data_bus[368]), .A2(n10574), .B1(
        i_data_bus[272]), .B2(n10575), .ZN(n6262) );
  AOI22D1BWP30P140LVT U9199 ( .A1(i_data_bus[336]), .A2(n10576), .B1(
        i_data_bus[304]), .B2(n10573), .ZN(n6261) );
  ND2D1BWP30P140LVT U9200 ( .A1(n6262), .A2(n6261), .ZN(N4767) );
  AOI22D1BWP30P140LVT U9201 ( .A1(i_data_bus[364]), .A2(n10574), .B1(
        i_data_bus[268]), .B2(n10575), .ZN(n6264) );
  AOI22D1BWP30P140LVT U9202 ( .A1(i_data_bus[332]), .A2(n10576), .B1(
        i_data_bus[300]), .B2(n10573), .ZN(n6263) );
  ND2D1BWP30P140LVT U9203 ( .A1(n6264), .A2(n6263), .ZN(N4763) );
  AOI22D1BWP30P140LVT U9204 ( .A1(i_data_bus[350]), .A2(n10576), .B1(
        i_data_bus[286]), .B2(n10575), .ZN(n6266) );
  AOI22D1BWP30P140LVT U9205 ( .A1(i_data_bus[382]), .A2(n10574), .B1(
        i_data_bus[318]), .B2(n10573), .ZN(n6265) );
  ND2D1BWP30P140LVT U9206 ( .A1(n6266), .A2(n6265), .ZN(N4781) );
  AOI22D1BWP30P140LVT U9207 ( .A1(i_data_bus[280]), .A2(n10575), .B1(
        i_data_bus[344]), .B2(n10576), .ZN(n6268) );
  AOI22D1BWP30P140LVT U9208 ( .A1(i_data_bus[376]), .A2(n10574), .B1(
        i_data_bus[312]), .B2(n10573), .ZN(n6267) );
  ND2D1BWP30P140LVT U9209 ( .A1(n6268), .A2(n6267), .ZN(N4775) );
  AOI22D1BWP30P140LVT U9210 ( .A1(i_data_bus[395]), .A2(n10441), .B1(
        i_data_bus[459]), .B2(n10442), .ZN(n6270) );
  AOI22D1BWP30P140LVT U9211 ( .A1(i_data_bus[427]), .A2(n10443), .B1(
        i_data_bus[491]), .B2(n10444), .ZN(n6269) );
  ND2D1BWP30P140LVT U9212 ( .A1(n6270), .A2(n6269), .ZN(N12474) );
  AOI22D1BWP30P140LVT U9213 ( .A1(i_data_bus[384]), .A2(n10441), .B1(
        i_data_bus[448]), .B2(n10442), .ZN(n6272) );
  AOI22D1BWP30P140LVT U9214 ( .A1(i_data_bus[416]), .A2(n10443), .B1(
        i_data_bus[480]), .B2(n10444), .ZN(n6271) );
  ND2D1BWP30P140LVT U9215 ( .A1(n6272), .A2(n6271), .ZN(N12463) );
  AOI22D1BWP30P140LVT U9216 ( .A1(i_data_bus[388]), .A2(n10441), .B1(
        i_data_bus[452]), .B2(n10442), .ZN(n6274) );
  AOI22D1BWP30P140LVT U9217 ( .A1(i_data_bus[420]), .A2(n10443), .B1(
        i_data_bus[484]), .B2(n10444), .ZN(n6273) );
  ND2D1BWP30P140LVT U9218 ( .A1(n6274), .A2(n6273), .ZN(N12467) );
  INR4D1BWP30P140LVT U9219 ( .A1(i_cmd[71]), .B1(i_cmd[87]), .B2(n9808), .B3(
        n6275), .ZN(n10415) );
  INR4D1BWP30P140LVT U9220 ( .A1(i_cmd[87]), .B1(i_cmd[71]), .B2(n9807), .B3(
        n6275), .ZN(n10413) );
  AOI22D1BWP30P140LVT U9221 ( .A1(i_data_bus[280]), .A2(n10415), .B1(
        i_data_bus[344]), .B2(n10413), .ZN(n6280) );
  NR4D1BWP30P140LVT U9222 ( .A1(i_cmd[79]), .A2(n6276), .A3(n9812), .A4(n6277), 
        .ZN(n10416) );
  NR4D1BWP30P140LVT U9223 ( .A1(i_cmd[95]), .A2(n9813), .A3(n6278), .A4(n6277), 
        .ZN(n10414) );
  AOI22D1BWP30P140LVT U9224 ( .A1(i_data_bus[376]), .A2(n10416), .B1(
        i_data_bus[312]), .B2(n10414), .ZN(n6279) );
  ND2D1BWP30P140LVT U9225 ( .A1(n6280), .A2(n6279), .ZN(N14145) );
  AOI22D1BWP30P140LVT U9226 ( .A1(i_data_bus[364]), .A2(n10416), .B1(
        i_data_bus[332]), .B2(n10413), .ZN(n6282) );
  AOI22D1BWP30P140LVT U9227 ( .A1(i_data_bus[268]), .A2(n10415), .B1(
        i_data_bus[300]), .B2(n10414), .ZN(n6281) );
  ND2D1BWP30P140LVT U9228 ( .A1(n6282), .A2(n6281), .ZN(N14133) );
  NR4D1BWP30P140LVT U9229 ( .A1(i_cmd[125]), .A2(n6283), .A3(n9760), .A4(n6285), .ZN(n10474) );
  INR4D1BWP30P140LVT U9230 ( .A1(i_cmd[101]), .B1(i_cmd[117]), .B2(n9758), 
        .B3(n6284), .ZN(n10473) );
  AOI22D1BWP30P140LVT U9231 ( .A1(i_data_bus[422]), .A2(n10474), .B1(
        i_data_bus[390]), .B2(n10473), .ZN(n6288) );
  INR4D1BWP30P140LVT U9232 ( .A1(i_cmd[117]), .B1(i_cmd[101]), .B2(n9761), 
        .B3(n6284), .ZN(n10476) );
  NR4D1BWP30P140LVT U9233 ( .A1(i_cmd[109]), .A2(n9764), .A3(n6286), .A4(n6285), .ZN(n10475) );
  AOI22D1BWP30P140LVT U9234 ( .A1(i_data_bus[454]), .A2(n10476), .B1(
        i_data_bus[486]), .B2(n10475), .ZN(n6287) );
  ND2D1BWP30P140LVT U9235 ( .A1(n6288), .A2(n6287), .ZN(N10595) );
  AOI22D1BWP30P140LVT U9236 ( .A1(i_data_bus[336]), .A2(n10413), .B1(
        i_data_bus[272]), .B2(n10415), .ZN(n6290) );
  AOI22D1BWP30P140LVT U9237 ( .A1(i_data_bus[368]), .A2(n10416), .B1(
        i_data_bus[304]), .B2(n10414), .ZN(n6289) );
  ND2D1BWP30P140LVT U9238 ( .A1(n6290), .A2(n6289), .ZN(N14137) );
  AOI22D1BWP30P140LVT U9239 ( .A1(i_data_bus[365]), .A2(n10416), .B1(
        i_data_bus[269]), .B2(n10415), .ZN(n6292) );
  AOI22D1BWP30P140LVT U9240 ( .A1(i_data_bus[333]), .A2(n10413), .B1(
        i_data_bus[301]), .B2(n10414), .ZN(n6291) );
  ND2D1BWP30P140LVT U9241 ( .A1(n6292), .A2(n6291), .ZN(N14134) );
  INR4D1BWP30P140LVT U9242 ( .A1(i_cmd[111]), .B1(i_cmd[127]), .B2(n9760), 
        .B3(n6293), .ZN(n10411) );
  INR4D1BWP30P140LVT U9243 ( .A1(i_cmd[127]), .B1(i_cmd[111]), .B2(n9764), 
        .B3(n6293), .ZN(n10412) );
  AOI22D1BWP30P140LVT U9244 ( .A1(i_data_bus[447]), .A2(n10411), .B1(
        i_data_bus[511]), .B2(n10412), .ZN(n6298) );
  NR4D1BWP30P140LVT U9245 ( .A1(i_cmd[103]), .A2(n6294), .A3(n9761), .A4(n6295), .ZN(n10410) );
  NR4D1BWP30P140LVT U9246 ( .A1(i_cmd[119]), .A2(n9758), .A3(n6296), .A4(n6295), .ZN(n10409) );
  AOI22D1BWP30P140LVT U9247 ( .A1(i_data_bus[479]), .A2(n10410), .B1(
        i_data_bus[415]), .B2(n10409), .ZN(n6297) );
  ND2D1BWP30P140LVT U9248 ( .A1(n6298), .A2(n6297), .ZN(N14368) );
  NR4D1BWP30P140LVT U9249 ( .A1(i_cmd[121]), .A2(n6299), .A3(n9760), .A4(n6301), .ZN(n10601) );
  INR4D1BWP30P140LVT U9250 ( .A1(i_cmd[97]), .B1(i_cmd[113]), .B2(n9758), .B3(
        n6300), .ZN(n10603) );
  AOI22D1BWP30P140LVT U9251 ( .A1(i_data_bus[422]), .A2(n10601), .B1(
        i_data_bus[390]), .B2(n10603), .ZN(n6304) );
  INR4D1BWP30P140LVT U9252 ( .A1(i_cmd[113]), .B1(i_cmd[97]), .B2(n9761), .B3(
        n6300), .ZN(n10604) );
  NR4D1BWP30P140LVT U9253 ( .A1(i_cmd[105]), .A2(n9764), .A3(n6302), .A4(n6301), .ZN(n10602) );
  AOI22D1BWP30P140LVT U9254 ( .A1(i_data_bus[454]), .A2(n10604), .B1(
        i_data_bus[486]), .B2(n10602), .ZN(n6303) );
  ND2D1BWP30P140LVT U9255 ( .A1(n6304), .A2(n6303), .ZN(N3099) );
  AOI22D1BWP30P140LVT U9256 ( .A1(i_data_bus[479]), .A2(n10604), .B1(
        i_data_bus[415]), .B2(n10603), .ZN(n6306) );
  AOI22D1BWP30P140LVT U9257 ( .A1(i_data_bus[447]), .A2(n10601), .B1(
        i_data_bus[511]), .B2(n10602), .ZN(n6305) );
  ND2D1BWP30P140LVT U9258 ( .A1(n6306), .A2(n6305), .ZN(N3124) );
  AOI22D1BWP30P140LVT U9259 ( .A1(i_data_bus[471]), .A2(n10604), .B1(
        i_data_bus[407]), .B2(n10603), .ZN(n6308) );
  AOI22D1BWP30P140LVT U9260 ( .A1(i_data_bus[439]), .A2(n10601), .B1(
        i_data_bus[503]), .B2(n10602), .ZN(n6307) );
  ND2D1BWP30P140LVT U9261 ( .A1(n6308), .A2(n6307), .ZN(N3116) );
  AOI22D1BWP30P140LVT U9262 ( .A1(i_data_bus[203]), .A2(n10610), .B1(
        i_data_bus[139]), .B2(n10612), .ZN(n6310) );
  AOI22D1BWP30P140LVT U9263 ( .A1(i_data_bus[235]), .A2(n10611), .B1(
        i_data_bus[171]), .B2(n10609), .ZN(n6309) );
  ND2D1BWP30P140LVT U9264 ( .A1(n6310), .A2(n6309), .ZN(N2672) );
  AOI22D1BWP30P140LVT U9265 ( .A1(i_data_bus[156]), .A2(n10612), .B1(
        i_data_bus[220]), .B2(n10610), .ZN(n6312) );
  AOI22D1BWP30P140LVT U9266 ( .A1(i_data_bus[252]), .A2(n10611), .B1(
        i_data_bus[188]), .B2(n10609), .ZN(n6311) );
  ND2D1BWP30P140LVT U9267 ( .A1(n6312), .A2(n6311), .ZN(N2689) );
  AOI22D1BWP30P140LVT U9268 ( .A1(i_data_bus[229]), .A2(n10611), .B1(
        i_data_bus[197]), .B2(n10610), .ZN(n6314) );
  AOI22D1BWP30P140LVT U9269 ( .A1(i_data_bus[133]), .A2(n10612), .B1(
        i_data_bus[165]), .B2(n10609), .ZN(n6313) );
  ND2D1BWP30P140LVT U9270 ( .A1(n6314), .A2(n6313), .ZN(N2666) );
  AOI22D1BWP30P140LVT U9271 ( .A1(i_data_bus[248]), .A2(n10611), .B1(
        i_data_bus[152]), .B2(n10612), .ZN(n6316) );
  AOI22D1BWP30P140LVT U9272 ( .A1(i_data_bus[216]), .A2(n10610), .B1(
        i_data_bus[184]), .B2(n10609), .ZN(n6315) );
  ND2D1BWP30P140LVT U9273 ( .A1(n6316), .A2(n6315), .ZN(N2685) );
  INR4D1BWP30P140LVT U9274 ( .A1(i_cmd[37]), .B1(i_cmd[53]), .B2(n9857), .B3(
        n6317), .ZN(n10481) );
  INR4D1BWP30P140LVT U9275 ( .A1(i_cmd[53]), .B1(i_cmd[37]), .B2(n9854), .B3(
        n6317), .ZN(n10482) );
  AOI22D1BWP30P140LVT U9276 ( .A1(i_data_bus[128]), .A2(n10481), .B1(
        i_data_bus[192]), .B2(n10482), .ZN(n6322) );
  NR4D1BWP30P140LVT U9277 ( .A1(i_cmd[45]), .A2(n6318), .A3(n9860), .A4(n6319), 
        .ZN(n10484) );
  NR4D1BWP30P140LVT U9278 ( .A1(i_cmd[61]), .A2(n9853), .A3(n6320), .A4(n6319), 
        .ZN(n10483) );
  AOI22D1BWP30P140LVT U9279 ( .A1(i_data_bus[224]), .A2(n10484), .B1(
        i_data_bus[160]), .B2(n10483), .ZN(n6321) );
  ND2D1BWP30P140LVT U9280 ( .A1(n6322), .A2(n6321), .ZN(N10157) );
  AOI22D1BWP30P140LVT U9281 ( .A1(i_data_bus[156]), .A2(n10481), .B1(
        i_data_bus[220]), .B2(n10482), .ZN(n6324) );
  AOI22D1BWP30P140LVT U9282 ( .A1(i_data_bus[252]), .A2(n10484), .B1(
        i_data_bus[188]), .B2(n10483), .ZN(n6323) );
  ND2D1BWP30P140LVT U9283 ( .A1(n6324), .A2(n6323), .ZN(N10185) );
  INR4D1BWP30P140LVT U9284 ( .A1(i_cmd[213]), .B1(i_cmd[197]), .B2(n9741), 
        .B3(n6326), .ZN(n10463) );
  NR4D1BWP30P140LVT U9285 ( .A1(i_cmd[221]), .A2(n9743), .A3(n6325), .A4(n6327), .ZN(n10464) );
  AOI22D1BWP30P140LVT U9286 ( .A1(i_data_bus[843]), .A2(n10463), .B1(
        i_data_bus[811]), .B2(n10464), .ZN(n6330) );
  INR4D1BWP30P140LVT U9287 ( .A1(i_cmd[197]), .B1(i_cmd[213]), .B2(n9744), 
        .B3(n6326), .ZN(n10462) );
  NR4D1BWP30P140LVT U9288 ( .A1(i_cmd[205]), .A2(n6328), .A3(n9747), .A4(n6327), .ZN(n10461) );
  AOI22D1BWP30P140LVT U9289 ( .A1(i_data_bus[779]), .A2(n10462), .B1(
        i_data_bus[875]), .B2(n10461), .ZN(n6329) );
  ND2D1BWP30P140LVT U9290 ( .A1(n6330), .A2(n6329), .ZN(N11248) );
  AOI22D1BWP30P140LVT U9291 ( .A1(i_data_bus[454]), .A2(n10508), .B1(
        i_data_bus[390]), .B2(n10505), .ZN(n6332) );
  AOI22D1BWP30P140LVT U9292 ( .A1(i_data_bus[422]), .A2(n10507), .B1(
        i_data_bus[486]), .B2(n10506), .ZN(n6331) );
  ND2D1BWP30P140LVT U9293 ( .A1(n6332), .A2(n6331), .ZN(N8721) );
  AOI22D1BWP30P140LVT U9294 ( .A1(i_data_bus[479]), .A2(n10508), .B1(
        i_data_bus[415]), .B2(n10505), .ZN(n6334) );
  AOI22D1BWP30P140LVT U9295 ( .A1(i_data_bus[447]), .A2(n10507), .B1(
        i_data_bus[511]), .B2(n10506), .ZN(n6333) );
  ND2D1BWP30P140LVT U9296 ( .A1(n6334), .A2(n6333), .ZN(N8746) );
  AOI22D1BWP30P140LVT U9297 ( .A1(i_data_bus[409]), .A2(n10572), .B1(
        i_data_bus[441]), .B2(n10569), .ZN(n6336) );
  AOI22D1BWP30P140LVT U9298 ( .A1(i_data_bus[473]), .A2(n10570), .B1(
        i_data_bus[505]), .B2(n10571), .ZN(n6335) );
  ND2D1BWP30P140LVT U9299 ( .A1(n6336), .A2(n6335), .ZN(N4992) );
  AOI22D1BWP30P140LVT U9300 ( .A1(i_data_bus[408]), .A2(n10572), .B1(
        i_data_bus[440]), .B2(n10569), .ZN(n6338) );
  AOI22D1BWP30P140LVT U9301 ( .A1(i_data_bus[472]), .A2(n10570), .B1(
        i_data_bus[504]), .B2(n10571), .ZN(n6337) );
  ND2D1BWP30P140LVT U9302 ( .A1(n6338), .A2(n6337), .ZN(N4991) );
  AOI22D1BWP30P140LVT U9303 ( .A1(i_data_bus[398]), .A2(n10572), .B1(
        i_data_bus[462]), .B2(n10570), .ZN(n6340) );
  AOI22D1BWP30P140LVT U9304 ( .A1(i_data_bus[430]), .A2(n10569), .B1(
        i_data_bus[494]), .B2(n10571), .ZN(n6339) );
  ND2D1BWP30P140LVT U9305 ( .A1(n6340), .A2(n6339), .ZN(N4981) );
  AOI22D1BWP30P140LVT U9306 ( .A1(i_data_bus[416]), .A2(n10569), .B1(
        i_data_bus[448]), .B2(n10570), .ZN(n6342) );
  AOI22D1BWP30P140LVT U9307 ( .A1(i_data_bus[384]), .A2(n10572), .B1(
        i_data_bus[480]), .B2(n10571), .ZN(n6341) );
  ND2D1BWP30P140LVT U9308 ( .A1(n6342), .A2(n6341), .ZN(N4967) );
  AOI22D1BWP30P140LVT U9309 ( .A1(i_data_bus[405]), .A2(n10572), .B1(
        i_data_bus[469]), .B2(n10570), .ZN(n6344) );
  AOI22D1BWP30P140LVT U9310 ( .A1(i_data_bus[437]), .A2(n10569), .B1(
        i_data_bus[501]), .B2(n10571), .ZN(n6343) );
  ND2D1BWP30P140LVT U9311 ( .A1(n6344), .A2(n6343), .ZN(N4988) );
  AOI22D1BWP30P140LVT U9312 ( .A1(i_data_bus[411]), .A2(n10572), .B1(
        i_data_bus[475]), .B2(n10570), .ZN(n6346) );
  AOI22D1BWP30P140LVT U9313 ( .A1(i_data_bus[443]), .A2(n10569), .B1(
        i_data_bus[507]), .B2(n10571), .ZN(n6345) );
  ND2D1BWP30P140LVT U9314 ( .A1(n6346), .A2(n6345), .ZN(N4994) );
  AOI22D1BWP30P140LVT U9315 ( .A1(i_data_bus[388]), .A2(n10572), .B1(
        i_data_bus[420]), .B2(n10569), .ZN(n6348) );
  AOI22D1BWP30P140LVT U9316 ( .A1(i_data_bus[452]), .A2(n10570), .B1(
        i_data_bus[484]), .B2(n10571), .ZN(n6347) );
  ND2D1BWP30P140LVT U9317 ( .A1(n6348), .A2(n6347), .ZN(N4971) );
  AOI22D1BWP30P140LVT U9318 ( .A1(i_data_bus[385]), .A2(n10572), .B1(
        i_data_bus[449]), .B2(n10570), .ZN(n6350) );
  AOI22D1BWP30P140LVT U9319 ( .A1(i_data_bus[417]), .A2(n10569), .B1(
        i_data_bus[481]), .B2(n10571), .ZN(n6349) );
  ND2D1BWP30P140LVT U9320 ( .A1(n6350), .A2(n6349), .ZN(N4968) );
  AOI22D1BWP30P140LVT U9321 ( .A1(i_data_bus[427]), .A2(n10569), .B1(
        i_data_bus[459]), .B2(n10570), .ZN(n6352) );
  AOI22D1BWP30P140LVT U9322 ( .A1(i_data_bus[395]), .A2(n10572), .B1(
        i_data_bus[491]), .B2(n10571), .ZN(n6351) );
  ND2D1BWP30P140LVT U9323 ( .A1(n6352), .A2(n6351), .ZN(N4978) );
  AOI22D1BWP30P140LVT U9324 ( .A1(i_data_bus[439]), .A2(n10569), .B1(
        i_data_bus[407]), .B2(n10572), .ZN(n6354) );
  AOI22D1BWP30P140LVT U9325 ( .A1(i_data_bus[471]), .A2(n10570), .B1(
        i_data_bus[503]), .B2(n10571), .ZN(n6353) );
  ND2D1BWP30P140LVT U9326 ( .A1(n6354), .A2(n6353), .ZN(N4990) );
  AOI22D1BWP30P140LVT U9327 ( .A1(i_data_bus[422]), .A2(n10569), .B1(
        i_data_bus[390]), .B2(n10572), .ZN(n6356) );
  AOI22D1BWP30P140LVT U9328 ( .A1(i_data_bus[454]), .A2(n10570), .B1(
        i_data_bus[486]), .B2(n10571), .ZN(n6355) );
  ND2D1BWP30P140LVT U9329 ( .A1(n6356), .A2(n6355), .ZN(N4973) );
  INR4D1BWP30P140LVT U9330 ( .A1(i_cmd[194]), .B1(i_cmd[210]), .B2(n9744), 
        .B3(n6357), .ZN(n10558) );
  INR4D1BWP30P140LVT U9331 ( .A1(i_cmd[210]), .B1(i_cmd[194]), .B2(n9741), 
        .B3(n6357), .ZN(n10557) );
  AOI22D1BWP30P140LVT U9332 ( .A1(i_data_bus[780]), .A2(n10558), .B1(
        i_data_bus[844]), .B2(n10557), .ZN(n6362) );
  NR4D1BWP30P140LVT U9333 ( .A1(i_cmd[218]), .A2(n6360), .A3(n9743), .A4(n6358), .ZN(n10560) );
  NR4D1BWP30P140LVT U9334 ( .A1(i_cmd[202]), .A2(n6360), .A3(n9747), .A4(n6359), .ZN(n10559) );
  AOI22D1BWP30P140LVT U9335 ( .A1(i_data_bus[812]), .A2(n10560), .B1(
        i_data_bus[876]), .B2(n10559), .ZN(n6361) );
  ND2D1BWP30P140LVT U9336 ( .A1(n6362), .A2(n6361), .ZN(N5627) );
  AOI22D1BWP30P140LVT U9337 ( .A1(i_data_bus[476]), .A2(n10410), .B1(
        i_data_bus[412]), .B2(n10409), .ZN(n6364) );
  AOI22D1BWP30P140LVT U9338 ( .A1(i_data_bus[444]), .A2(n10411), .B1(
        i_data_bus[508]), .B2(n10412), .ZN(n6363) );
  ND2D1BWP30P140LVT U9339 ( .A1(n6364), .A2(n6363), .ZN(N14365) );
  AOI22D1BWP30P140LVT U9340 ( .A1(i_data_bus[422]), .A2(n10411), .B1(
        i_data_bus[390]), .B2(n10409), .ZN(n6366) );
  AOI22D1BWP30P140LVT U9341 ( .A1(i_data_bus[454]), .A2(n10410), .B1(
        i_data_bus[486]), .B2(n10412), .ZN(n6365) );
  ND2D1BWP30P140LVT U9342 ( .A1(n6366), .A2(n6365), .ZN(N14343) );
  NR4D1BWP30P140LVT U9343 ( .A1(i_cmd[55]), .A2(n6367), .A3(n9857), .A4(n6369), 
        .ZN(n10417) );
  INR4D1BWP30P140LVT U9344 ( .A1(i_cmd[47]), .B1(i_cmd[63]), .B2(n9853), .B3(
        n6368), .ZN(n10420) );
  AOI22D1BWP30P140LVT U9345 ( .A1(i_data_bus[156]), .A2(n10417), .B1(
        i_data_bus[188]), .B2(n10420), .ZN(n6372) );
  INR4D1BWP30P140LVT U9346 ( .A1(i_cmd[63]), .B1(i_cmd[47]), .B2(n9860), .B3(
        n6368), .ZN(n10418) );
  NR4D1BWP30P140LVT U9347 ( .A1(i_cmd[39]), .A2(n9854), .A3(n6370), .A4(n6369), 
        .ZN(n10419) );
  AOI22D1BWP30P140LVT U9348 ( .A1(i_data_bus[252]), .A2(n10418), .B1(
        i_data_bus[220]), .B2(n10419), .ZN(n6371) );
  ND2D1BWP30P140LVT U9349 ( .A1(n6372), .A2(n6371), .ZN(N13933) );
  AOI22D1BWP30P140LVT U9350 ( .A1(i_data_bus[228]), .A2(n10418), .B1(
        i_data_bus[164]), .B2(n10420), .ZN(n6374) );
  AOI22D1BWP30P140LVT U9351 ( .A1(i_data_bus[132]), .A2(n10417), .B1(
        i_data_bus[196]), .B2(n10419), .ZN(n6373) );
  ND2D1BWP30P140LVT U9352 ( .A1(n6374), .A2(n6373), .ZN(N13909) );
  INR4D1BWP30P140LVT U9353 ( .A1(i_cmd[60]), .B1(i_cmd[44]), .B2(n9860), .B3(
        n6375), .ZN(n10516) );
  INR4D1BWP30P140LVT U9354 ( .A1(i_cmd[44]), .B1(i_cmd[60]), .B2(n9853), .B3(
        n6375), .ZN(n10515) );
  AOI22D1BWP30P140LVT U9355 ( .A1(i_data_bus[228]), .A2(n10516), .B1(
        i_data_bus[164]), .B2(n10515), .ZN(n6380) );
  NR4D1BWP30P140LVT U9356 ( .A1(i_cmd[52]), .A2(n6376), .A3(n9857), .A4(n6377), 
        .ZN(n10513) );
  NR4D1BWP30P140LVT U9357 ( .A1(i_cmd[36]), .A2(n9854), .A3(n6378), .A4(n6377), 
        .ZN(n10514) );
  AOI22D1BWP30P140LVT U9358 ( .A1(i_data_bus[132]), .A2(n10513), .B1(
        i_data_bus[196]), .B2(n10514), .ZN(n6379) );
  ND2D1BWP30P140LVT U9359 ( .A1(n6380), .A2(n6379), .ZN(N8287) );
  INR4D1BWP30P140LVT U9360 ( .A1(i_cmd[86]), .B1(i_cmd[70]), .B2(n9807), .B3(
        n6381), .ZN(n10446) );
  INR4D1BWP30P140LVT U9361 ( .A1(i_cmd[70]), .B1(i_cmd[86]), .B2(n9808), .B3(
        n6381), .ZN(n10447) );
  AOI22D1BWP30P140LVT U9362 ( .A1(i_data_bus[338]), .A2(n10446), .B1(
        i_data_bus[274]), .B2(n10447), .ZN(n6386) );
  NR4D1BWP30P140LVT U9363 ( .A1(i_cmd[78]), .A2(n6382), .A3(n9812), .A4(n6383), 
        .ZN(n10445) );
  NR4D1BWP30P140LVT U9364 ( .A1(i_cmd[94]), .A2(n9813), .A3(n6384), .A4(n6383), 
        .ZN(n10448) );
  AOI22D1BWP30P140LVT U9365 ( .A1(i_data_bus[370]), .A2(n10445), .B1(
        i_data_bus[306]), .B2(n10448), .ZN(n6385) );
  ND2D1BWP30P140LVT U9366 ( .A1(n6386), .A2(n6385), .ZN(N12265) );
  AOI22D1BWP30P140LVT U9367 ( .A1(i_data_bus[350]), .A2(n10446), .B1(
        i_data_bus[286]), .B2(n10447), .ZN(n6388) );
  AOI22D1BWP30P140LVT U9368 ( .A1(i_data_bus[382]), .A2(n10445), .B1(
        i_data_bus[318]), .B2(n10448), .ZN(n6387) );
  ND2D1BWP30P140LVT U9369 ( .A1(n6388), .A2(n6387), .ZN(N12277) );
  AOI22D1BWP30P140LVT U9370 ( .A1(i_data_bus[340]), .A2(n10446), .B1(
        i_data_bus[276]), .B2(n10447), .ZN(n6390) );
  AOI22D1BWP30P140LVT U9371 ( .A1(i_data_bus[372]), .A2(n10445), .B1(
        i_data_bus[308]), .B2(n10448), .ZN(n6389) );
  ND2D1BWP30P140LVT U9372 ( .A1(n6390), .A2(n6389), .ZN(N12267) );
  AOI22D1BWP30P140LVT U9373 ( .A1(i_data_bus[673]), .A2(n10404), .B1(
        i_data_bus[705]), .B2(n10402), .ZN(n6392) );
  AOI22D1BWP30P140LVT U9374 ( .A1(i_data_bus[641]), .A2(n10401), .B1(
        i_data_bus[737]), .B2(n10403), .ZN(n6391) );
  ND2D1BWP30P140LVT U9375 ( .A1(n6392), .A2(n6391), .ZN(N14770) );
  AOI22D1BWP30P140LVT U9376 ( .A1(i_data_bus[409]), .A2(n10441), .B1(
        i_data_bus[441]), .B2(n10443), .ZN(n6394) );
  AOI22D1BWP30P140LVT U9377 ( .A1(i_data_bus[473]), .A2(n10442), .B1(
        i_data_bus[505]), .B2(n10444), .ZN(n6393) );
  ND2D1BWP30P140LVT U9378 ( .A1(n6394), .A2(n6393), .ZN(N12488) );
  AOI22D1BWP30P140LVT U9379 ( .A1(i_data_bus[394]), .A2(n10441), .B1(
        i_data_bus[426]), .B2(n10443), .ZN(n6396) );
  AOI22D1BWP30P140LVT U9380 ( .A1(i_data_bus[458]), .A2(n10442), .B1(
        i_data_bus[490]), .B2(n10444), .ZN(n6395) );
  ND2D1BWP30P140LVT U9381 ( .A1(n6396), .A2(n6395), .ZN(N12473) );
  AOI22D1BWP30P140LVT U9382 ( .A1(i_data_bus[472]), .A2(n10442), .B1(
        i_data_bus[440]), .B2(n10443), .ZN(n6398) );
  AOI22D1BWP30P140LVT U9383 ( .A1(i_data_bus[408]), .A2(n10441), .B1(
        i_data_bus[504]), .B2(n10444), .ZN(n6397) );
  ND2D1BWP30P140LVT U9384 ( .A1(n6398), .A2(n6397), .ZN(N12487) );
  NR4D1BWP30P140LVT U9385 ( .A1(i_cmd[65]), .A2(n6399), .A3(n9807), .A4(n6401), 
        .ZN(n10607) );
  INR4D1BWP30P140LVT U9386 ( .A1(i_cmd[73]), .B1(i_cmd[89]), .B2(n9813), .B3(
        n6400), .ZN(n10606) );
  AOI22D1BWP30P140LVT U9387 ( .A1(i_data_bus[348]), .A2(n10607), .B1(
        i_data_bus[316]), .B2(n10606), .ZN(n6404) );
  INR4D1BWP30P140LVT U9388 ( .A1(i_cmd[89]), .B1(i_cmd[73]), .B2(n9812), .B3(
        n6400), .ZN(n10608) );
  NR4D1BWP30P140LVT U9389 ( .A1(i_cmd[81]), .A2(n9808), .A3(n6402), .A4(n6401), 
        .ZN(n10605) );
  AOI22D1BWP30P140LVT U9390 ( .A1(i_data_bus[380]), .A2(n10608), .B1(
        i_data_bus[284]), .B2(n10605), .ZN(n6403) );
  ND2D1BWP30P140LVT U9391 ( .A1(n6404), .A2(n6403), .ZN(N2905) );
  AOI22D1BWP30P140LVT U9392 ( .A1(i_data_bus[350]), .A2(n10607), .B1(
        i_data_bus[318]), .B2(n10606), .ZN(n6406) );
  AOI22D1BWP30P140LVT U9393 ( .A1(i_data_bus[382]), .A2(n10608), .B1(
        i_data_bus[286]), .B2(n10605), .ZN(n6405) );
  ND2D1BWP30P140LVT U9394 ( .A1(n6406), .A2(n6405), .ZN(N2907) );
  AOI22D1BWP30P140LVT U9395 ( .A1(i_data_bus[368]), .A2(n10608), .B1(
        i_data_bus[304]), .B2(n10606), .ZN(n6408) );
  AOI22D1BWP30P140LVT U9396 ( .A1(i_data_bus[336]), .A2(n10607), .B1(
        i_data_bus[272]), .B2(n10605), .ZN(n6407) );
  ND2D1BWP30P140LVT U9397 ( .A1(n6408), .A2(n6407), .ZN(N2893) );
  NR4D1BWP30P140LVT U9398 ( .A1(i_cmd[77]), .A2(n6409), .A3(n9812), .A4(n6411), 
        .ZN(n10479) );
  INR4D1BWP30P140LVT U9399 ( .A1(i_cmd[85]), .B1(i_cmd[69]), .B2(n9807), .B3(
        n6410), .ZN(n10478) );
  AOI22D1BWP30P140LVT U9400 ( .A1(i_data_bus[364]), .A2(n10479), .B1(
        i_data_bus[332]), .B2(n10478), .ZN(n6414) );
  INR4D1BWP30P140LVT U9401 ( .A1(i_cmd[69]), .B1(i_cmd[85]), .B2(n9808), .B3(
        n6410), .ZN(n10480) );
  NR4D1BWP30P140LVT U9402 ( .A1(i_cmd[93]), .A2(n9813), .A3(n6412), .A4(n6411), 
        .ZN(n10477) );
  AOI22D1BWP30P140LVT U9403 ( .A1(i_data_bus[268]), .A2(n10480), .B1(
        i_data_bus[300]), .B2(n10477), .ZN(n6413) );
  ND2D1BWP30P140LVT U9404 ( .A1(n6414), .A2(n6413), .ZN(N10385) );
  AOI22D1BWP30P140LVT U9405 ( .A1(i_data_bus[128]), .A2(n10417), .B1(
        i_data_bus[224]), .B2(n10418), .ZN(n6416) );
  AOI22D1BWP30P140LVT U9406 ( .A1(i_data_bus[160]), .A2(n10420), .B1(
        i_data_bus[192]), .B2(n10419), .ZN(n6415) );
  ND2D1BWP30P140LVT U9407 ( .A1(n6416), .A2(n6415), .ZN(N13905) );
  AOI22D1BWP30P140LVT U9408 ( .A1(i_data_bus[363]), .A2(n10445), .B1(
        i_data_bus[331]), .B2(n10446), .ZN(n6418) );
  AOI22D1BWP30P140LVT U9409 ( .A1(i_data_bus[267]), .A2(n10447), .B1(
        i_data_bus[299]), .B2(n10448), .ZN(n6417) );
  ND2D1BWP30P140LVT U9410 ( .A1(n6418), .A2(n6417), .ZN(N12258) );
  AOI22D1BWP30P140LVT U9411 ( .A1(i_data_bus[268]), .A2(n10447), .B1(
        i_data_bus[332]), .B2(n10446), .ZN(n6420) );
  AOI22D1BWP30P140LVT U9412 ( .A1(i_data_bus[364]), .A2(n10445), .B1(
        i_data_bus[300]), .B2(n10448), .ZN(n6419) );
  ND2D1BWP30P140LVT U9413 ( .A1(n6420), .A2(n6419), .ZN(N12259) );
  AOI22D1BWP30P140LVT U9414 ( .A1(i_data_bus[990]), .A2(n10426), .B1(
        i_data_bus[1022]), .B2(n10427), .ZN(n6422) );
  AOI22D1BWP30P140LVT U9415 ( .A1(i_data_bus[958]), .A2(n10428), .B1(
        i_data_bus[926]), .B2(n10425), .ZN(n6421) );
  ND2D1BWP30P140LVT U9416 ( .A1(n6422), .A2(n6421), .ZN(N13357) );
  AOI22D1BWP30P140LVT U9417 ( .A1(i_data_bus[978]), .A2(n10426), .B1(
        i_data_bus[946]), .B2(n10428), .ZN(n6424) );
  AOI22D1BWP30P140LVT U9418 ( .A1(i_data_bus[1010]), .A2(n10427), .B1(
        i_data_bus[914]), .B2(n10425), .ZN(n6423) );
  ND2D1BWP30P140LVT U9419 ( .A1(n6424), .A2(n6423), .ZN(N13345) );
  AOI22D1BWP30P140LVT U9420 ( .A1(i_data_bus[936]), .A2(n10428), .B1(
        i_data_bus[1000]), .B2(n10427), .ZN(n6426) );
  AOI22D1BWP30P140LVT U9421 ( .A1(i_data_bus[968]), .A2(n10426), .B1(
        i_data_bus[904]), .B2(n10425), .ZN(n6425) );
  ND2D1BWP30P140LVT U9422 ( .A1(n6426), .A2(n6425), .ZN(N13335) );
  AOI22D1BWP30P140LVT U9423 ( .A1(i_data_bus[408]), .A2(n10473), .B1(
        i_data_bus[472]), .B2(n10476), .ZN(n6428) );
  AOI22D1BWP30P140LVT U9424 ( .A1(i_data_bus[440]), .A2(n10474), .B1(
        i_data_bus[504]), .B2(n10475), .ZN(n6427) );
  ND2D1BWP30P140LVT U9425 ( .A1(n6428), .A2(n6427), .ZN(N10613) );
  AOI22D1BWP30P140LVT U9426 ( .A1(i_data_bus[429]), .A2(n10474), .B1(
        i_data_bus[461]), .B2(n10476), .ZN(n6430) );
  AOI22D1BWP30P140LVT U9427 ( .A1(i_data_bus[397]), .A2(n10473), .B1(
        i_data_bus[493]), .B2(n10475), .ZN(n6429) );
  ND2D1BWP30P140LVT U9428 ( .A1(n6430), .A2(n6429), .ZN(N10602) );
  INR4D1BWP30P140LVT U9429 ( .A1(i_cmd[20]), .B1(i_cmd[4]), .B2(n10014), .B3(
        n6432), .ZN(n10517) );
  NR4D1BWP30P140LVT U9430 ( .A1(i_cmd[12]), .A2(n6431), .A3(n10019), .A4(n6433), .ZN(n10519) );
  AOI22D1BWP30P140LVT U9431 ( .A1(i_data_bus[73]), .A2(n10517), .B1(
        i_data_bus[105]), .B2(n10519), .ZN(n6436) );
  INR4D1BWP30P140LVT U9432 ( .A1(i_cmd[4]), .B1(i_cmd[20]), .B2(n10013), .B3(
        n6432), .ZN(n10520) );
  NR4D1BWP30P140LVT U9433 ( .A1(i_cmd[28]), .A2(n10018), .A3(n6434), .A4(n6433), .ZN(n10518) );
  AOI22D1BWP30P140LVT U9434 ( .A1(i_data_bus[9]), .A2(n10520), .B1(
        i_data_bus[41]), .B2(n10518), .ZN(n6435) );
  ND2D1BWP30P140LVT U9435 ( .A1(n6436), .A2(n6435), .ZN(N8076) );
  AOI22D1BWP30P140LVT U9436 ( .A1(i_data_bus[114]), .A2(n10519), .B1(
        i_data_bus[82]), .B2(n10517), .ZN(n6438) );
  AOI22D1BWP30P140LVT U9437 ( .A1(i_data_bus[18]), .A2(n10520), .B1(
        i_data_bus[50]), .B2(n10518), .ZN(n6437) );
  ND2D1BWP30P140LVT U9438 ( .A1(n6438), .A2(n6437), .ZN(N8085) );
  AOI22D1BWP30P140LVT U9439 ( .A1(i_data_bus[15]), .A2(n10520), .B1(
        i_data_bus[79]), .B2(n10517), .ZN(n6440) );
  AOI22D1BWP30P140LVT U9440 ( .A1(i_data_bus[111]), .A2(n10519), .B1(
        i_data_bus[47]), .B2(n10518), .ZN(n6439) );
  ND2D1BWP30P140LVT U9441 ( .A1(n6440), .A2(n6439), .ZN(N8082) );
  INR4D1BWP30P140LVT U9442 ( .A1(i_cmd[193]), .B1(i_cmd[209]), .B2(n9744), 
        .B3(n6441), .ZN(n10589) );
  INR4D1BWP30P140LVT U9443 ( .A1(i_cmd[209]), .B1(i_cmd[193]), .B2(n9741), 
        .B3(n6441), .ZN(n10590) );
  AOI22D1BWP30P140LVT U9444 ( .A1(i_data_bus[769]), .A2(n10589), .B1(
        i_data_bus[833]), .B2(n10590), .ZN(n6446) );
  NR4D1BWP30P140LVT U9445 ( .A1(i_cmd[217]), .A2(n6444), .A3(n9743), .A4(n6442), .ZN(n10592) );
  NR4D1BWP30P140LVT U9446 ( .A1(i_cmd[201]), .A2(n6444), .A3(n9747), .A4(n6443), .ZN(n10591) );
  AOI22D1BWP30P140LVT U9447 ( .A1(i_data_bus[801]), .A2(n10592), .B1(
        i_data_bus[865]), .B2(n10591), .ZN(n6445) );
  ND2D1BWP30P140LVT U9448 ( .A1(n6446), .A2(n6445), .ZN(N3742) );
  AOI22D1BWP30P140LVT U9449 ( .A1(i_data_bus[788]), .A2(n10589), .B1(
        i_data_bus[852]), .B2(n10590), .ZN(n6448) );
  AOI22D1BWP30P140LVT U9450 ( .A1(i_data_bus[820]), .A2(n10592), .B1(
        i_data_bus[884]), .B2(n10591), .ZN(n6447) );
  ND2D1BWP30P140LVT U9451 ( .A1(n6448), .A2(n6447), .ZN(N3761) );
  AOI22D1BWP30P140LVT U9452 ( .A1(i_data_bus[860]), .A2(n10463), .B1(
        i_data_bus[796]), .B2(n10462), .ZN(n6450) );
  AOI22D1BWP30P140LVT U9453 ( .A1(i_data_bus[828]), .A2(n10464), .B1(
        i_data_bus[892]), .B2(n10461), .ZN(n6449) );
  ND2D1BWP30P140LVT U9454 ( .A1(n6450), .A2(n6449), .ZN(N11265) );
  AOI22D1BWP30P140LVT U9455 ( .A1(i_data_bus[825]), .A2(n10464), .B1(
        i_data_bus[793]), .B2(n10462), .ZN(n6452) );
  AOI22D1BWP30P140LVT U9456 ( .A1(i_data_bus[857]), .A2(n10463), .B1(
        i_data_bus[889]), .B2(n10461), .ZN(n6451) );
  ND2D1BWP30P140LVT U9457 ( .A1(n6452), .A2(n6451), .ZN(N11262) );
  AOI22D1BWP30P140LVT U9458 ( .A1(i_data_bus[599]), .A2(n10536), .B1(
        i_data_bus[535]), .B2(n10533), .ZN(n6454) );
  AOI22D1BWP30P140LVT U9459 ( .A1(i_data_bus[631]), .A2(n10534), .B1(
        i_data_bus[567]), .B2(n10535), .ZN(n6453) );
  ND2D1BWP30P140LVT U9460 ( .A1(n6454), .A2(n6453), .ZN(N7080) );
  AOI22D1BWP30P140LVT U9461 ( .A1(i_data_bus[516]), .A2(n10533), .B1(
        i_data_bus[580]), .B2(n10536), .ZN(n6456) );
  AOI22D1BWP30P140LVT U9462 ( .A1(i_data_bus[612]), .A2(n10534), .B1(
        i_data_bus[548]), .B2(n10535), .ZN(n6455) );
  ND2D1BWP30P140LVT U9463 ( .A1(n6456), .A2(n6455), .ZN(N7061) );
  AOI22D1BWP30P140LVT U9464 ( .A1(i_data_bus[387]), .A2(n10603), .B1(
        i_data_bus[419]), .B2(n10601), .ZN(n6458) );
  AOI22D1BWP30P140LVT U9465 ( .A1(i_data_bus[451]), .A2(n10604), .B1(
        i_data_bus[483]), .B2(n10602), .ZN(n6457) );
  ND2D1BWP30P140LVT U9466 ( .A1(n6458), .A2(n6457), .ZN(N3096) );
  AOI22D1BWP30P140LVT U9467 ( .A1(i_data_bus[394]), .A2(n10603), .B1(
        i_data_bus[426]), .B2(n10601), .ZN(n6460) );
  AOI22D1BWP30P140LVT U9468 ( .A1(i_data_bus[458]), .A2(n10604), .B1(
        i_data_bus[490]), .B2(n10602), .ZN(n6459) );
  ND2D1BWP30P140LVT U9469 ( .A1(n6460), .A2(n6459), .ZN(N3103) );
  AOI22D1BWP30P140LVT U9470 ( .A1(i_data_bus[355]), .A2(n10608), .B1(
        i_data_bus[323]), .B2(n10607), .ZN(n6462) );
  AOI22D1BWP30P140LVT U9471 ( .A1(i_data_bus[291]), .A2(n10606), .B1(
        i_data_bus[259]), .B2(n10605), .ZN(n6461) );
  ND2D1BWP30P140LVT U9472 ( .A1(n6462), .A2(n6461), .ZN(N2880) );
  AOI22D1BWP30P140LVT U9473 ( .A1(i_data_bus[315]), .A2(n10606), .B1(
        i_data_bus[347]), .B2(n10607), .ZN(n6464) );
  AOI22D1BWP30P140LVT U9474 ( .A1(i_data_bus[379]), .A2(n10608), .B1(
        i_data_bus[283]), .B2(n10605), .ZN(n6463) );
  ND2D1BWP30P140LVT U9475 ( .A1(n6464), .A2(n6463), .ZN(N2904) );
  INR4D1BWP30P140LVT U9476 ( .A1(i_cmd[68]), .B1(i_cmd[84]), .B2(n9808), .B3(
        n6465), .ZN(n10510) );
  INR4D1BWP30P140LVT U9477 ( .A1(i_cmd[84]), .B1(i_cmd[68]), .B2(n9807), .B3(
        n6465), .ZN(n10509) );
  AOI22D1BWP30P140LVT U9478 ( .A1(i_data_bus[259]), .A2(n10510), .B1(
        i_data_bus[323]), .B2(n10509), .ZN(n6470) );
  NR4D1BWP30P140LVT U9479 ( .A1(i_cmd[76]), .A2(n6466), .A3(n9812), .A4(n6467), 
        .ZN(n10511) );
  NR4D1BWP30P140LVT U9480 ( .A1(i_cmd[92]), .A2(n9813), .A3(n6468), .A4(n6467), 
        .ZN(n10512) );
  AOI22D1BWP30P140LVT U9481 ( .A1(i_data_bus[355]), .A2(n10511), .B1(
        i_data_bus[291]), .B2(n10512), .ZN(n6469) );
  ND2D1BWP30P140LVT U9482 ( .A1(n6470), .A2(n6469), .ZN(N8502) );
  AOI22D1BWP30P140LVT U9483 ( .A1(i_data_bus[336]), .A2(n10509), .B1(
        i_data_bus[272]), .B2(n10510), .ZN(n6472) );
  AOI22D1BWP30P140LVT U9484 ( .A1(i_data_bus[368]), .A2(n10511), .B1(
        i_data_bus[304]), .B2(n10512), .ZN(n6471) );
  ND2D1BWP30P140LVT U9485 ( .A1(n6472), .A2(n6471), .ZN(N8515) );
  AOI22D1BWP30P140LVT U9486 ( .A1(i_data_bus[370]), .A2(n10511), .B1(
        i_data_bus[274]), .B2(n10510), .ZN(n6474) );
  AOI22D1BWP30P140LVT U9487 ( .A1(i_data_bus[338]), .A2(n10509), .B1(
        i_data_bus[306]), .B2(n10512), .ZN(n6473) );
  ND2D1BWP30P140LVT U9488 ( .A1(n6474), .A2(n6473), .ZN(N8517) );
  AOI22D1BWP30P140LVT U9489 ( .A1(i_data_bus[320]), .A2(n10509), .B1(
        i_data_bus[256]), .B2(n10510), .ZN(n6476) );
  AOI22D1BWP30P140LVT U9490 ( .A1(i_data_bus[352]), .A2(n10511), .B1(
        i_data_bus[288]), .B2(n10512), .ZN(n6475) );
  ND2D1BWP30P140LVT U9491 ( .A1(n6476), .A2(n6475), .ZN(N8499) );
  AOI22D1BWP30P140LVT U9492 ( .A1(i_data_bus[270]), .A2(n10510), .B1(
        i_data_bus[334]), .B2(n10509), .ZN(n6478) );
  AOI22D1BWP30P140LVT U9493 ( .A1(i_data_bus[366]), .A2(n10511), .B1(
        i_data_bus[302]), .B2(n10512), .ZN(n6477) );
  ND2D1BWP30P140LVT U9494 ( .A1(n6478), .A2(n6477), .ZN(N8513) );
  AOI22D1BWP30P140LVT U9495 ( .A1(i_data_bus[365]), .A2(n10511), .B1(
        i_data_bus[333]), .B2(n10509), .ZN(n6480) );
  AOI22D1BWP30P140LVT U9496 ( .A1(i_data_bus[269]), .A2(n10510), .B1(
        i_data_bus[301]), .B2(n10512), .ZN(n6479) );
  ND2D1BWP30P140LVT U9497 ( .A1(n6480), .A2(n6479), .ZN(N8512) );
  AOI22D1BWP30P140LVT U9498 ( .A1(i_data_bus[262]), .A2(n10510), .B1(
        i_data_bus[326]), .B2(n10509), .ZN(n6482) );
  AOI22D1BWP30P140LVT U9499 ( .A1(i_data_bus[358]), .A2(n10511), .B1(
        i_data_bus[294]), .B2(n10512), .ZN(n6481) );
  ND2D1BWP30P140LVT U9500 ( .A1(n6482), .A2(n6481), .ZN(N8505) );
  AOI22D1BWP30P140LVT U9501 ( .A1(i_data_bus[325]), .A2(n10509), .B1(
        i_data_bus[261]), .B2(n10510), .ZN(n6484) );
  AOI22D1BWP30P140LVT U9502 ( .A1(i_data_bus[357]), .A2(n10511), .B1(
        i_data_bus[293]), .B2(n10512), .ZN(n6483) );
  ND2D1BWP30P140LVT U9503 ( .A1(n6484), .A2(n6483), .ZN(N8504) );
  AOI22D1BWP30P140LVT U9504 ( .A1(i_data_bus[376]), .A2(n10511), .B1(
        i_data_bus[344]), .B2(n10509), .ZN(n6486) );
  AOI22D1BWP30P140LVT U9505 ( .A1(i_data_bus[280]), .A2(n10510), .B1(
        i_data_bus[312]), .B2(n10512), .ZN(n6485) );
  ND2D1BWP30P140LVT U9506 ( .A1(n6486), .A2(n6485), .ZN(N8523) );
  AOI22D1BWP30P140LVT U9507 ( .A1(i_data_bus[367]), .A2(n10511), .B1(
        i_data_bus[335]), .B2(n10509), .ZN(n6488) );
  AOI22D1BWP30P140LVT U9508 ( .A1(i_data_bus[271]), .A2(n10510), .B1(
        i_data_bus[303]), .B2(n10512), .ZN(n6487) );
  ND2D1BWP30P140LVT U9509 ( .A1(n6488), .A2(n6487), .ZN(N8514) );
  AOI22D1BWP30P140LVT U9510 ( .A1(i_data_bus[350]), .A2(n10509), .B1(
        i_data_bus[286]), .B2(n10510), .ZN(n6490) );
  AOI22D1BWP30P140LVT U9511 ( .A1(i_data_bus[382]), .A2(n10511), .B1(
        i_data_bus[318]), .B2(n10512), .ZN(n6489) );
  ND2D1BWP30P140LVT U9512 ( .A1(n6490), .A2(n6489), .ZN(N8529) );
  AOI22D1BWP30P140LVT U9513 ( .A1(i_data_bus[813]), .A2(n10592), .B1(
        i_data_bus[781]), .B2(n10589), .ZN(n6492) );
  AOI22D1BWP30P140LVT U9514 ( .A1(i_data_bus[845]), .A2(n10590), .B1(
        i_data_bus[877]), .B2(n10591), .ZN(n6491) );
  ND2D1BWP30P140LVT U9515 ( .A1(n6492), .A2(n6491), .ZN(N3754) );
  AOI22D1BWP30P140LVT U9516 ( .A1(i_data_bus[832]), .A2(n10590), .B1(
        i_data_bus[768]), .B2(n10589), .ZN(n6494) );
  AOI22D1BWP30P140LVT U9517 ( .A1(i_data_bus[800]), .A2(n10592), .B1(
        i_data_bus[864]), .B2(n10591), .ZN(n6493) );
  ND2D1BWP30P140LVT U9518 ( .A1(n6494), .A2(n6493), .ZN(N3741) );
  INR4D1BWP30P140LVT U9519 ( .A1(i_cmd[190]), .B1(i_cmd[174]), .B2(n9844), 
        .B3(n6495), .ZN(n10433) );
  INR4D1BWP30P140LVT U9520 ( .A1(i_cmd[174]), .B1(i_cmd[190]), .B2(n9847), 
        .B3(n6495), .ZN(n10436) );
  AOI22D1BWP30P140LVT U9521 ( .A1(i_data_bus[744]), .A2(n10433), .B1(
        i_data_bus[680]), .B2(n10436), .ZN(n6500) );
  NR4D1BWP30P140LVT U9522 ( .A1(i_cmd[182]), .A2(n6496), .A3(n9843), .A4(n6497), .ZN(n10435) );
  NR4D1BWP30P140LVT U9523 ( .A1(i_cmd[166]), .A2(n9850), .A3(n6498), .A4(n6497), .ZN(n10434) );
  AOI22D1BWP30P140LVT U9524 ( .A1(i_data_bus[648]), .A2(n10435), .B1(
        i_data_bus[712]), .B2(n10434), .ZN(n6499) );
  ND2D1BWP30P140LVT U9525 ( .A1(n6500), .A2(n6499), .ZN(N12903) );
  AOI22D1BWP30P140LVT U9526 ( .A1(i_data_bus[644]), .A2(n10435), .B1(
        i_data_bus[676]), .B2(n10436), .ZN(n6502) );
  AOI22D1BWP30P140LVT U9527 ( .A1(i_data_bus[740]), .A2(n10433), .B1(
        i_data_bus[708]), .B2(n10434), .ZN(n6501) );
  ND2D1BWP30P140LVT U9528 ( .A1(n6502), .A2(n6501), .ZN(N12899) );
  AOI22D1BWP30P140LVT U9529 ( .A1(i_data_bus[659]), .A2(n10435), .B1(
        i_data_bus[691]), .B2(n10436), .ZN(n6504) );
  AOI22D1BWP30P140LVT U9530 ( .A1(i_data_bus[755]), .A2(n10433), .B1(
        i_data_bus[723]), .B2(n10434), .ZN(n6503) );
  ND2D1BWP30P140LVT U9531 ( .A1(n6504), .A2(n6503), .ZN(N12914) );
  AOI22D1BWP30P140LVT U9532 ( .A1(i_data_bus[749]), .A2(n10433), .B1(
        i_data_bus[685]), .B2(n10436), .ZN(n6506) );
  AOI22D1BWP30P140LVT U9533 ( .A1(i_data_bus[653]), .A2(n10435), .B1(
        i_data_bus[717]), .B2(n10434), .ZN(n6505) );
  ND2D1BWP30P140LVT U9534 ( .A1(n6506), .A2(n6505), .ZN(N12908) );
  AOI22D1BWP30P140LVT U9535 ( .A1(i_data_bus[753]), .A2(n10433), .B1(
        i_data_bus[689]), .B2(n10436), .ZN(n6508) );
  AOI22D1BWP30P140LVT U9536 ( .A1(i_data_bus[657]), .A2(n10435), .B1(
        i_data_bus[721]), .B2(n10434), .ZN(n6507) );
  ND2D1BWP30P140LVT U9537 ( .A1(n6508), .A2(n6507), .ZN(N12912) );
  NR4D1BWP30P140LVT U9538 ( .A1(i_cmd[137]), .A2(n6509), .A3(n9837), .A4(n6511), .ZN(n10599) );
  INR4D1BWP30P140LVT U9539 ( .A1(i_cmd[145]), .B1(i_cmd[129]), .B2(n9834), 
        .B3(n6510), .ZN(n10600) );
  AOI22D1BWP30P140LVT U9540 ( .A1(i_data_bus[612]), .A2(n10599), .B1(
        i_data_bus[580]), .B2(n10600), .ZN(n6514) );
  INR4D1BWP30P140LVT U9541 ( .A1(i_cmd[129]), .B1(i_cmd[145]), .B2(n9839), 
        .B3(n6510), .ZN(n10597) );
  NR4D1BWP30P140LVT U9542 ( .A1(i_cmd[153]), .A2(n9833), .A3(n6512), .A4(n6511), .ZN(n10598) );
  AOI22D1BWP30P140LVT U9543 ( .A1(i_data_bus[516]), .A2(n10597), .B1(
        i_data_bus[548]), .B2(n10598), .ZN(n6513) );
  ND2D1BWP30P140LVT U9544 ( .A1(n6514), .A2(n6513), .ZN(N3313) );
  AOI22D1BWP30P140LVT U9545 ( .A1(i_data_bus[611]), .A2(n10599), .B1(
        i_data_bus[579]), .B2(n10600), .ZN(n6516) );
  AOI22D1BWP30P140LVT U9546 ( .A1(i_data_bus[515]), .A2(n10597), .B1(
        i_data_bus[547]), .B2(n10598), .ZN(n6515) );
  ND2D1BWP30P140LVT U9547 ( .A1(n6516), .A2(n6515), .ZN(N3312) );
  AOI22D1BWP30P140LVT U9548 ( .A1(i_data_bus[521]), .A2(n10597), .B1(
        i_data_bus[585]), .B2(n10600), .ZN(n6518) );
  AOI22D1BWP30P140LVT U9549 ( .A1(i_data_bus[617]), .A2(n10599), .B1(
        i_data_bus[553]), .B2(n10598), .ZN(n6517) );
  ND2D1BWP30P140LVT U9550 ( .A1(n6518), .A2(n6517), .ZN(N3318) );
  AOI22D1BWP30P140LVT U9551 ( .A1(i_data_bus[610]), .A2(n10599), .B1(
        i_data_bus[514]), .B2(n10597), .ZN(n6520) );
  AOI22D1BWP30P140LVT U9552 ( .A1(i_data_bus[578]), .A2(n10600), .B1(
        i_data_bus[546]), .B2(n10598), .ZN(n6519) );
  ND2D1BWP30P140LVT U9553 ( .A1(n6520), .A2(n6519), .ZN(N3311) );
  AOI22D1BWP30P140LVT U9554 ( .A1(i_data_bus[637]), .A2(n10599), .B1(
        i_data_bus[541]), .B2(n10597), .ZN(n6522) );
  AOI22D1BWP30P140LVT U9555 ( .A1(i_data_bus[605]), .A2(n10600), .B1(
        i_data_bus[573]), .B2(n10598), .ZN(n6521) );
  ND2D1BWP30P140LVT U9556 ( .A1(n6522), .A2(n6521), .ZN(N3338) );
  AOI22D1BWP30P140LVT U9557 ( .A1(i_data_bus[636]), .A2(n10599), .B1(
        i_data_bus[540]), .B2(n10597), .ZN(n6524) );
  AOI22D1BWP30P140LVT U9558 ( .A1(i_data_bus[604]), .A2(n10600), .B1(
        i_data_bus[572]), .B2(n10598), .ZN(n6523) );
  ND2D1BWP30P140LVT U9559 ( .A1(n6524), .A2(n6523), .ZN(N3337) );
  AOI22D1BWP30P140LVT U9560 ( .A1(i_data_bus[711]), .A2(n10465), .B1(
        i_data_bus[743]), .B2(n10466), .ZN(n6526) );
  AOI22D1BWP30P140LVT U9561 ( .A1(i_data_bus[679]), .A2(n10468), .B1(
        i_data_bus[647]), .B2(n10467), .ZN(n6525) );
  ND2D1BWP30P140LVT U9562 ( .A1(n6526), .A2(n6525), .ZN(N11028) );
  AOI22D1BWP30P140LVT U9563 ( .A1(i_data_bus[704]), .A2(n10465), .B1(
        i_data_bus[736]), .B2(n10466), .ZN(n6528) );
  AOI22D1BWP30P140LVT U9564 ( .A1(i_data_bus[672]), .A2(n10468), .B1(
        i_data_bus[640]), .B2(n10467), .ZN(n6527) );
  ND2D1BWP30P140LVT U9565 ( .A1(n6528), .A2(n6527), .ZN(N11021) );
  AOI22D1BWP30P140LVT U9566 ( .A1(i_data_bus[687]), .A2(n10468), .B1(
        i_data_bus[751]), .B2(n10466), .ZN(n6530) );
  AOI22D1BWP30P140LVT U9567 ( .A1(i_data_bus[719]), .A2(n10465), .B1(
        i_data_bus[655]), .B2(n10467), .ZN(n6529) );
  ND2D1BWP30P140LVT U9568 ( .A1(n6530), .A2(n6529), .ZN(N11036) );
  AOI22D1BWP30P140LVT U9569 ( .A1(i_data_bus[730]), .A2(n10465), .B1(
        i_data_bus[762]), .B2(n10466), .ZN(n6532) );
  AOI22D1BWP30P140LVT U9570 ( .A1(i_data_bus[698]), .A2(n10468), .B1(
        i_data_bus[666]), .B2(n10467), .ZN(n6531) );
  ND2D1BWP30P140LVT U9571 ( .A1(n6532), .A2(n6531), .ZN(N11047) );
  AOI22D1BWP30P140LVT U9572 ( .A1(i_data_bus[720]), .A2(n10465), .B1(
        i_data_bus[688]), .B2(n10468), .ZN(n6534) );
  AOI22D1BWP30P140LVT U9573 ( .A1(i_data_bus[752]), .A2(n10466), .B1(
        i_data_bus[656]), .B2(n10467), .ZN(n6533) );
  ND2D1BWP30P140LVT U9574 ( .A1(n6534), .A2(n6533), .ZN(N11037) );
  AOI22D1BWP30P140LVT U9575 ( .A1(i_data_bus[454]), .A2(n10538), .B1(
        i_data_bus[390]), .B2(n10537), .ZN(n6536) );
  AOI22D1BWP30P140LVT U9576 ( .A1(i_data_bus[422]), .A2(n10540), .B1(
        i_data_bus[486]), .B2(n10539), .ZN(n6535) );
  ND2D1BWP30P140LVT U9577 ( .A1(n6536), .A2(n6535), .ZN(N6847) );
  NR4D1BWP30P140LVT U9578 ( .A1(i_cmd[236]), .A2(n6537), .A3(n10030), .A4(
        n6539), .ZN(n10489) );
  INR4D1BWP30P140LVT U9579 ( .A1(i_cmd[228]), .B1(i_cmd[244]), .B2(n10028), 
        .B3(n6538), .ZN(n10492) );
  AOI22D1BWP30P140LVT U9580 ( .A1(i_data_bus[1001]), .A2(n10489), .B1(
        i_data_bus[905]), .B2(n10492), .ZN(n6542) );
  INR4D1BWP30P140LVT U9581 ( .A1(i_cmd[244]), .B1(i_cmd[228]), .B2(n10024), 
        .B3(n6538), .ZN(n10490) );
  NR4D1BWP30P140LVT U9582 ( .A1(i_cmd[252]), .A2(n10023), .A3(n6540), .A4(
        n6539), .ZN(n10491) );
  AOI22D1BWP30P140LVT U9583 ( .A1(i_data_bus[969]), .A2(n10490), .B1(
        i_data_bus[937]), .B2(n10491), .ZN(n6541) );
  ND2D1BWP30P140LVT U9584 ( .A1(n6542), .A2(n6541), .ZN(N9588) );
  AOI22D1BWP30P140LVT U9585 ( .A1(i_data_bus[981]), .A2(n10490), .B1(
        i_data_bus[917]), .B2(n10492), .ZN(n6544) );
  AOI22D1BWP30P140LVT U9586 ( .A1(i_data_bus[1013]), .A2(n10489), .B1(
        i_data_bus[949]), .B2(n10491), .ZN(n6543) );
  ND2D1BWP30P140LVT U9587 ( .A1(n6544), .A2(n6543), .ZN(N9600) );
  AOI22D1BWP30P140LVT U9588 ( .A1(i_data_bus[980]), .A2(n10490), .B1(
        i_data_bus[916]), .B2(n10492), .ZN(n6546) );
  AOI22D1BWP30P140LVT U9589 ( .A1(i_data_bus[1012]), .A2(n10489), .B1(
        i_data_bus[948]), .B2(n10491), .ZN(n6545) );
  ND2D1BWP30P140LVT U9590 ( .A1(n6546), .A2(n6545), .ZN(N9599) );
  AOI22D1BWP30P140LVT U9591 ( .A1(i_data_bus[988]), .A2(n10490), .B1(
        i_data_bus[924]), .B2(n10492), .ZN(n6548) );
  AOI22D1BWP30P140LVT U9592 ( .A1(i_data_bus[1020]), .A2(n10489), .B1(
        i_data_bus[956]), .B2(n10491), .ZN(n6547) );
  ND2D1BWP30P140LVT U9593 ( .A1(n6548), .A2(n6547), .ZN(N9607) );
  AOI22D1BWP30P140LVT U9594 ( .A1(i_data_bus[769]), .A2(n10397), .B1(
        i_data_bus[833]), .B2(n10399), .ZN(n6550) );
  AOI22D1BWP30P140LVT U9595 ( .A1(i_data_bus[801]), .A2(n10400), .B1(
        i_data_bus[865]), .B2(n10398), .ZN(n6549) );
  ND2D1BWP30P140LVT U9596 ( .A1(n6550), .A2(n6549), .ZN(N14986) );
  AOI22D1BWP30P140LVT U9597 ( .A1(i_data_bus[790]), .A2(n10397), .B1(
        i_data_bus[854]), .B2(n10399), .ZN(n6552) );
  AOI22D1BWP30P140LVT U9598 ( .A1(i_data_bus[822]), .A2(n10400), .B1(
        i_data_bus[886]), .B2(n10398), .ZN(n6551) );
  ND2D1BWP30P140LVT U9599 ( .A1(n6552), .A2(n6551), .ZN(N15007) );
  AOI22D1BWP30P140LVT U9600 ( .A1(i_data_bus[860]), .A2(n10495), .B1(
        i_data_bus[796]), .B2(n10493), .ZN(n6554) );
  AOI22D1BWP30P140LVT U9601 ( .A1(i_data_bus[828]), .A2(n10496), .B1(
        i_data_bus[892]), .B2(n10494), .ZN(n6553) );
  ND2D1BWP30P140LVT U9602 ( .A1(n6554), .A2(n6553), .ZN(N9391) );
  AOI22D1BWP30P140LVT U9603 ( .A1(i_data_bus[471]), .A2(n10410), .B1(
        i_data_bus[439]), .B2(n10411), .ZN(n6556) );
  AOI22D1BWP30P140LVT U9604 ( .A1(i_data_bus[503]), .A2(n10412), .B1(
        i_data_bus[407]), .B2(n10409), .ZN(n6555) );
  ND2D1BWP30P140LVT U9605 ( .A1(n6556), .A2(n6555), .ZN(N14360) );
  AOI22D1BWP30P140LVT U9606 ( .A1(i_data_bus[499]), .A2(n10412), .B1(
        i_data_bus[435]), .B2(n10411), .ZN(n6558) );
  AOI22D1BWP30P140LVT U9607 ( .A1(i_data_bus[467]), .A2(n10410), .B1(
        i_data_bus[403]), .B2(n10409), .ZN(n6557) );
  ND2D1BWP30P140LVT U9608 ( .A1(n6558), .A2(n6557), .ZN(N14356) );
  AOI22D1BWP30P140LVT U9609 ( .A1(i_data_bus[460]), .A2(n10410), .B1(
        i_data_bus[428]), .B2(n10411), .ZN(n6560) );
  AOI22D1BWP30P140LVT U9610 ( .A1(i_data_bus[492]), .A2(n10412), .B1(
        i_data_bus[396]), .B2(n10409), .ZN(n6559) );
  ND2D1BWP30P140LVT U9611 ( .A1(n6560), .A2(n6559), .ZN(N14349) );
  AOI22D1BWP30P140LVT U9612 ( .A1(i_data_bus[404]), .A2(n10603), .B1(
        i_data_bus[468]), .B2(n10604), .ZN(n6562) );
  AOI22D1BWP30P140LVT U9613 ( .A1(i_data_bus[436]), .A2(n10601), .B1(
        i_data_bus[500]), .B2(n10602), .ZN(n6561) );
  ND2D1BWP30P140LVT U9614 ( .A1(n6562), .A2(n6561), .ZN(N3113) );
  AOI22D1BWP30P140LVT U9615 ( .A1(i_data_bus[408]), .A2(n10603), .B1(
        i_data_bus[472]), .B2(n10604), .ZN(n6564) );
  AOI22D1BWP30P140LVT U9616 ( .A1(i_data_bus[440]), .A2(n10601), .B1(
        i_data_bus[504]), .B2(n10602), .ZN(n6563) );
  ND2D1BWP30P140LVT U9617 ( .A1(n6564), .A2(n6563), .ZN(N3117) );
  AOI22D1BWP30P140LVT U9618 ( .A1(i_data_bus[433]), .A2(n10601), .B1(
        i_data_bus[465]), .B2(n10604), .ZN(n6566) );
  AOI22D1BWP30P140LVT U9619 ( .A1(i_data_bus[401]), .A2(n10603), .B1(
        i_data_bus[497]), .B2(n10602), .ZN(n6565) );
  ND2D1BWP30P140LVT U9620 ( .A1(n6566), .A2(n6565), .ZN(N3110) );
  AOI22D1BWP30P140LVT U9621 ( .A1(i_data_bus[388]), .A2(n10603), .B1(
        i_data_bus[452]), .B2(n10604), .ZN(n6568) );
  AOI22D1BWP30P140LVT U9622 ( .A1(i_data_bus[420]), .A2(n10601), .B1(
        i_data_bus[484]), .B2(n10602), .ZN(n6567) );
  ND2D1BWP30P140LVT U9623 ( .A1(n6568), .A2(n6567), .ZN(N3097) );
  AOI22D1BWP30P140LVT U9624 ( .A1(i_data_bus[411]), .A2(n10603), .B1(
        i_data_bus[475]), .B2(n10604), .ZN(n6570) );
  AOI22D1BWP30P140LVT U9625 ( .A1(i_data_bus[443]), .A2(n10601), .B1(
        i_data_bus[507]), .B2(n10602), .ZN(n6569) );
  ND2D1BWP30P140LVT U9626 ( .A1(n6570), .A2(n6569), .ZN(N3120) );
  AOI22D1BWP30P140LVT U9627 ( .A1(i_data_bus[399]), .A2(n10603), .B1(
        i_data_bus[463]), .B2(n10604), .ZN(n6572) );
  AOI22D1BWP30P140LVT U9628 ( .A1(i_data_bus[431]), .A2(n10601), .B1(
        i_data_bus[495]), .B2(n10602), .ZN(n6571) );
  ND2D1BWP30P140LVT U9629 ( .A1(n6572), .A2(n6571), .ZN(N3108) );
  AOI22D1BWP30P140LVT U9630 ( .A1(i_data_bus[394]), .A2(n10409), .B1(
        i_data_bus[426]), .B2(n10411), .ZN(n6574) );
  AOI22D1BWP30P140LVT U9631 ( .A1(i_data_bus[458]), .A2(n10410), .B1(
        i_data_bus[490]), .B2(n10412), .ZN(n6573) );
  ND2D1BWP30P140LVT U9632 ( .A1(n6574), .A2(n6573), .ZN(N14347) );
  AOI22D1BWP30P140LVT U9633 ( .A1(i_data_bus[408]), .A2(n10409), .B1(
        i_data_bus[440]), .B2(n10411), .ZN(n6576) );
  AOI22D1BWP30P140LVT U9634 ( .A1(i_data_bus[472]), .A2(n10410), .B1(
        i_data_bus[504]), .B2(n10412), .ZN(n6575) );
  ND2D1BWP30P140LVT U9635 ( .A1(n6576), .A2(n6575), .ZN(N14361) );
  AOI22D1BWP30P140LVT U9636 ( .A1(i_data_bus[391]), .A2(n10409), .B1(
        i_data_bus[423]), .B2(n10411), .ZN(n6578) );
  AOI22D1BWP30P140LVT U9637 ( .A1(i_data_bus[455]), .A2(n10410), .B1(
        i_data_bus[487]), .B2(n10412), .ZN(n6577) );
  ND2D1BWP30P140LVT U9638 ( .A1(n6578), .A2(n6577), .ZN(N14344) );
  AOI22D1BWP30P140LVT U9639 ( .A1(i_data_bus[452]), .A2(n10410), .B1(
        i_data_bus[420]), .B2(n10411), .ZN(n6580) );
  AOI22D1BWP30P140LVT U9640 ( .A1(i_data_bus[388]), .A2(n10409), .B1(
        i_data_bus[484]), .B2(n10412), .ZN(n6579) );
  ND2D1BWP30P140LVT U9641 ( .A1(n6580), .A2(n6579), .ZN(N14341) );
  INR4D1BWP30P140LVT U9642 ( .A1(i_cmd[26]), .B1(i_cmd[10]), .B2(n10019), .B3(
        n6581), .ZN(n10584) );
  INR4D1BWP30P140LVT U9643 ( .A1(i_cmd[10]), .B1(i_cmd[26]), .B2(n10018), .B3(
        n6581), .ZN(n10583) );
  AOI22D1BWP30P140LVT U9644 ( .A1(i_data_bus[117]), .A2(n10584), .B1(
        i_data_bus[53]), .B2(n10583), .ZN(n6586) );
  NR4D1BWP30P140LVT U9645 ( .A1(i_cmd[18]), .A2(n6582), .A3(n10013), .A4(n6583), .ZN(n10581) );
  NR4D1BWP30P140LVT U9646 ( .A1(i_cmd[2]), .A2(n10014), .A3(n6584), .A4(n6583), 
        .ZN(n10582) );
  AOI22D1BWP30P140LVT U9647 ( .A1(i_data_bus[21]), .A2(n10581), .B1(
        i_data_bus[85]), .B2(n10582), .ZN(n6585) );
  ND2D1BWP30P140LVT U9648 ( .A1(n6586), .A2(n6585), .ZN(N4340) );
  AOI22D1BWP30P140LVT U9649 ( .A1(i_data_bus[14]), .A2(n10581), .B1(
        i_data_bus[46]), .B2(n10583), .ZN(n6588) );
  AOI22D1BWP30P140LVT U9650 ( .A1(i_data_bus[110]), .A2(n10584), .B1(
        i_data_bus[78]), .B2(n10582), .ZN(n6587) );
  ND2D1BWP30P140LVT U9651 ( .A1(n6588), .A2(n6587), .ZN(N4333) );
  AOI22D1BWP30P140LVT U9652 ( .A1(i_data_bus[15]), .A2(n10581), .B1(
        i_data_bus[47]), .B2(n10583), .ZN(n6590) );
  AOI22D1BWP30P140LVT U9653 ( .A1(i_data_bus[111]), .A2(n10584), .B1(
        i_data_bus[79]), .B2(n10582), .ZN(n6589) );
  ND2D1BWP30P140LVT U9654 ( .A1(n6590), .A2(n6589), .ZN(N4334) );
  AOI22D1BWP30P140LVT U9655 ( .A1(i_data_bus[120]), .A2(n10584), .B1(
        i_data_bus[56]), .B2(n10583), .ZN(n6592) );
  AOI22D1BWP30P140LVT U9656 ( .A1(i_data_bus[24]), .A2(n10581), .B1(
        i_data_bus[88]), .B2(n10582), .ZN(n6591) );
  ND2D1BWP30P140LVT U9657 ( .A1(n6592), .A2(n6591), .ZN(N4343) );
  AOI22D1BWP30P140LVT U9658 ( .A1(i_data_bus[29]), .A2(n10581), .B1(
        i_data_bus[125]), .B2(n10584), .ZN(n6594) );
  AOI22D1BWP30P140LVT U9659 ( .A1(i_data_bus[61]), .A2(n10583), .B1(
        i_data_bus[93]), .B2(n10582), .ZN(n6593) );
  ND2D1BWP30P140LVT U9660 ( .A1(n6594), .A2(n6593), .ZN(N4348) );
  AOI22D1BWP30P140LVT U9661 ( .A1(i_data_bus[756]), .A2(n10466), .B1(
        i_data_bus[724]), .B2(n10465), .ZN(n6596) );
  AOI22D1BWP30P140LVT U9662 ( .A1(i_data_bus[692]), .A2(n10468), .B1(
        i_data_bus[660]), .B2(n10467), .ZN(n6595) );
  ND2D1BWP30P140LVT U9663 ( .A1(n6596), .A2(n6595), .ZN(N11041) );
  AOI22D1BWP30P140LVT U9664 ( .A1(i_data_bus[737]), .A2(n10466), .B1(
        i_data_bus[705]), .B2(n10465), .ZN(n6598) );
  AOI22D1BWP30P140LVT U9665 ( .A1(i_data_bus[673]), .A2(n10468), .B1(
        i_data_bus[641]), .B2(n10467), .ZN(n6597) );
  ND2D1BWP30P140LVT U9666 ( .A1(n6598), .A2(n6597), .ZN(N11022) );
  AOI22D1BWP30P140LVT U9667 ( .A1(i_data_bus[758]), .A2(n10466), .B1(
        i_data_bus[726]), .B2(n10465), .ZN(n6600) );
  AOI22D1BWP30P140LVT U9668 ( .A1(i_data_bus[694]), .A2(n10468), .B1(
        i_data_bus[662]), .B2(n10467), .ZN(n6599) );
  ND2D1BWP30P140LVT U9669 ( .A1(n6600), .A2(n6599), .ZN(N11043) );
  AOI22D1BWP30P140LVT U9670 ( .A1(i_data_bus[648]), .A2(n10467), .B1(
        i_data_bus[712]), .B2(n10465), .ZN(n6602) );
  AOI22D1BWP30P140LVT U9671 ( .A1(i_data_bus[744]), .A2(n10466), .B1(
        i_data_bus[680]), .B2(n10468), .ZN(n6601) );
  ND2D1BWP30P140LVT U9672 ( .A1(n6602), .A2(n6601), .ZN(N11029) );
  AOI22D1BWP30P140LVT U9673 ( .A1(i_data_bus[691]), .A2(n10468), .B1(
        i_data_bus[723]), .B2(n10465), .ZN(n6604) );
  AOI22D1BWP30P140LVT U9674 ( .A1(i_data_bus[659]), .A2(n10467), .B1(
        i_data_bus[755]), .B2(n10466), .ZN(n6603) );
  ND2D1BWP30P140LVT U9675 ( .A1(n6604), .A2(n6603), .ZN(N11040) );
  AOI22D1BWP30P140LVT U9676 ( .A1(i_data_bus[753]), .A2(n10466), .B1(
        i_data_bus[721]), .B2(n10465), .ZN(n6606) );
  AOI22D1BWP30P140LVT U9677 ( .A1(i_data_bus[657]), .A2(n10467), .B1(
        i_data_bus[689]), .B2(n10468), .ZN(n6605) );
  ND2D1BWP30P140LVT U9678 ( .A1(n6606), .A2(n6605), .ZN(N11038) );
  AOI22D1BWP30P140LVT U9679 ( .A1(i_data_bus[695]), .A2(n10468), .B1(
        i_data_bus[727]), .B2(n10465), .ZN(n6608) );
  AOI22D1BWP30P140LVT U9680 ( .A1(i_data_bus[663]), .A2(n10467), .B1(
        i_data_bus[759]), .B2(n10466), .ZN(n6607) );
  ND2D1BWP30P140LVT U9681 ( .A1(n6608), .A2(n6607), .ZN(N11044) );
  AOI22D1BWP30P140LVT U9682 ( .A1(i_data_bus[513]), .A2(n10405), .B1(
        i_data_bus[577]), .B2(n10408), .ZN(n6610) );
  AOI22D1BWP30P140LVT U9683 ( .A1(i_data_bus[609]), .A2(n10407), .B1(
        i_data_bus[545]), .B2(n10406), .ZN(n6609) );
  ND2D1BWP30P140LVT U9684 ( .A1(n6610), .A2(n6609), .ZN(N14554) );
  AOI22D1BWP30P140LVT U9685 ( .A1(i_data_bus[613]), .A2(n10407), .B1(
        i_data_bus[581]), .B2(n10408), .ZN(n6612) );
  AOI22D1BWP30P140LVT U9686 ( .A1(i_data_bus[517]), .A2(n10405), .B1(
        i_data_bus[549]), .B2(n10406), .ZN(n6611) );
  ND2D1BWP30P140LVT U9687 ( .A1(n6612), .A2(n6611), .ZN(N14558) );
  AOI22D1BWP30P140LVT U9688 ( .A1(i_data_bus[631]), .A2(n10407), .B1(
        i_data_bus[535]), .B2(n10405), .ZN(n6614) );
  AOI22D1BWP30P140LVT U9689 ( .A1(i_data_bus[599]), .A2(n10408), .B1(
        i_data_bus[567]), .B2(n10406), .ZN(n6613) );
  ND2D1BWP30P140LVT U9690 ( .A1(n6614), .A2(n6613), .ZN(N14576) );
  AOI22D1BWP30P140LVT U9691 ( .A1(i_data_bus[636]), .A2(n10407), .B1(
        i_data_bus[540]), .B2(n10405), .ZN(n6616) );
  AOI22D1BWP30P140LVT U9692 ( .A1(i_data_bus[604]), .A2(n10408), .B1(
        i_data_bus[572]), .B2(n10406), .ZN(n6615) );
  ND2D1BWP30P140LVT U9693 ( .A1(n6616), .A2(n6615), .ZN(N14581) );
  AOI22D1BWP30P140LVT U9694 ( .A1(i_data_bus[637]), .A2(n10407), .B1(
        i_data_bus[541]), .B2(n10405), .ZN(n6618) );
  AOI22D1BWP30P140LVT U9695 ( .A1(i_data_bus[605]), .A2(n10408), .B1(
        i_data_bus[573]), .B2(n10406), .ZN(n6617) );
  ND2D1BWP30P140LVT U9696 ( .A1(n6618), .A2(n6617), .ZN(N14582) );
  NR4D1BWP30P140LVT U9697 ( .A1(i_cmd[9]), .A2(n6619), .A3(n10019), .A4(n6621), 
        .ZN(n10616) );
  INR4D1BWP30P140LVT U9698 ( .A1(i_cmd[17]), .B1(i_cmd[1]), .B2(n10014), .B3(
        n6620), .ZN(n10613) );
  AOI22D1BWP30P140LVT U9699 ( .A1(i_data_bus[117]), .A2(n10616), .B1(
        i_data_bus[85]), .B2(n10613), .ZN(n6624) );
  INR4D1BWP30P140LVT U9700 ( .A1(i_cmd[1]), .B1(i_cmd[17]), .B2(n10013), .B3(
        n6620), .ZN(n10615) );
  NR4D1BWP30P140LVT U9701 ( .A1(i_cmd[25]), .A2(n10018), .A3(n6622), .A4(n6621), .ZN(n10614) );
  AOI22D1BWP30P140LVT U9702 ( .A1(i_data_bus[21]), .A2(n10615), .B1(
        i_data_bus[53]), .B2(n10614), .ZN(n6623) );
  ND2D1BWP30P140LVT U9703 ( .A1(n6624), .A2(n6623), .ZN(N2466) );
  AOI22D1BWP30P140LVT U9704 ( .A1(i_data_bus[110]), .A2(n10616), .B1(
        i_data_bus[78]), .B2(n10613), .ZN(n6626) );
  AOI22D1BWP30P140LVT U9705 ( .A1(i_data_bus[14]), .A2(n10615), .B1(
        i_data_bus[46]), .B2(n10614), .ZN(n6625) );
  ND2D1BWP30P140LVT U9706 ( .A1(n6626), .A2(n6625), .ZN(N2459) );
  AOI22D1BWP30P140LVT U9707 ( .A1(i_data_bus[73]), .A2(n10613), .B1(
        i_data_bus[105]), .B2(n10616), .ZN(n6628) );
  AOI22D1BWP30P140LVT U9708 ( .A1(i_data_bus[9]), .A2(n10615), .B1(
        i_data_bus[41]), .B2(n10614), .ZN(n6627) );
  ND2D1BWP30P140LVT U9709 ( .A1(n6628), .A2(n6627), .ZN(N2454) );
  AOI22D1BWP30P140LVT U9710 ( .A1(i_data_bus[673]), .A2(n10436), .B1(
        i_data_bus[737]), .B2(n10433), .ZN(n6630) );
  AOI22D1BWP30P140LVT U9711 ( .A1(i_data_bus[641]), .A2(n10435), .B1(
        i_data_bus[705]), .B2(n10434), .ZN(n6629) );
  ND2D1BWP30P140LVT U9712 ( .A1(n6630), .A2(n6629), .ZN(N12896) );
  AOI22D1BWP30P140LVT U9713 ( .A1(i_data_bus[667]), .A2(n10435), .B1(
        i_data_bus[763]), .B2(n10433), .ZN(n6632) );
  AOI22D1BWP30P140LVT U9714 ( .A1(i_data_bus[699]), .A2(n10436), .B1(
        i_data_bus[731]), .B2(n10434), .ZN(n6631) );
  ND2D1BWP30P140LVT U9715 ( .A1(n6632), .A2(n6631), .ZN(N12922) );
  AOI22D1BWP30P140LVT U9716 ( .A1(i_data_bus[663]), .A2(n10435), .B1(
        i_data_bus[759]), .B2(n10433), .ZN(n6634) );
  AOI22D1BWP30P140LVT U9717 ( .A1(i_data_bus[695]), .A2(n10436), .B1(
        i_data_bus[727]), .B2(n10434), .ZN(n6633) );
  ND2D1BWP30P140LVT U9718 ( .A1(n6634), .A2(n6633), .ZN(N12918) );
  AOI22D1BWP30P140LVT U9719 ( .A1(i_data_bus[482]), .A2(n10539), .B1(
        i_data_bus[386]), .B2(n10537), .ZN(n6636) );
  AOI22D1BWP30P140LVT U9720 ( .A1(i_data_bus[418]), .A2(n10540), .B1(
        i_data_bus[450]), .B2(n10538), .ZN(n6635) );
  ND2D1BWP30P140LVT U9721 ( .A1(n6636), .A2(n6635), .ZN(N6843) );
  AOI22D1BWP30P140LVT U9722 ( .A1(i_data_bus[508]), .A2(n10539), .B1(
        i_data_bus[412]), .B2(n10537), .ZN(n6638) );
  AOI22D1BWP30P140LVT U9723 ( .A1(i_data_bus[444]), .A2(n10540), .B1(
        i_data_bus[476]), .B2(n10538), .ZN(n6637) );
  ND2D1BWP30P140LVT U9724 ( .A1(n6638), .A2(n6637), .ZN(N6869) );
  AOI22D1BWP30P140LVT U9725 ( .A1(i_data_bus[433]), .A2(n10540), .B1(
        i_data_bus[497]), .B2(n10539), .ZN(n6640) );
  AOI22D1BWP30P140LVT U9726 ( .A1(i_data_bus[401]), .A2(n10537), .B1(
        i_data_bus[465]), .B2(n10538), .ZN(n6639) );
  ND2D1BWP30P140LVT U9727 ( .A1(n6640), .A2(n6639), .ZN(N6858) );
  AOI22D1BWP30P140LVT U9728 ( .A1(i_data_bus[427]), .A2(n10540), .B1(
        i_data_bus[395]), .B2(n10537), .ZN(n6642) );
  AOI22D1BWP30P140LVT U9729 ( .A1(i_data_bus[491]), .A2(n10539), .B1(
        i_data_bus[459]), .B2(n10538), .ZN(n6641) );
  ND2D1BWP30P140LVT U9730 ( .A1(n6642), .A2(n6641), .ZN(N6852) );
  AOI22D1BWP30P140LVT U9731 ( .A1(i_data_bus[507]), .A2(n10539), .B1(
        i_data_bus[411]), .B2(n10537), .ZN(n6644) );
  AOI22D1BWP30P140LVT U9732 ( .A1(i_data_bus[443]), .A2(n10540), .B1(
        i_data_bus[475]), .B2(n10538), .ZN(n6643) );
  ND2D1BWP30P140LVT U9733 ( .A1(n6644), .A2(n6643), .ZN(N6868) );
  AOI22D1BWP30P140LVT U9734 ( .A1(i_data_bus[431]), .A2(n10540), .B1(
        i_data_bus[399]), .B2(n10537), .ZN(n6646) );
  AOI22D1BWP30P140LVT U9735 ( .A1(i_data_bus[495]), .A2(n10539), .B1(
        i_data_bus[463]), .B2(n10538), .ZN(n6645) );
  ND2D1BWP30P140LVT U9736 ( .A1(n6646), .A2(n6645), .ZN(N6856) );
  INR4D1BWP30P140LVT U9737 ( .A1(i_cmd[22]), .B1(i_cmd[6]), .B2(n10014), .B3(
        n6648), .ZN(n10454) );
  NR4D1BWP30P140LVT U9738 ( .A1(i_cmd[30]), .A2(n6647), .A3(n10018), .A4(n6649), .ZN(n10453) );
  AOI22D1BWP30P140LVT U9739 ( .A1(i_data_bus[87]), .A2(n10454), .B1(
        i_data_bus[55]), .B2(n10453), .ZN(n6652) );
  INR4D1BWP30P140LVT U9740 ( .A1(i_cmd[6]), .B1(i_cmd[22]), .B2(n10013), .B3(
        n6648), .ZN(n10456) );
  NR4D1BWP30P140LVT U9741 ( .A1(i_cmd[14]), .A2(n10019), .A3(n6650), .A4(n6649), .ZN(n10455) );
  AOI22D1BWP30P140LVT U9742 ( .A1(i_data_bus[23]), .A2(n10456), .B1(
        i_data_bus[119]), .B2(n10455), .ZN(n6651) );
  ND2D1BWP30P140LVT U9743 ( .A1(n6652), .A2(n6651), .ZN(N11838) );
  INR4D1BWP30P140LVT U9744 ( .A1(i_cmd[239]), .B1(i_cmd[255]), .B2(n10023), 
        .B3(n6653), .ZN(n10394) );
  INR4D1BWP30P140LVT U9745 ( .A1(i_cmd[255]), .B1(i_cmd[239]), .B2(n10030), 
        .B3(n6653), .ZN(n10393) );
  AOI22D1BWP30P140LVT U9746 ( .A1(i_data_bus[939]), .A2(n10394), .B1(
        i_data_bus[1003]), .B2(n10393), .ZN(n6658) );
  NR4D1BWP30P140LVT U9747 ( .A1(i_cmd[231]), .A2(n6654), .A3(n10024), .A4(
        n6655), .ZN(n10396) );
  NR4D1BWP30P140LVT U9748 ( .A1(i_cmd[247]), .A2(n10028), .A3(n6656), .A4(
        n6655), .ZN(n10395) );
  AOI22D1BWP30P140LVT U9749 ( .A1(i_data_bus[971]), .A2(n10396), .B1(
        i_data_bus[907]), .B2(n10395), .ZN(n6657) );
  ND2D1BWP30P140LVT U9750 ( .A1(n6658), .A2(n6657), .ZN(N15212) );
  AOI22D1BWP30P140LVT U9751 ( .A1(i_data_bus[986]), .A2(n10396), .B1(
        i_data_bus[1018]), .B2(n10393), .ZN(n6660) );
  AOI22D1BWP30P140LVT U9752 ( .A1(i_data_bus[954]), .A2(n10394), .B1(
        i_data_bus[922]), .B2(n10395), .ZN(n6659) );
  ND2D1BWP30P140LVT U9753 ( .A1(n6660), .A2(n6659), .ZN(N15227) );
  AOI22D1BWP30P140LVT U9754 ( .A1(i_data_bus[978]), .A2(n10396), .B1(
        i_data_bus[1010]), .B2(n10393), .ZN(n6662) );
  AOI22D1BWP30P140LVT U9755 ( .A1(i_data_bus[946]), .A2(n10394), .B1(
        i_data_bus[914]), .B2(n10395), .ZN(n6661) );
  ND2D1BWP30P140LVT U9756 ( .A1(n6662), .A2(n6661), .ZN(N15219) );
  AOI22D1BWP30P140LVT U9757 ( .A1(i_data_bus[953]), .A2(n10394), .B1(
        i_data_bus[1017]), .B2(n10393), .ZN(n6664) );
  AOI22D1BWP30P140LVT U9758 ( .A1(i_data_bus[985]), .A2(n10396), .B1(
        i_data_bus[921]), .B2(n10395), .ZN(n6663) );
  ND2D1BWP30P140LVT U9759 ( .A1(n6664), .A2(n6663), .ZN(N15226) );
  AOI22D1BWP30P140LVT U9760 ( .A1(i_data_bus[1013]), .A2(n10393), .B1(
        i_data_bus[949]), .B2(n10394), .ZN(n6666) );
  AOI22D1BWP30P140LVT U9761 ( .A1(i_data_bus[981]), .A2(n10396), .B1(
        i_data_bus[917]), .B2(n10395), .ZN(n6665) );
  ND2D1BWP30P140LVT U9762 ( .A1(n6666), .A2(n6665), .ZN(N15222) );
  AOI22D1BWP30P140LVT U9763 ( .A1(i_data_bus[980]), .A2(n10396), .B1(
        i_data_bus[948]), .B2(n10394), .ZN(n6668) );
  AOI22D1BWP30P140LVT U9764 ( .A1(i_data_bus[1012]), .A2(n10393), .B1(
        i_data_bus[916]), .B2(n10395), .ZN(n6667) );
  ND2D1BWP30P140LVT U9765 ( .A1(n6668), .A2(n6667), .ZN(N15221) );
  AOI22D1BWP30P140LVT U9766 ( .A1(i_data_bus[795]), .A2(n10462), .B1(
        i_data_bus[859]), .B2(n10463), .ZN(n6670) );
  AOI22D1BWP30P140LVT U9767 ( .A1(i_data_bus[827]), .A2(n10464), .B1(
        i_data_bus[891]), .B2(n10461), .ZN(n6669) );
  ND2D1BWP30P140LVT U9768 ( .A1(n6670), .A2(n6669), .ZN(N11264) );
  AOI22D1BWP30P140LVT U9769 ( .A1(i_data_bus[813]), .A2(n10464), .B1(
        i_data_bus[845]), .B2(n10463), .ZN(n6672) );
  AOI22D1BWP30P140LVT U9770 ( .A1(i_data_bus[781]), .A2(n10462), .B1(
        i_data_bus[877]), .B2(n10461), .ZN(n6671) );
  ND2D1BWP30P140LVT U9771 ( .A1(n6672), .A2(n6671), .ZN(N11250) );
  AOI22D1BWP30P140LVT U9772 ( .A1(i_data_bus[812]), .A2(n10464), .B1(
        i_data_bus[844]), .B2(n10463), .ZN(n6674) );
  AOI22D1BWP30P140LVT U9773 ( .A1(i_data_bus[780]), .A2(n10462), .B1(
        i_data_bus[876]), .B2(n10461), .ZN(n6673) );
  ND2D1BWP30P140LVT U9774 ( .A1(n6674), .A2(n6673), .ZN(N11249) );
  AOI22D1BWP30P140LVT U9775 ( .A1(i_data_bus[790]), .A2(n10462), .B1(
        i_data_bus[854]), .B2(n10463), .ZN(n6676) );
  AOI22D1BWP30P140LVT U9776 ( .A1(i_data_bus[822]), .A2(n10464), .B1(
        i_data_bus[886]), .B2(n10461), .ZN(n6675) );
  ND2D1BWP30P140LVT U9777 ( .A1(n6676), .A2(n6675), .ZN(N11259) );
  AOI22D1BWP30P140LVT U9778 ( .A1(i_data_bus[451]), .A2(n10508), .B1(
        i_data_bus[483]), .B2(n10506), .ZN(n6678) );
  AOI22D1BWP30P140LVT U9779 ( .A1(i_data_bus[387]), .A2(n10505), .B1(
        i_data_bus[419]), .B2(n10507), .ZN(n6677) );
  ND2D1BWP30P140LVT U9780 ( .A1(n6678), .A2(n6677), .ZN(N8718) );
  AOI22D1BWP30P140LVT U9781 ( .A1(i_data_bus[460]), .A2(n10508), .B1(
        i_data_bus[396]), .B2(n10505), .ZN(n6680) );
  AOI22D1BWP30P140LVT U9782 ( .A1(i_data_bus[492]), .A2(n10506), .B1(
        i_data_bus[428]), .B2(n10507), .ZN(n6679) );
  ND2D1BWP30P140LVT U9783 ( .A1(n6680), .A2(n6679), .ZN(N8727) );
  AOI22D1BWP30P140LVT U9784 ( .A1(i_data_bus[408]), .A2(n10505), .B1(
        i_data_bus[504]), .B2(n10506), .ZN(n6682) );
  AOI22D1BWP30P140LVT U9785 ( .A1(i_data_bus[472]), .A2(n10508), .B1(
        i_data_bus[440]), .B2(n10507), .ZN(n6681) );
  ND2D1BWP30P140LVT U9786 ( .A1(n6682), .A2(n6681), .ZN(N8739) );
  AOI22D1BWP30P140LVT U9787 ( .A1(i_data_bus[468]), .A2(n10508), .B1(
        i_data_bus[500]), .B2(n10506), .ZN(n6684) );
  AOI22D1BWP30P140LVT U9788 ( .A1(i_data_bus[404]), .A2(n10505), .B1(
        i_data_bus[436]), .B2(n10507), .ZN(n6683) );
  ND2D1BWP30P140LVT U9789 ( .A1(n6684), .A2(n6683), .ZN(N8735) );
  AOI22D1BWP30P140LVT U9790 ( .A1(i_data_bus[499]), .A2(n10506), .B1(
        i_data_bus[403]), .B2(n10505), .ZN(n6686) );
  AOI22D1BWP30P140LVT U9791 ( .A1(i_data_bus[467]), .A2(n10508), .B1(
        i_data_bus[435]), .B2(n10507), .ZN(n6685) );
  ND2D1BWP30P140LVT U9792 ( .A1(n6686), .A2(n6685), .ZN(N8734) );
  AOI22D1BWP30P140LVT U9793 ( .A1(i_data_bus[493]), .A2(n10412), .B1(
        i_data_bus[461]), .B2(n10410), .ZN(n6688) );
  AOI22D1BWP30P140LVT U9794 ( .A1(i_data_bus[429]), .A2(n10411), .B1(
        i_data_bus[397]), .B2(n10409), .ZN(n6687) );
  ND2D1BWP30P140LVT U9795 ( .A1(n6688), .A2(n6687), .ZN(N14350) );
  AOI22D1BWP30P140LVT U9796 ( .A1(i_data_bus[496]), .A2(n10412), .B1(
        i_data_bus[464]), .B2(n10410), .ZN(n6690) );
  AOI22D1BWP30P140LVT U9797 ( .A1(i_data_bus[432]), .A2(n10411), .B1(
        i_data_bus[400]), .B2(n10409), .ZN(n6689) );
  ND2D1BWP30P140LVT U9798 ( .A1(n6690), .A2(n6689), .ZN(N14353) );
  AOI22D1BWP30P140LVT U9799 ( .A1(i_data_bus[507]), .A2(n10412), .B1(
        i_data_bus[475]), .B2(n10410), .ZN(n6692) );
  AOI22D1BWP30P140LVT U9800 ( .A1(i_data_bus[443]), .A2(n10411), .B1(
        i_data_bus[411]), .B2(n10409), .ZN(n6691) );
  ND2D1BWP30P140LVT U9801 ( .A1(n6692), .A2(n6691), .ZN(N14364) );
  AOI22D1BWP30P140LVT U9802 ( .A1(i_data_bus[401]), .A2(n10409), .B1(
        i_data_bus[465]), .B2(n10410), .ZN(n6694) );
  AOI22D1BWP30P140LVT U9803 ( .A1(i_data_bus[433]), .A2(n10411), .B1(
        i_data_bus[497]), .B2(n10412), .ZN(n6693) );
  ND2D1BWP30P140LVT U9804 ( .A1(n6694), .A2(n6693), .ZN(N14354) );
  AOI22D1BWP30P140LVT U9805 ( .A1(i_data_bus[384]), .A2(n10409), .B1(
        i_data_bus[448]), .B2(n10410), .ZN(n6696) );
  AOI22D1BWP30P140LVT U9806 ( .A1(i_data_bus[416]), .A2(n10411), .B1(
        i_data_bus[480]), .B2(n10412), .ZN(n6695) );
  ND2D1BWP30P140LVT U9807 ( .A1(n6696), .A2(n6695), .ZN(N14337) );
  AOI22D1BWP30P140LVT U9808 ( .A1(i_data_bus[446]), .A2(n10411), .B1(
        i_data_bus[478]), .B2(n10410), .ZN(n6698) );
  AOI22D1BWP30P140LVT U9809 ( .A1(i_data_bus[414]), .A2(n10409), .B1(
        i_data_bus[510]), .B2(n10412), .ZN(n6697) );
  ND2D1BWP30P140LVT U9810 ( .A1(n6698), .A2(n6697), .ZN(N14367) );
  AOI22D1BWP30P140LVT U9811 ( .A1(i_data_bus[399]), .A2(n10409), .B1(
        i_data_bus[463]), .B2(n10410), .ZN(n6700) );
  AOI22D1BWP30P140LVT U9812 ( .A1(i_data_bus[431]), .A2(n10411), .B1(
        i_data_bus[495]), .B2(n10412), .ZN(n6699) );
  ND2D1BWP30P140LVT U9813 ( .A1(n6700), .A2(n6699), .ZN(N14352) );
  NR4D1BWP30P140LVT U9814 ( .A1(i_cmd[227]), .A2(n6703), .A3(n10024), .A4(
        n6701), .ZN(n10522) );
  INR4D1BWP30P140LVT U9815 ( .A1(i_cmd[251]), .B1(i_cmd[235]), .B2(n10030), 
        .B3(n6704), .ZN(n10523) );
  AOI22D1BWP30P140LVT U9816 ( .A1(i_data_bus[988]), .A2(n10522), .B1(
        i_data_bus[1020]), .B2(n10523), .ZN(n6706) );
  NR4D1BWP30P140LVT U9817 ( .A1(i_cmd[243]), .A2(n6703), .A3(n10028), .A4(
        n6702), .ZN(n10524) );
  INR4D1BWP30P140LVT U9818 ( .A1(i_cmd[235]), .B1(i_cmd[251]), .B2(n10023), 
        .B3(n6704), .ZN(n10521) );
  AOI22D1BWP30P140LVT U9819 ( .A1(i_data_bus[924]), .A2(n10524), .B1(
        i_data_bus[956]), .B2(n10521), .ZN(n6705) );
  ND2D1BWP30P140LVT U9820 ( .A1(n6706), .A2(n6705), .ZN(N7733) );
  AOI22D1BWP30P140LVT U9821 ( .A1(i_data_bus[925]), .A2(n10524), .B1(
        i_data_bus[1021]), .B2(n10523), .ZN(n6708) );
  AOI22D1BWP30P140LVT U9822 ( .A1(i_data_bus[989]), .A2(n10522), .B1(
        i_data_bus[957]), .B2(n10521), .ZN(n6707) );
  ND2D1BWP30P140LVT U9823 ( .A1(n6708), .A2(n6707), .ZN(N7734) );
  AOI22D1BWP30P140LVT U9824 ( .A1(i_data_bus[962]), .A2(n10522), .B1(
        i_data_bus[994]), .B2(n10523), .ZN(n6710) );
  AOI22D1BWP30P140LVT U9825 ( .A1(i_data_bus[898]), .A2(n10524), .B1(
        i_data_bus[930]), .B2(n10521), .ZN(n6709) );
  ND2D1BWP30P140LVT U9826 ( .A1(n6710), .A2(n6709), .ZN(N7707) );
  AOI22D1BWP30P140LVT U9827 ( .A1(i_data_bus[970]), .A2(n10522), .B1(
        i_data_bus[1002]), .B2(n10523), .ZN(n6712) );
  AOI22D1BWP30P140LVT U9828 ( .A1(i_data_bus[906]), .A2(n10524), .B1(
        i_data_bus[938]), .B2(n10521), .ZN(n6711) );
  ND2D1BWP30P140LVT U9829 ( .A1(n6712), .A2(n6711), .ZN(N7715) );
  AOI22D1BWP30P140LVT U9830 ( .A1(i_data_bus[980]), .A2(n10522), .B1(
        i_data_bus[1012]), .B2(n10523), .ZN(n6714) );
  AOI22D1BWP30P140LVT U9831 ( .A1(i_data_bus[916]), .A2(n10524), .B1(
        i_data_bus[948]), .B2(n10521), .ZN(n6713) );
  ND2D1BWP30P140LVT U9832 ( .A1(n6714), .A2(n6713), .ZN(N7725) );
  INR4D1BWP30P140LVT U9833 ( .A1(i_cmd[170]), .B1(i_cmd[186]), .B2(n9847), 
        .B3(n6715), .ZN(n10564) );
  INR4D1BWP30P140LVT U9834 ( .A1(i_cmd[186]), .B1(i_cmd[170]), .B2(n9844), 
        .B3(n6715), .ZN(n10562) );
  AOI22D1BWP30P140LVT U9835 ( .A1(i_data_bus[703]), .A2(n10564), .B1(
        i_data_bus[767]), .B2(n10562), .ZN(n6720) );
  NR4D1BWP30P140LVT U9836 ( .A1(i_cmd[162]), .A2(n6716), .A3(n9850), .A4(n6717), .ZN(n10561) );
  NR4D1BWP30P140LVT U9837 ( .A1(i_cmd[178]), .A2(n9843), .A3(n6718), .A4(n6717), .ZN(n10563) );
  AOI22D1BWP30P140LVT U9838 ( .A1(i_data_bus[735]), .A2(n10561), .B1(
        i_data_bus[671]), .B2(n10563), .ZN(n6719) );
  ND2D1BWP30P140LVT U9839 ( .A1(n6720), .A2(n6719), .ZN(N5430) );
  AOI22D1BWP30P140LVT U9840 ( .A1(i_data_bus[709]), .A2(n10561), .B1(
        i_data_bus[741]), .B2(n10562), .ZN(n6722) );
  AOI22D1BWP30P140LVT U9841 ( .A1(i_data_bus[677]), .A2(n10564), .B1(
        i_data_bus[645]), .B2(n10563), .ZN(n6721) );
  ND2D1BWP30P140LVT U9842 ( .A1(n6722), .A2(n6721), .ZN(N5404) );
  AOI22D1BWP30P140LVT U9843 ( .A1(i_data_bus[679]), .A2(n10564), .B1(
        i_data_bus[743]), .B2(n10562), .ZN(n6724) );
  AOI22D1BWP30P140LVT U9844 ( .A1(i_data_bus[711]), .A2(n10561), .B1(
        i_data_bus[647]), .B2(n10563), .ZN(n6723) );
  ND2D1BWP30P140LVT U9845 ( .A1(n6724), .A2(n6723), .ZN(N5406) );
  AOI22D1BWP30P140LVT U9846 ( .A1(i_data_bus[686]), .A2(n10564), .B1(
        i_data_bus[718]), .B2(n10561), .ZN(n6726) );
  AOI22D1BWP30P140LVT U9847 ( .A1(i_data_bus[750]), .A2(n10562), .B1(
        i_data_bus[654]), .B2(n10563), .ZN(n6725) );
  ND2D1BWP30P140LVT U9848 ( .A1(n6726), .A2(n6725), .ZN(N5413) );
  AOI22D1BWP30P140LVT U9849 ( .A1(i_data_bus[704]), .A2(n10561), .B1(
        i_data_bus[736]), .B2(n10562), .ZN(n6728) );
  AOI22D1BWP30P140LVT U9850 ( .A1(i_data_bus[672]), .A2(n10564), .B1(
        i_data_bus[640]), .B2(n10563), .ZN(n6727) );
  ND2D1BWP30P140LVT U9851 ( .A1(n6728), .A2(n6727), .ZN(N5399) );
  AOI22D1BWP30P140LVT U9852 ( .A1(i_data_bus[740]), .A2(n10562), .B1(
        i_data_bus[676]), .B2(n10564), .ZN(n6730) );
  AOI22D1BWP30P140LVT U9853 ( .A1(i_data_bus[708]), .A2(n10561), .B1(
        i_data_bus[644]), .B2(n10563), .ZN(n6729) );
  ND2D1BWP30P140LVT U9854 ( .A1(n6730), .A2(n6729), .ZN(N5403) );
  AOI22D1BWP30P140LVT U9855 ( .A1(i_data_bus[725]), .A2(n10561), .B1(
        i_data_bus[693]), .B2(n10564), .ZN(n6732) );
  AOI22D1BWP30P140LVT U9856 ( .A1(i_data_bus[757]), .A2(n10562), .B1(
        i_data_bus[661]), .B2(n10563), .ZN(n6731) );
  ND2D1BWP30P140LVT U9857 ( .A1(n6732), .A2(n6731), .ZN(N5420) );
  AOI22D1BWP30P140LVT U9858 ( .A1(i_data_bus[694]), .A2(n10564), .B1(
        i_data_bus[758]), .B2(n10562), .ZN(n6734) );
  AOI22D1BWP30P140LVT U9859 ( .A1(i_data_bus[726]), .A2(n10561), .B1(
        i_data_bus[662]), .B2(n10563), .ZN(n6733) );
  ND2D1BWP30P140LVT U9860 ( .A1(n6734), .A2(n6733), .ZN(N5421) );
  AOI22D1BWP30P140LVT U9861 ( .A1(i_data_bus[754]), .A2(n10562), .B1(
        i_data_bus[690]), .B2(n10564), .ZN(n6736) );
  AOI22D1BWP30P140LVT U9862 ( .A1(i_data_bus[722]), .A2(n10561), .B1(
        i_data_bus[658]), .B2(n10563), .ZN(n6735) );
  ND2D1BWP30P140LVT U9863 ( .A1(n6736), .A2(n6735), .ZN(N5417) );
  AOI22D1BWP30P140LVT U9864 ( .A1(i_data_bus[752]), .A2(n10562), .B1(
        i_data_bus[688]), .B2(n10564), .ZN(n6738) );
  AOI22D1BWP30P140LVT U9865 ( .A1(i_data_bus[720]), .A2(n10561), .B1(
        i_data_bus[656]), .B2(n10563), .ZN(n6737) );
  ND2D1BWP30P140LVT U9866 ( .A1(n6738), .A2(n6737), .ZN(N5415) );
  INR4D1BWP30P140LVT U9867 ( .A1(i_cmd[187]), .B1(i_cmd[171]), .B2(n9844), 
        .B3(n6739), .ZN(n10530) );
  INR4D1BWP30P140LVT U9868 ( .A1(i_cmd[171]), .B1(i_cmd[187]), .B2(n9847), 
        .B3(n6739), .ZN(n10532) );
  AOI22D1BWP30P140LVT U9869 ( .A1(i_data_bus[763]), .A2(n10530), .B1(
        i_data_bus[699]), .B2(n10532), .ZN(n6744) );
  NR4D1BWP30P140LVT U9870 ( .A1(i_cmd[179]), .A2(n6740), .A3(n9843), .A4(n6741), .ZN(n10529) );
  NR4D1BWP30P140LVT U9871 ( .A1(i_cmd[163]), .A2(n9850), .A3(n6742), .A4(n6741), .ZN(n10531) );
  AOI22D1BWP30P140LVT U9872 ( .A1(i_data_bus[667]), .A2(n10529), .B1(
        i_data_bus[731]), .B2(n10531), .ZN(n6743) );
  ND2D1BWP30P140LVT U9873 ( .A1(n6744), .A2(n6743), .ZN(N7300) );
  AOI22D1BWP30P140LVT U9874 ( .A1(i_data_bus[640]), .A2(n10529), .B1(
        i_data_bus[736]), .B2(n10530), .ZN(n6746) );
  AOI22D1BWP30P140LVT U9875 ( .A1(i_data_bus[672]), .A2(n10532), .B1(
        i_data_bus[704]), .B2(n10531), .ZN(n6745) );
  ND2D1BWP30P140LVT U9876 ( .A1(n6746), .A2(n6745), .ZN(N7273) );
  AOI22D1BWP30P140LVT U9877 ( .A1(i_data_bus[673]), .A2(n10532), .B1(
        i_data_bus[641]), .B2(n10529), .ZN(n6748) );
  AOI22D1BWP30P140LVT U9878 ( .A1(i_data_bus[737]), .A2(n10530), .B1(
        i_data_bus[705]), .B2(n10531), .ZN(n6747) );
  ND2D1BWP30P140LVT U9879 ( .A1(n6748), .A2(n6747), .ZN(N7274) );
  AOI22D1BWP30P140LVT U9880 ( .A1(i_data_bus[675]), .A2(n10532), .B1(
        i_data_bus[739]), .B2(n10530), .ZN(n6750) );
  AOI22D1BWP30P140LVT U9881 ( .A1(i_data_bus[643]), .A2(n10529), .B1(
        i_data_bus[707]), .B2(n10531), .ZN(n6749) );
  ND2D1BWP30P140LVT U9882 ( .A1(n6750), .A2(n6749), .ZN(N7276) );
  AOI22D1BWP30P140LVT U9883 ( .A1(i_data_bus[653]), .A2(n10529), .B1(
        i_data_bus[685]), .B2(n10532), .ZN(n6752) );
  AOI22D1BWP30P140LVT U9884 ( .A1(i_data_bus[749]), .A2(n10530), .B1(
        i_data_bus[717]), .B2(n10531), .ZN(n6751) );
  ND2D1BWP30P140LVT U9885 ( .A1(n6752), .A2(n6751), .ZN(N7286) );
  AOI22D1BWP30P140LVT U9886 ( .A1(i_data_bus[753]), .A2(n10530), .B1(
        i_data_bus[689]), .B2(n10532), .ZN(n6754) );
  AOI22D1BWP30P140LVT U9887 ( .A1(i_data_bus[657]), .A2(n10529), .B1(
        i_data_bus[721]), .B2(n10531), .ZN(n6753) );
  ND2D1BWP30P140LVT U9888 ( .A1(n6754), .A2(n6753), .ZN(N7290) );
  AOI22D1BWP30P140LVT U9889 ( .A1(i_data_bus[230]), .A2(n10484), .B1(
        i_data_bus[134]), .B2(n10481), .ZN(n6756) );
  AOI22D1BWP30P140LVT U9890 ( .A1(i_data_bus[198]), .A2(n10482), .B1(
        i_data_bus[166]), .B2(n10483), .ZN(n6755) );
  ND2D1BWP30P140LVT U9891 ( .A1(n6756), .A2(n6755), .ZN(N10163) );
  AOI22D1BWP30P140LVT U9892 ( .A1(i_data_bus[253]), .A2(n10484), .B1(
        i_data_bus[157]), .B2(n10481), .ZN(n6758) );
  AOI22D1BWP30P140LVT U9893 ( .A1(i_data_bus[221]), .A2(n10482), .B1(
        i_data_bus[189]), .B2(n10483), .ZN(n6757) );
  ND2D1BWP30P140LVT U9894 ( .A1(n6758), .A2(n6757), .ZN(N10186) );
  AOI22D1BWP30P140LVT U9895 ( .A1(i_data_bus[38]), .A2(n10453), .B1(
        i_data_bus[70]), .B2(n10454), .ZN(n6760) );
  AOI22D1BWP30P140LVT U9896 ( .A1(i_data_bus[6]), .A2(n10456), .B1(
        i_data_bus[102]), .B2(n10455), .ZN(n6759) );
  ND2D1BWP30P140LVT U9897 ( .A1(n6760), .A2(n6759), .ZN(N11821) );
  AOI22D1BWP30P140LVT U9898 ( .A1(i_data_bus[17]), .A2(n10456), .B1(
        i_data_bus[81]), .B2(n10454), .ZN(n6762) );
  AOI22D1BWP30P140LVT U9899 ( .A1(i_data_bus[49]), .A2(n10453), .B1(
        i_data_bus[113]), .B2(n10455), .ZN(n6761) );
  ND2D1BWP30P140LVT U9900 ( .A1(n6762), .A2(n6761), .ZN(N11832) );
  AOI22D1BWP30P140LVT U9901 ( .A1(i_data_bus[47]), .A2(n10453), .B1(
        i_data_bus[79]), .B2(n10454), .ZN(n6764) );
  AOI22D1BWP30P140LVT U9902 ( .A1(i_data_bus[15]), .A2(n10456), .B1(
        i_data_bus[111]), .B2(n10455), .ZN(n6763) );
  ND2D1BWP30P140LVT U9903 ( .A1(n6764), .A2(n6763), .ZN(N11830) );
  AOI22D1BWP30P140LVT U9904 ( .A1(i_data_bus[410]), .A2(n10537), .B1(
        i_data_bus[442]), .B2(n10540), .ZN(n6766) );
  AOI22D1BWP30P140LVT U9905 ( .A1(i_data_bus[506]), .A2(n10539), .B1(
        i_data_bus[474]), .B2(n10538), .ZN(n6765) );
  ND2D1BWP30P140LVT U9906 ( .A1(n6766), .A2(n6765), .ZN(N6867) );
  AOI22D1BWP30P140LVT U9907 ( .A1(i_data_bus[414]), .A2(n10537), .B1(
        i_data_bus[446]), .B2(n10540), .ZN(n6768) );
  AOI22D1BWP30P140LVT U9908 ( .A1(i_data_bus[510]), .A2(n10539), .B1(
        i_data_bus[478]), .B2(n10538), .ZN(n6767) );
  ND2D1BWP30P140LVT U9909 ( .A1(n6768), .A2(n6767), .ZN(N6871) );
  AOI22D1BWP30P140LVT U9910 ( .A1(i_data_bus[406]), .A2(n10537), .B1(
        i_data_bus[438]), .B2(n10540), .ZN(n6770) );
  AOI22D1BWP30P140LVT U9911 ( .A1(i_data_bus[502]), .A2(n10539), .B1(
        i_data_bus[470]), .B2(n10538), .ZN(n6769) );
  ND2D1BWP30P140LVT U9912 ( .A1(n6770), .A2(n6769), .ZN(N6863) );
  AOI22D1BWP30P140LVT U9913 ( .A1(i_data_bus[452]), .A2(n10538), .B1(
        i_data_bus[420]), .B2(n10540), .ZN(n6772) );
  AOI22D1BWP30P140LVT U9914 ( .A1(i_data_bus[388]), .A2(n10537), .B1(
        i_data_bus[484]), .B2(n10539), .ZN(n6771) );
  ND2D1BWP30P140LVT U9915 ( .A1(n6772), .A2(n6771), .ZN(N6845) );
  AOI22D1BWP30P140LVT U9916 ( .A1(i_data_bus[878]), .A2(n10398), .B1(
        i_data_bus[846]), .B2(n10399), .ZN(n6774) );
  AOI22D1BWP30P140LVT U9917 ( .A1(i_data_bus[814]), .A2(n10400), .B1(
        i_data_bus[782]), .B2(n10397), .ZN(n6773) );
  ND2D1BWP30P140LVT U9918 ( .A1(n6774), .A2(n6773), .ZN(N14999) );
  AOI22D1BWP30P140LVT U9919 ( .A1(i_data_bus[871]), .A2(n10398), .B1(
        i_data_bus[839]), .B2(n10399), .ZN(n6776) );
  AOI22D1BWP30P140LVT U9920 ( .A1(i_data_bus[807]), .A2(n10400), .B1(
        i_data_bus[775]), .B2(n10397), .ZN(n6775) );
  ND2D1BWP30P140LVT U9921 ( .A1(n6776), .A2(n6775), .ZN(N14992) );
  AOI22D1BWP30P140LVT U9922 ( .A1(i_data_bus[827]), .A2(n10400), .B1(
        i_data_bus[859]), .B2(n10399), .ZN(n6778) );
  AOI22D1BWP30P140LVT U9923 ( .A1(i_data_bus[891]), .A2(n10398), .B1(
        i_data_bus[795]), .B2(n10397), .ZN(n6777) );
  ND2D1BWP30P140LVT U9924 ( .A1(n6778), .A2(n6777), .ZN(N15012) );
  AOI22D1BWP30P140LVT U9925 ( .A1(i_data_bus[820]), .A2(n10400), .B1(
        i_data_bus[852]), .B2(n10399), .ZN(n6780) );
  AOI22D1BWP30P140LVT U9926 ( .A1(i_data_bus[884]), .A2(n10398), .B1(
        i_data_bus[788]), .B2(n10397), .ZN(n6779) );
  ND2D1BWP30P140LVT U9927 ( .A1(n6780), .A2(n6779), .ZN(N15005) );
  AOI22D1BWP30P140LVT U9928 ( .A1(i_data_bus[813]), .A2(n10400), .B1(
        i_data_bus[877]), .B2(n10398), .ZN(n6782) );
  AOI22D1BWP30P140LVT U9929 ( .A1(i_data_bus[845]), .A2(n10399), .B1(
        i_data_bus[781]), .B2(n10397), .ZN(n6781) );
  ND2D1BWP30P140LVT U9930 ( .A1(n6782), .A2(n6781), .ZN(N14998) );
  INR4D1BWP30P140LVT U9931 ( .A1(i_cmd[59]), .B1(i_cmd[43]), .B2(n9860), .B3(
        n6786), .ZN(n10547) );
  NR4D1BWP30P140LVT U9932 ( .A1(i_cmd[35]), .A2(n6785), .A3(n9854), .A4(n6783), 
        .ZN(n10548) );
  AOI22D1BWP30P140LVT U9933 ( .A1(i_data_bus[229]), .A2(n10547), .B1(
        i_data_bus[197]), .B2(n10548), .ZN(n6788) );
  NR4D1BWP30P140LVT U9934 ( .A1(i_cmd[51]), .A2(n6785), .A3(n9857), .A4(n6784), 
        .ZN(n10546) );
  INR4D1BWP30P140LVT U9935 ( .A1(i_cmd[43]), .B1(i_cmd[59]), .B2(n9853), .B3(
        n6786), .ZN(n10545) );
  AOI22D1BWP30P140LVT U9936 ( .A1(i_data_bus[133]), .A2(n10546), .B1(
        i_data_bus[165]), .B2(n10545), .ZN(n6787) );
  ND2D1BWP30P140LVT U9937 ( .A1(n6788), .A2(n6787), .ZN(N6414) );
  AOI22D1BWP30P140LVT U9938 ( .A1(i_data_bus[832]), .A2(n10557), .B1(
        i_data_bus[768]), .B2(n10558), .ZN(n6790) );
  AOI22D1BWP30P140LVT U9939 ( .A1(i_data_bus[800]), .A2(n10560), .B1(
        i_data_bus[864]), .B2(n10559), .ZN(n6789) );
  ND2D1BWP30P140LVT U9940 ( .A1(n6790), .A2(n6789), .ZN(N5615) );
  AOI22D1BWP30P140LVT U9941 ( .A1(i_data_bus[813]), .A2(n10560), .B1(
        i_data_bus[781]), .B2(n10558), .ZN(n6792) );
  AOI22D1BWP30P140LVT U9942 ( .A1(i_data_bus[845]), .A2(n10557), .B1(
        i_data_bus[877]), .B2(n10559), .ZN(n6791) );
  ND2D1BWP30P140LVT U9943 ( .A1(n6792), .A2(n6791), .ZN(N5628) );
  AOI22D1BWP30P140LVT U9944 ( .A1(i_data_bus[857]), .A2(n10557), .B1(
        i_data_bus[793]), .B2(n10558), .ZN(n6794) );
  AOI22D1BWP30P140LVT U9945 ( .A1(i_data_bus[825]), .A2(n10560), .B1(
        i_data_bus[889]), .B2(n10559), .ZN(n6793) );
  ND2D1BWP30P140LVT U9946 ( .A1(n6794), .A2(n6793), .ZN(N5640) );
  AOI22D1BWP30P140LVT U9947 ( .A1(i_data_bus[1005]), .A2(n10457), .B1(
        i_data_bus[941]), .B2(n10460), .ZN(n6796) );
  AOI22D1BWP30P140LVT U9948 ( .A1(i_data_bus[973]), .A2(n10459), .B1(
        i_data_bus[909]), .B2(n10458), .ZN(n6795) );
  ND2D1BWP30P140LVT U9949 ( .A1(n6796), .A2(n6795), .ZN(N11466) );
  AOI22D1BWP30P140LVT U9950 ( .A1(i_data_bus[976]), .A2(n10459), .B1(
        i_data_bus[944]), .B2(n10460), .ZN(n6798) );
  AOI22D1BWP30P140LVT U9951 ( .A1(i_data_bus[1008]), .A2(n10457), .B1(
        i_data_bus[912]), .B2(n10458), .ZN(n6797) );
  ND2D1BWP30P140LVT U9952 ( .A1(n6798), .A2(n6797), .ZN(N11469) );
  AOI22D1BWP30P140LVT U9953 ( .A1(i_data_bus[968]), .A2(n10459), .B1(
        i_data_bus[1000]), .B2(n10457), .ZN(n6800) );
  AOI22D1BWP30P140LVT U9954 ( .A1(i_data_bus[936]), .A2(n10460), .B1(
        i_data_bus[904]), .B2(n10458), .ZN(n6799) );
  ND2D1BWP30P140LVT U9955 ( .A1(n6800), .A2(n6799), .ZN(N11461) );
  AOI22D1BWP30P140LVT U9956 ( .A1(i_data_bus[987]), .A2(n10459), .B1(
        i_data_bus[1019]), .B2(n10457), .ZN(n6802) );
  AOI22D1BWP30P140LVT U9957 ( .A1(i_data_bus[955]), .A2(n10460), .B1(
        i_data_bus[923]), .B2(n10458), .ZN(n6801) );
  ND2D1BWP30P140LVT U9958 ( .A1(n6802), .A2(n6801), .ZN(N11480) );
  AOI22D1BWP30P140LVT U9959 ( .A1(i_data_bus[1013]), .A2(n10457), .B1(
        i_data_bus[949]), .B2(n10460), .ZN(n6804) );
  AOI22D1BWP30P140LVT U9960 ( .A1(i_data_bus[981]), .A2(n10459), .B1(
        i_data_bus[917]), .B2(n10458), .ZN(n6803) );
  ND2D1BWP30P140LVT U9961 ( .A1(n6804), .A2(n6803), .ZN(N11474) );
  AOI22D1BWP30P140LVT U9962 ( .A1(i_data_bus[990]), .A2(n10459), .B1(
        i_data_bus[1022]), .B2(n10457), .ZN(n6806) );
  AOI22D1BWP30P140LVT U9963 ( .A1(i_data_bus[958]), .A2(n10460), .B1(
        i_data_bus[926]), .B2(n10458), .ZN(n6805) );
  ND2D1BWP30P140LVT U9964 ( .A1(n6806), .A2(n6805), .ZN(N11483) );
  AOI22D1BWP30P140LVT U9965 ( .A1(i_data_bus[980]), .A2(n10459), .B1(
        i_data_bus[948]), .B2(n10460), .ZN(n6808) );
  AOI22D1BWP30P140LVT U9966 ( .A1(i_data_bus[1012]), .A2(n10457), .B1(
        i_data_bus[916]), .B2(n10458), .ZN(n6807) );
  ND2D1BWP30P140LVT U9967 ( .A1(n6808), .A2(n6807), .ZN(N11473) );
  AOI22D1BWP30P140LVT U9968 ( .A1(i_data_bus[978]), .A2(n10459), .B1(
        i_data_bus[1010]), .B2(n10457), .ZN(n6810) );
  AOI22D1BWP30P140LVT U9969 ( .A1(i_data_bus[946]), .A2(n10460), .B1(
        i_data_bus[914]), .B2(n10458), .ZN(n6809) );
  ND2D1BWP30P140LVT U9970 ( .A1(n6810), .A2(n6809), .ZN(N11471) );
  AOI22D1BWP30P140LVT U9971 ( .A1(i_data_bus[372]), .A2(n10511), .B1(
        i_data_bus[340]), .B2(n10509), .ZN(n6812) );
  AOI22D1BWP30P140LVT U9972 ( .A1(i_data_bus[308]), .A2(n10512), .B1(
        i_data_bus[276]), .B2(n10510), .ZN(n6811) );
  ND2D1BWP30P140LVT U9973 ( .A1(n6812), .A2(n6811), .ZN(N8519) );
  AOI22D1BWP30P140LVT U9974 ( .A1(i_data_bus[328]), .A2(n10509), .B1(
        i_data_bus[296]), .B2(n10512), .ZN(n6814) );
  AOI22D1BWP30P140LVT U9975 ( .A1(i_data_bus[360]), .A2(n10511), .B1(
        i_data_bus[264]), .B2(n10510), .ZN(n6813) );
  ND2D1BWP30P140LVT U9976 ( .A1(n6814), .A2(n6813), .ZN(N8507) );
  INR4D1BWP30P140LVT U9977 ( .A1(i_cmd[249]), .B1(i_cmd[233]), .B2(n10030), 
        .B3(n6818), .ZN(n10585) );
  NR4D1BWP30P140LVT U9978 ( .A1(i_cmd[241]), .A2(n6815), .A3(n10028), .A4(
        n6816), .ZN(n10587) );
  AOI22D1BWP30P140LVT U9979 ( .A1(i_data_bus[1001]), .A2(n10585), .B1(
        i_data_bus[905]), .B2(n10587), .ZN(n6820) );
  NR4D1BWP30P140LVT U9980 ( .A1(i_cmd[225]), .A2(n10024), .A3(n6817), .A4(
        n6816), .ZN(n10586) );
  INR4D1BWP30P140LVT U9981 ( .A1(i_cmd[233]), .B1(i_cmd[249]), .B2(n10023), 
        .B3(n6818), .ZN(n10588) );
  AOI22D1BWP30P140LVT U9982 ( .A1(i_data_bus[969]), .A2(n10586), .B1(
        i_data_bus[937]), .B2(n10588), .ZN(n6819) );
  ND2D1BWP30P140LVT U9983 ( .A1(n6820), .A2(n6819), .ZN(N3966) );
  AOI22D1BWP30P140LVT U9984 ( .A1(i_data_bus[921]), .A2(n10587), .B1(
        i_data_bus[1017]), .B2(n10585), .ZN(n6822) );
  AOI22D1BWP30P140LVT U9985 ( .A1(i_data_bus[985]), .A2(n10586), .B1(
        i_data_bus[953]), .B2(n10588), .ZN(n6821) );
  ND2D1BWP30P140LVT U9986 ( .A1(n6822), .A2(n6821), .ZN(N3982) );
  AOI22D1BWP30P140LVT U9987 ( .A1(i_data_bus[906]), .A2(n10587), .B1(
        i_data_bus[1002]), .B2(n10585), .ZN(n6824) );
  AOI22D1BWP30P140LVT U9988 ( .A1(i_data_bus[970]), .A2(n10586), .B1(
        i_data_bus[938]), .B2(n10588), .ZN(n6823) );
  ND2D1BWP30P140LVT U9989 ( .A1(n6824), .A2(n6823), .ZN(N3967) );
  AOI22D1BWP30P140LVT U9990 ( .A1(i_data_bus[992]), .A2(n10585), .B1(
        i_data_bus[960]), .B2(n10586), .ZN(n6826) );
  AOI22D1BWP30P140LVT U9991 ( .A1(i_data_bus[896]), .A2(n10587), .B1(
        i_data_bus[928]), .B2(n10588), .ZN(n6825) );
  ND2D1BWP30P140LVT U9992 ( .A1(n6826), .A2(n6825), .ZN(N3957) );
  AOI22D1BWP30P140LVT U9993 ( .A1(i_data_bus[898]), .A2(n10587), .B1(
        i_data_bus[962]), .B2(n10586), .ZN(n6828) );
  AOI22D1BWP30P140LVT U9994 ( .A1(i_data_bus[994]), .A2(n10585), .B1(
        i_data_bus[930]), .B2(n10588), .ZN(n6827) );
  ND2D1BWP30P140LVT U9995 ( .A1(n6828), .A2(n6827), .ZN(N3959) );
  AOI22D1BWP30P140LVT U9996 ( .A1(i_data_bus[980]), .A2(n10586), .B1(
        i_data_bus[1012]), .B2(n10585), .ZN(n6830) );
  AOI22D1BWP30P140LVT U9997 ( .A1(i_data_bus[916]), .A2(n10587), .B1(
        i_data_bus[948]), .B2(n10588), .ZN(n6829) );
  ND2D1BWP30P140LVT U9998 ( .A1(n6830), .A2(n6829), .ZN(N3977) );
  AOI22D1BWP30P140LVT U9999 ( .A1(i_data_bus[910]), .A2(n10587), .B1(
        i_data_bus[1006]), .B2(n10585), .ZN(n6832) );
  AOI22D1BWP30P140LVT U10000 ( .A1(i_data_bus[974]), .A2(n10586), .B1(
        i_data_bus[942]), .B2(n10588), .ZN(n6831) );
  ND2D1BWP30P140LVT U10001 ( .A1(n6832), .A2(n6831), .ZN(N3971) );
  AOI22D1BWP30P140LVT U10002 ( .A1(i_data_bus[405]), .A2(n10505), .B1(
        i_data_bus[469]), .B2(n10508), .ZN(n6834) );
  AOI22D1BWP30P140LVT U10003 ( .A1(i_data_bus[437]), .A2(n10507), .B1(
        i_data_bus[501]), .B2(n10506), .ZN(n6833) );
  ND2D1BWP30P140LVT U10004 ( .A1(n6834), .A2(n6833), .ZN(N8736) );
  AOI22D1BWP30P140LVT U10005 ( .A1(i_data_bus[427]), .A2(n10507), .B1(
        i_data_bus[459]), .B2(n10508), .ZN(n6836) );
  AOI22D1BWP30P140LVT U10006 ( .A1(i_data_bus[395]), .A2(n10505), .B1(
        i_data_bus[491]), .B2(n10506), .ZN(n6835) );
  ND2D1BWP30P140LVT U10007 ( .A1(n6836), .A2(n6835), .ZN(N8726) );
  INR4D1BWP30P140LVT U10008 ( .A1(i_cmd[42]), .B1(i_cmd[58]), .B2(n9853), .B3(
        n6837), .ZN(n10579) );
  INR4D1BWP30P140LVT U10009 ( .A1(i_cmd[58]), .B1(i_cmd[42]), .B2(n9860), .B3(
        n6837), .ZN(n10580) );
  AOI22D1BWP30P140LVT U10010 ( .A1(i_data_bus[187]), .A2(n10579), .B1(
        i_data_bus[251]), .B2(n10580), .ZN(n6842) );
  NR4D1BWP30P140LVT U10011 ( .A1(i_cmd[50]), .A2(n6838), .A3(n9857), .A4(n6839), .ZN(n10577) );
  NR4D1BWP30P140LVT U10012 ( .A1(i_cmd[34]), .A2(n9854), .A3(n6840), .A4(n6839), .ZN(n10578) );
  AOI22D1BWP30P140LVT U10013 ( .A1(i_data_bus[155]), .A2(n10577), .B1(
        i_data_bus[219]), .B2(n10578), .ZN(n6841) );
  ND2D1BWP30P140LVT U10014 ( .A1(n6842), .A2(n6841), .ZN(N4562) );
  AOI22D1BWP30P140LVT U10015 ( .A1(i_data_bus[149]), .A2(n10577), .B1(
        i_data_bus[245]), .B2(n10580), .ZN(n6844) );
  AOI22D1BWP30P140LVT U10016 ( .A1(i_data_bus[181]), .A2(n10579), .B1(
        i_data_bus[213]), .B2(n10578), .ZN(n6843) );
  ND2D1BWP30P140LVT U10017 ( .A1(n6844), .A2(n6843), .ZN(N4556) );
  AOI22D1BWP30P140LVT U10018 ( .A1(i_data_bus[375]), .A2(n10608), .B1(
        i_data_bus[343]), .B2(n10607), .ZN(n6846) );
  AOI22D1BWP30P140LVT U10019 ( .A1(i_data_bus[279]), .A2(n10605), .B1(
        i_data_bus[311]), .B2(n10606), .ZN(n6845) );
  ND2D1BWP30P140LVT U10020 ( .A1(n6846), .A2(n6845), .ZN(N2900) );
  AOI22D1BWP30P140LVT U10021 ( .A1(i_data_bus[340]), .A2(n10607), .B1(
        i_data_bus[276]), .B2(n10605), .ZN(n6848) );
  AOI22D1BWP30P140LVT U10022 ( .A1(i_data_bus[372]), .A2(n10608), .B1(
        i_data_bus[308]), .B2(n10606), .ZN(n6847) );
  ND2D1BWP30P140LVT U10023 ( .A1(n6848), .A2(n6847), .ZN(N2897) );
  AOI22D1BWP30P140LVT U10024 ( .A1(i_data_bus[365]), .A2(n10608), .B1(
        i_data_bus[333]), .B2(n10607), .ZN(n6850) );
  AOI22D1BWP30P140LVT U10025 ( .A1(i_data_bus[269]), .A2(n10605), .B1(
        i_data_bus[301]), .B2(n10606), .ZN(n6849) );
  ND2D1BWP30P140LVT U10026 ( .A1(n6850), .A2(n6849), .ZN(N2890) );
  AOI22D1BWP30P140LVT U10027 ( .A1(i_data_bus[481]), .A2(n10506), .B1(
        i_data_bus[449]), .B2(n10508), .ZN(n6852) );
  AOI22D1BWP30P140LVT U10028 ( .A1(i_data_bus[385]), .A2(n10505), .B1(
        i_data_bus[417]), .B2(n10507), .ZN(n6851) );
  ND2D1BWP30P140LVT U10029 ( .A1(n6852), .A2(n6851), .ZN(N8716) );
  AOI22D1BWP30P140LVT U10030 ( .A1(i_data_bus[510]), .A2(n10506), .B1(
        i_data_bus[478]), .B2(n10508), .ZN(n6854) );
  AOI22D1BWP30P140LVT U10031 ( .A1(i_data_bus[414]), .A2(n10505), .B1(
        i_data_bus[446]), .B2(n10507), .ZN(n6853) );
  ND2D1BWP30P140LVT U10032 ( .A1(n6854), .A2(n6853), .ZN(N8745) );
  AOI22D1BWP30P140LVT U10033 ( .A1(i_data_bus[338]), .A2(n10607), .B1(
        i_data_bus[274]), .B2(n10605), .ZN(n6856) );
  AOI22D1BWP30P140LVT U10034 ( .A1(i_data_bus[370]), .A2(n10608), .B1(
        i_data_bus[306]), .B2(n10606), .ZN(n6855) );
  ND2D1BWP30P140LVT U10035 ( .A1(n6856), .A2(n6855), .ZN(N2895) );
  AOI22D1BWP30P140LVT U10036 ( .A1(i_data_bus[262]), .A2(n10605), .B1(
        i_data_bus[326]), .B2(n10607), .ZN(n6858) );
  AOI22D1BWP30P140LVT U10037 ( .A1(i_data_bus[358]), .A2(n10608), .B1(
        i_data_bus[294]), .B2(n10606), .ZN(n6857) );
  ND2D1BWP30P140LVT U10038 ( .A1(n6858), .A2(n6857), .ZN(N2883) );
  AOI22D1BWP30P140LVT U10039 ( .A1(i_data_bus[357]), .A2(n10608), .B1(
        i_data_bus[261]), .B2(n10605), .ZN(n6860) );
  AOI22D1BWP30P140LVT U10040 ( .A1(i_data_bus[325]), .A2(n10607), .B1(
        i_data_bus[293]), .B2(n10606), .ZN(n6859) );
  ND2D1BWP30P140LVT U10041 ( .A1(n6860), .A2(n6859), .ZN(N2882) );
  AOI22D1BWP30P140LVT U10042 ( .A1(i_data_bus[360]), .A2(n10608), .B1(
        i_data_bus[264]), .B2(n10605), .ZN(n6862) );
  AOI22D1BWP30P140LVT U10043 ( .A1(i_data_bus[328]), .A2(n10607), .B1(
        i_data_bus[296]), .B2(n10606), .ZN(n6861) );
  ND2D1BWP30P140LVT U10044 ( .A1(n6862), .A2(n6861), .ZN(N2885) );
  AOI22D1BWP30P140LVT U10045 ( .A1(i_data_bus[389]), .A2(n10505), .B1(
        i_data_bus[453]), .B2(n10508), .ZN(n6864) );
  AOI22D1BWP30P140LVT U10046 ( .A1(i_data_bus[485]), .A2(n10506), .B1(
        i_data_bus[421]), .B2(n10507), .ZN(n6863) );
  ND2D1BWP30P140LVT U10047 ( .A1(n6864), .A2(n6863), .ZN(N8720) );
  AOI22D1BWP30P140LVT U10048 ( .A1(i_data_bus[392]), .A2(n10505), .B1(
        i_data_bus[456]), .B2(n10508), .ZN(n6866) );
  AOI22D1BWP30P140LVT U10049 ( .A1(i_data_bus[488]), .A2(n10506), .B1(
        i_data_bus[424]), .B2(n10507), .ZN(n6865) );
  ND2D1BWP30P140LVT U10050 ( .A1(n6866), .A2(n6865), .ZN(N8723) );
  AOI22D1BWP30P140LVT U10051 ( .A1(i_data_bus[406]), .A2(n10505), .B1(
        i_data_bus[470]), .B2(n10508), .ZN(n6868) );
  AOI22D1BWP30P140LVT U10052 ( .A1(i_data_bus[502]), .A2(n10506), .B1(
        i_data_bus[438]), .B2(n10507), .ZN(n6867) );
  ND2D1BWP30P140LVT U10053 ( .A1(n6868), .A2(n6867), .ZN(N8737) );
  AOI22D1BWP30P140LVT U10054 ( .A1(i_data_bus[997]), .A2(n10523), .B1(
        i_data_bus[901]), .B2(n10524), .ZN(n6870) );
  AOI22D1BWP30P140LVT U10055 ( .A1(i_data_bus[965]), .A2(n10522), .B1(
        i_data_bus[933]), .B2(n10521), .ZN(n6869) );
  ND2D1BWP30P140LVT U10056 ( .A1(n6870), .A2(n6869), .ZN(N7710) );
  AOI22D1BWP30P140LVT U10057 ( .A1(i_data_bus[981]), .A2(n10522), .B1(
        i_data_bus[917]), .B2(n10524), .ZN(n6872) );
  AOI22D1BWP30P140LVT U10058 ( .A1(i_data_bus[1013]), .A2(n10523), .B1(
        i_data_bus[949]), .B2(n10521), .ZN(n6871) );
  ND2D1BWP30P140LVT U10059 ( .A1(n6872), .A2(n6871), .ZN(N7726) );
  AOI22D1BWP30P140LVT U10060 ( .A1(i_data_bus[1000]), .A2(n10523), .B1(
        i_data_bus[904]), .B2(n10524), .ZN(n6874) );
  AOI22D1BWP30P140LVT U10061 ( .A1(i_data_bus[968]), .A2(n10522), .B1(
        i_data_bus[936]), .B2(n10521), .ZN(n6873) );
  ND2D1BWP30P140LVT U10062 ( .A1(n6874), .A2(n6873), .ZN(N7713) );
  AOI22D1BWP30P140LVT U10063 ( .A1(i_data_bus[1001]), .A2(n10523), .B1(
        i_data_bus[905]), .B2(n10524), .ZN(n6876) );
  AOI22D1BWP30P140LVT U10064 ( .A1(i_data_bus[969]), .A2(n10522), .B1(
        i_data_bus[937]), .B2(n10521), .ZN(n6875) );
  ND2D1BWP30P140LVT U10065 ( .A1(n6876), .A2(n6875), .ZN(N7714) );
  INR4D1BWP30P140LVT U10066 ( .A1(i_cmd[38]), .B1(i_cmd[54]), .B2(n9857), .B3(
        n6877), .ZN(n10452) );
  INR4D1BWP30P140LVT U10067 ( .A1(i_cmd[54]), .B1(i_cmd[38]), .B2(n9854), .B3(
        n6877), .ZN(n10451) );
  AOI22D1BWP30P140LVT U10068 ( .A1(i_data_bus[155]), .A2(n10452), .B1(
        i_data_bus[219]), .B2(n10451), .ZN(n6882) );
  NR4D1BWP30P140LVT U10069 ( .A1(i_cmd[62]), .A2(n6878), .A3(n9853), .A4(n6879), .ZN(n10450) );
  NR4D1BWP30P140LVT U10070 ( .A1(i_cmd[46]), .A2(n9860), .A3(n6880), .A4(n6879), .ZN(n10449) );
  AOI22D1BWP30P140LVT U10071 ( .A1(i_data_bus[187]), .A2(n10450), .B1(
        i_data_bus[251]), .B2(n10449), .ZN(n6881) );
  ND2D1BWP30P140LVT U10072 ( .A1(n6882), .A2(n6881), .ZN(N12058) );
  AOI22D1BWP30P140LVT U10073 ( .A1(i_data_bus[148]), .A2(n10452), .B1(
        i_data_bus[180]), .B2(n10450), .ZN(n6884) );
  AOI22D1BWP30P140LVT U10074 ( .A1(i_data_bus[212]), .A2(n10451), .B1(
        i_data_bus[244]), .B2(n10449), .ZN(n6883) );
  ND2D1BWP30P140LVT U10075 ( .A1(n6884), .A2(n6883), .ZN(N12051) );
  AOI22D1BWP30P140LVT U10076 ( .A1(i_data_bus[151]), .A2(n10452), .B1(
        i_data_bus[215]), .B2(n10451), .ZN(n6886) );
  AOI22D1BWP30P140LVT U10077 ( .A1(i_data_bus[183]), .A2(n10450), .B1(
        i_data_bus[247]), .B2(n10449), .ZN(n6885) );
  ND2D1BWP30P140LVT U10078 ( .A1(n6886), .A2(n6885), .ZN(N12054) );
  AOI22D1BWP30P140LVT U10079 ( .A1(i_data_bus[207]), .A2(n10451), .B1(
        i_data_bus[175]), .B2(n10450), .ZN(n6888) );
  AOI22D1BWP30P140LVT U10080 ( .A1(i_data_bus[143]), .A2(n10452), .B1(
        i_data_bus[239]), .B2(n10449), .ZN(n6887) );
  ND2D1BWP30P140LVT U10081 ( .A1(n6888), .A2(n6887), .ZN(N12046) );
  AOI22D1BWP30P140LVT U10082 ( .A1(i_data_bus[194]), .A2(n10451), .B1(
        i_data_bus[162]), .B2(n10450), .ZN(n6890) );
  AOI22D1BWP30P140LVT U10083 ( .A1(i_data_bus[130]), .A2(n10452), .B1(
        i_data_bus[226]), .B2(n10449), .ZN(n6889) );
  ND2D1BWP30P140LVT U10084 ( .A1(n6890), .A2(n6889), .ZN(N12033) );
  AOI22D1BWP30P140LVT U10085 ( .A1(i_data_bus[196]), .A2(n10451), .B1(
        i_data_bus[164]), .B2(n10450), .ZN(n6892) );
  AOI22D1BWP30P140LVT U10086 ( .A1(i_data_bus[132]), .A2(n10452), .B1(
        i_data_bus[228]), .B2(n10449), .ZN(n6891) );
  ND2D1BWP30P140LVT U10087 ( .A1(n6892), .A2(n6891), .ZN(N12035) );
  AOI22D1BWP30P140LVT U10088 ( .A1(i_data_bus[161]), .A2(n10450), .B1(
        i_data_bus[193]), .B2(n10451), .ZN(n6894) );
  AOI22D1BWP30P140LVT U10089 ( .A1(i_data_bus[129]), .A2(n10452), .B1(
        i_data_bus[225]), .B2(n10449), .ZN(n6893) );
  ND2D1BWP30P140LVT U10090 ( .A1(n6894), .A2(n6893), .ZN(N12032) );
  AOI22D1BWP30P140LVT U10091 ( .A1(i_data_bus[200]), .A2(n10451), .B1(
        i_data_bus[168]), .B2(n10450), .ZN(n6896) );
  AOI22D1BWP30P140LVT U10092 ( .A1(i_data_bus[136]), .A2(n10452), .B1(
        i_data_bus[232]), .B2(n10449), .ZN(n6895) );
  ND2D1BWP30P140LVT U10093 ( .A1(n6896), .A2(n6895), .ZN(N12039) );
  AOI22D1BWP30P140LVT U10094 ( .A1(i_data_bus[179]), .A2(n10450), .B1(
        i_data_bus[147]), .B2(n10452), .ZN(n6898) );
  AOI22D1BWP30P140LVT U10095 ( .A1(i_data_bus[211]), .A2(n10451), .B1(
        i_data_bus[243]), .B2(n10449), .ZN(n6897) );
  ND2D1BWP30P140LVT U10096 ( .A1(n6898), .A2(n6897), .ZN(N12050) );
  AOI22D1BWP30P140LVT U10097 ( .A1(i_data_bus[206]), .A2(n10451), .B1(
        i_data_bus[142]), .B2(n10452), .ZN(n6900) );
  AOI22D1BWP30P140LVT U10098 ( .A1(i_data_bus[174]), .A2(n10450), .B1(
        i_data_bus[238]), .B2(n10449), .ZN(n6899) );
  ND2D1BWP30P140LVT U10099 ( .A1(n6900), .A2(n6899), .ZN(N12045) );
  AOI22D1BWP30P140LVT U10100 ( .A1(i_data_bus[202]), .A2(n10451), .B1(
        i_data_bus[138]), .B2(n10452), .ZN(n6902) );
  AOI22D1BWP30P140LVT U10101 ( .A1(i_data_bus[170]), .A2(n10450), .B1(
        i_data_bus[234]), .B2(n10449), .ZN(n6901) );
  ND2D1BWP30P140LVT U10102 ( .A1(n6902), .A2(n6901), .ZN(N12041) );
  AOI22D1BWP30P140LVT U10103 ( .A1(i_data_bus[209]), .A2(n10451), .B1(
        i_data_bus[145]), .B2(n10452), .ZN(n6904) );
  AOI22D1BWP30P140LVT U10104 ( .A1(i_data_bus[177]), .A2(n10450), .B1(
        i_data_bus[241]), .B2(n10449), .ZN(n6903) );
  ND2D1BWP30P140LVT U10105 ( .A1(n6904), .A2(n6903), .ZN(N12048) );
  AOI22D1BWP30P140LVT U10106 ( .A1(i_data_bus[489]), .A2(n10571), .B1(
        i_data_bus[393]), .B2(n10572), .ZN(n6906) );
  AOI22D1BWP30P140LVT U10107 ( .A1(i_data_bus[457]), .A2(n10570), .B1(
        i_data_bus[425]), .B2(n10569), .ZN(n6905) );
  ND2D1BWP30P140LVT U10108 ( .A1(n6906), .A2(n6905), .ZN(N4976) );
  AOI22D1BWP30P140LVT U10109 ( .A1(i_data_bus[510]), .A2(n10571), .B1(
        i_data_bus[478]), .B2(n10570), .ZN(n6908) );
  AOI22D1BWP30P140LVT U10110 ( .A1(i_data_bus[414]), .A2(n10572), .B1(
        i_data_bus[446]), .B2(n10569), .ZN(n6907) );
  ND2D1BWP30P140LVT U10111 ( .A1(n6908), .A2(n6907), .ZN(N4997) );
  AOI22D1BWP30P140LVT U10112 ( .A1(i_data_bus[502]), .A2(n10571), .B1(
        i_data_bus[406]), .B2(n10572), .ZN(n6910) );
  AOI22D1BWP30P140LVT U10113 ( .A1(i_data_bus[470]), .A2(n10570), .B1(
        i_data_bus[438]), .B2(n10569), .ZN(n6909) );
  ND2D1BWP30P140LVT U10114 ( .A1(n6910), .A2(n6909), .ZN(N4989) );
  AOI22D1BWP30P140LVT U10115 ( .A1(i_data_bus[465]), .A2(n10570), .B1(
        i_data_bus[497]), .B2(n10571), .ZN(n6912) );
  AOI22D1BWP30P140LVT U10116 ( .A1(i_data_bus[401]), .A2(n10572), .B1(
        i_data_bus[433]), .B2(n10569), .ZN(n6911) );
  ND2D1BWP30P140LVT U10117 ( .A1(n6912), .A2(n6911), .ZN(N4984) );
  AOI22D1BWP30P140LVT U10118 ( .A1(i_data_bus[458]), .A2(n10570), .B1(
        i_data_bus[394]), .B2(n10572), .ZN(n6914) );
  AOI22D1BWP30P140LVT U10119 ( .A1(i_data_bus[490]), .A2(n10571), .B1(
        i_data_bus[426]), .B2(n10569), .ZN(n6913) );
  ND2D1BWP30P140LVT U10120 ( .A1(n6914), .A2(n6913), .ZN(N4977) );
  AOI22D1BWP30P140LVT U10121 ( .A1(i_data_bus[460]), .A2(n10570), .B1(
        i_data_bus[396]), .B2(n10572), .ZN(n6916) );
  AOI22D1BWP30P140LVT U10122 ( .A1(i_data_bus[492]), .A2(n10571), .B1(
        i_data_bus[428]), .B2(n10569), .ZN(n6915) );
  ND2D1BWP30P140LVT U10123 ( .A1(n6916), .A2(n6915), .ZN(N4979) );
  AOI22D1BWP30P140LVT U10124 ( .A1(i_data_bus[464]), .A2(n10570), .B1(
        i_data_bus[400]), .B2(n10572), .ZN(n6918) );
  AOI22D1BWP30P140LVT U10125 ( .A1(i_data_bus[496]), .A2(n10571), .B1(
        i_data_bus[432]), .B2(n10569), .ZN(n6917) );
  ND2D1BWP30P140LVT U10126 ( .A1(n6918), .A2(n6917), .ZN(N4983) );
  AOI22D1BWP30P140LVT U10127 ( .A1(i_data_bus[467]), .A2(n10570), .B1(
        i_data_bus[403]), .B2(n10572), .ZN(n6920) );
  AOI22D1BWP30P140LVT U10128 ( .A1(i_data_bus[499]), .A2(n10571), .B1(
        i_data_bus[435]), .B2(n10569), .ZN(n6919) );
  ND2D1BWP30P140LVT U10129 ( .A1(n6920), .A2(n6919), .ZN(N4986) );
  AOI22D1BWP30P140LVT U10130 ( .A1(i_data_bus[389]), .A2(n10572), .B1(
        i_data_bus[453]), .B2(n10570), .ZN(n6922) );
  AOI22D1BWP30P140LVT U10131 ( .A1(i_data_bus[485]), .A2(n10571), .B1(
        i_data_bus[421]), .B2(n10569), .ZN(n6921) );
  ND2D1BWP30P140LVT U10132 ( .A1(n6922), .A2(n6921), .ZN(N4972) );
  AOI22D1BWP30P140LVT U10133 ( .A1(i_data_bus[413]), .A2(n10572), .B1(
        i_data_bus[477]), .B2(n10570), .ZN(n6924) );
  AOI22D1BWP30P140LVT U10134 ( .A1(i_data_bus[509]), .A2(n10571), .B1(
        i_data_bus[445]), .B2(n10569), .ZN(n6923) );
  ND2D1BWP30P140LVT U10135 ( .A1(n6924), .A2(n6923), .ZN(N4996) );
  AOI22D1BWP30P140LVT U10136 ( .A1(i_data_bus[451]), .A2(n10570), .B1(
        i_data_bus[483]), .B2(n10571), .ZN(n6926) );
  AOI22D1BWP30P140LVT U10137 ( .A1(i_data_bus[387]), .A2(n10572), .B1(
        i_data_bus[419]), .B2(n10569), .ZN(n6925) );
  ND2D1BWP30P140LVT U10138 ( .A1(n6926), .A2(n6925), .ZN(N4970) );
  AOI22D1BWP30P140LVT U10139 ( .A1(i_data_bus[488]), .A2(n10571), .B1(
        i_data_bus[456]), .B2(n10570), .ZN(n6928) );
  AOI22D1BWP30P140LVT U10140 ( .A1(i_data_bus[392]), .A2(n10572), .B1(
        i_data_bus[424]), .B2(n10569), .ZN(n6927) );
  ND2D1BWP30P140LVT U10141 ( .A1(n6928), .A2(n6927), .ZN(N4975) );
  AOI22D1BWP30P140LVT U10142 ( .A1(i_data_bus[415]), .A2(n10572), .B1(
        i_data_bus[511]), .B2(n10571), .ZN(n6930) );
  AOI22D1BWP30P140LVT U10143 ( .A1(i_data_bus[479]), .A2(n10570), .B1(
        i_data_bus[447]), .B2(n10569), .ZN(n6929) );
  ND2D1BWP30P140LVT U10144 ( .A1(n6930), .A2(n6929), .ZN(N4998) );
  AOI22D1BWP30P140LVT U10145 ( .A1(i_data_bus[128]), .A2(n10513), .B1(
        i_data_bus[192]), .B2(n10514), .ZN(n6932) );
  AOI22D1BWP30P140LVT U10146 ( .A1(i_data_bus[224]), .A2(n10516), .B1(
        i_data_bus[160]), .B2(n10515), .ZN(n6931) );
  ND2D1BWP30P140LVT U10147 ( .A1(n6932), .A2(n6931), .ZN(N8283) );
  AOI22D1BWP30P140LVT U10148 ( .A1(i_data_bus[794]), .A2(n10429), .B1(
        i_data_bus[826]), .B2(n10430), .ZN(n6934) );
  AOI22D1BWP30P140LVT U10149 ( .A1(i_data_bus[858]), .A2(n10432), .B1(
        i_data_bus[890]), .B2(n10431), .ZN(n6933) );
  ND2D1BWP30P140LVT U10150 ( .A1(n6934), .A2(n6933), .ZN(N13137) );
  AOI22D1BWP30P140LVT U10151 ( .A1(i_data_bus[843]), .A2(n10432), .B1(
        i_data_bus[811]), .B2(n10430), .ZN(n6936) );
  AOI22D1BWP30P140LVT U10152 ( .A1(i_data_bus[779]), .A2(n10429), .B1(
        i_data_bus[875]), .B2(n10431), .ZN(n6935) );
  ND2D1BWP30P140LVT U10153 ( .A1(n6936), .A2(n6935), .ZN(N13122) );
  AOI22D1BWP30P140LVT U10154 ( .A1(i_data_bus[780]), .A2(n10429), .B1(
        i_data_bus[812]), .B2(n10430), .ZN(n6938) );
  AOI22D1BWP30P140LVT U10155 ( .A1(i_data_bus[844]), .A2(n10432), .B1(
        i_data_bus[876]), .B2(n10431), .ZN(n6937) );
  ND2D1BWP30P140LVT U10156 ( .A1(n6938), .A2(n6937), .ZN(N13123) );
  AOI22D1BWP30P140LVT U10157 ( .A1(i_data_bus[842]), .A2(n10432), .B1(
        i_data_bus[810]), .B2(n10430), .ZN(n6940) );
  AOI22D1BWP30P140LVT U10158 ( .A1(i_data_bus[778]), .A2(n10429), .B1(
        i_data_bus[874]), .B2(n10431), .ZN(n6939) );
  ND2D1BWP30P140LVT U10159 ( .A1(n6940), .A2(n6939), .ZN(N13121) );
  AOI22D1BWP30P140LVT U10160 ( .A1(i_data_bus[796]), .A2(n10429), .B1(
        i_data_bus[828]), .B2(n10430), .ZN(n6942) );
  AOI22D1BWP30P140LVT U10161 ( .A1(i_data_bus[860]), .A2(n10432), .B1(
        i_data_bus[892]), .B2(n10431), .ZN(n6941) );
  ND2D1BWP30P140LVT U10162 ( .A1(n6942), .A2(n6941), .ZN(N13139) );
  AOI22D1BWP30P140LVT U10163 ( .A1(i_data_bus[208]), .A2(n10610), .B1(
        i_data_bus[240]), .B2(n10611), .ZN(n6944) );
  AOI22D1BWP30P140LVT U10164 ( .A1(i_data_bus[144]), .A2(n10612), .B1(
        i_data_bus[176]), .B2(n10609), .ZN(n6943) );
  ND2D1BWP30P140LVT U10165 ( .A1(n6944), .A2(n6943), .ZN(N2677) );
  AOI22D1BWP30P140LVT U10166 ( .A1(i_data_bus[136]), .A2(n10612), .B1(
        i_data_bus[232]), .B2(n10611), .ZN(n6946) );
  AOI22D1BWP30P140LVT U10167 ( .A1(i_data_bus[200]), .A2(n10610), .B1(
        i_data_bus[168]), .B2(n10609), .ZN(n6945) );
  ND2D1BWP30P140LVT U10168 ( .A1(n6946), .A2(n6945), .ZN(N2669) );
  AOI22D1BWP30P140LVT U10169 ( .A1(i_data_bus[158]), .A2(n10612), .B1(
        i_data_bus[254]), .B2(n10611), .ZN(n6948) );
  AOI22D1BWP30P140LVT U10170 ( .A1(i_data_bus[222]), .A2(n10610), .B1(
        i_data_bus[190]), .B2(n10609), .ZN(n6947) );
  ND2D1BWP30P140LVT U10171 ( .A1(n6948), .A2(n6947), .ZN(N2691) );
  AOI22D1BWP30P140LVT U10172 ( .A1(i_data_bus[130]), .A2(n10612), .B1(
        i_data_bus[226]), .B2(n10611), .ZN(n6950) );
  AOI22D1BWP30P140LVT U10173 ( .A1(i_data_bus[194]), .A2(n10610), .B1(
        i_data_bus[162]), .B2(n10609), .ZN(n6949) );
  ND2D1BWP30P140LVT U10174 ( .A1(n6950), .A2(n6949), .ZN(N2663) );
  AOI22D1BWP30P140LVT U10175 ( .A1(i_data_bus[712]), .A2(n10402), .B1(
        i_data_bus[680]), .B2(n10404), .ZN(n6952) );
  AOI22D1BWP30P140LVT U10176 ( .A1(i_data_bus[744]), .A2(n10403), .B1(
        i_data_bus[648]), .B2(n10401), .ZN(n6951) );
  ND2D1BWP30P140LVT U10177 ( .A1(n6952), .A2(n6951), .ZN(N14777) );
  AOI22D1BWP30P140LVT U10178 ( .A1(i_data_bus[730]), .A2(n10402), .B1(
        i_data_bus[762]), .B2(n10403), .ZN(n6954) );
  AOI22D1BWP30P140LVT U10179 ( .A1(i_data_bus[698]), .A2(n10404), .B1(
        i_data_bus[666]), .B2(n10401), .ZN(n6953) );
  ND2D1BWP30P140LVT U10180 ( .A1(n6954), .A2(n6953), .ZN(N14795) );
  AOI22D1BWP30P140LVT U10181 ( .A1(i_data_bus[718]), .A2(n10402), .B1(
        i_data_bus[750]), .B2(n10403), .ZN(n6956) );
  AOI22D1BWP30P140LVT U10182 ( .A1(i_data_bus[686]), .A2(n10404), .B1(
        i_data_bus[654]), .B2(n10401), .ZN(n6955) );
  ND2D1BWP30P140LVT U10183 ( .A1(n6956), .A2(n6955), .ZN(N14783) );
  AOI22D1BWP30P140LVT U10184 ( .A1(i_data_bus[714]), .A2(n10402), .B1(
        i_data_bus[682]), .B2(n10404), .ZN(n6958) );
  AOI22D1BWP30P140LVT U10185 ( .A1(i_data_bus[746]), .A2(n10403), .B1(
        i_data_bus[650]), .B2(n10401), .ZN(n6957) );
  ND2D1BWP30P140LVT U10186 ( .A1(n6958), .A2(n6957), .ZN(N14779) );
  AOI22D1BWP30P140LVT U10187 ( .A1(i_data_bus[717]), .A2(n10402), .B1(
        i_data_bus[685]), .B2(n10404), .ZN(n6960) );
  AOI22D1BWP30P140LVT U10188 ( .A1(i_data_bus[749]), .A2(n10403), .B1(
        i_data_bus[653]), .B2(n10401), .ZN(n6959) );
  ND2D1BWP30P140LVT U10189 ( .A1(n6960), .A2(n6959), .ZN(N14782) );
  AOI22D1BWP30P140LVT U10190 ( .A1(i_data_bus[694]), .A2(n10404), .B1(
        i_data_bus[726]), .B2(n10402), .ZN(n6962) );
  AOI22D1BWP30P140LVT U10191 ( .A1(i_data_bus[758]), .A2(n10403), .B1(
        i_data_bus[662]), .B2(n10401), .ZN(n6961) );
  ND2D1BWP30P140LVT U10192 ( .A1(n6962), .A2(n6961), .ZN(N14791) );
  AOI22D1BWP30P140LVT U10193 ( .A1(i_data_bus[674]), .A2(n10404), .B1(
        i_data_bus[738]), .B2(n10403), .ZN(n6964) );
  AOI22D1BWP30P140LVT U10194 ( .A1(i_data_bus[706]), .A2(n10402), .B1(
        i_data_bus[642]), .B2(n10401), .ZN(n6963) );
  ND2D1BWP30P140LVT U10195 ( .A1(n6964), .A2(n6963), .ZN(N14771) );
  AOI22D1BWP30P140LVT U10196 ( .A1(i_data_bus[757]), .A2(n10403), .B1(
        i_data_bus[693]), .B2(n10404), .ZN(n6966) );
  AOI22D1BWP30P140LVT U10197 ( .A1(i_data_bus[725]), .A2(n10402), .B1(
        i_data_bus[661]), .B2(n10401), .ZN(n6965) );
  ND2D1BWP30P140LVT U10198 ( .A1(n6966), .A2(n6965), .ZN(N14790) );
  AOI22D1BWP30P140LVT U10199 ( .A1(i_data_bus[747]), .A2(n10403), .B1(
        i_data_bus[683]), .B2(n10404), .ZN(n6968) );
  AOI22D1BWP30P140LVT U10200 ( .A1(i_data_bus[715]), .A2(n10402), .B1(
        i_data_bus[651]), .B2(n10401), .ZN(n6967) );
  ND2D1BWP30P140LVT U10201 ( .A1(n6968), .A2(n6967), .ZN(N14780) );
  AOI22D1BWP30P140LVT U10202 ( .A1(i_data_bus[155]), .A2(n10612), .B1(
        i_data_bus[251]), .B2(n10611), .ZN(n6970) );
  AOI22D1BWP30P140LVT U10203 ( .A1(i_data_bus[187]), .A2(n10609), .B1(
        i_data_bus[219]), .B2(n10610), .ZN(n6969) );
  ND2D1BWP30P140LVT U10204 ( .A1(n6970), .A2(n6969), .ZN(N2688) );
  AOI22D1BWP30P140LVT U10205 ( .A1(i_data_bus[179]), .A2(n10609), .B1(
        i_data_bus[243]), .B2(n10611), .ZN(n6972) );
  AOI22D1BWP30P140LVT U10206 ( .A1(i_data_bus[147]), .A2(n10612), .B1(
        i_data_bus[211]), .B2(n10610), .ZN(n6971) );
  ND2D1BWP30P140LVT U10207 ( .A1(n6972), .A2(n6971), .ZN(N2680) );
  AOI22D1BWP30P140LVT U10208 ( .A1(i_data_bus[146]), .A2(n10612), .B1(
        i_data_bus[242]), .B2(n10611), .ZN(n6974) );
  AOI22D1BWP30P140LVT U10209 ( .A1(i_data_bus[178]), .A2(n10609), .B1(
        i_data_bus[210]), .B2(n10610), .ZN(n6973) );
  ND2D1BWP30P140LVT U10210 ( .A1(n6974), .A2(n6973), .ZN(N2679) );
  AOI22D1BWP30P140LVT U10211 ( .A1(i_data_bus[148]), .A2(n10612), .B1(
        i_data_bus[244]), .B2(n10611), .ZN(n6976) );
  AOI22D1BWP30P140LVT U10212 ( .A1(i_data_bus[180]), .A2(n10609), .B1(
        i_data_bus[212]), .B2(n10610), .ZN(n6975) );
  ND2D1BWP30P140LVT U10213 ( .A1(n6976), .A2(n6975), .ZN(N2681) );
  AOI22D1BWP30P140LVT U10214 ( .A1(i_data_bus[177]), .A2(n10609), .B1(
        i_data_bus[241]), .B2(n10611), .ZN(n6978) );
  AOI22D1BWP30P140LVT U10215 ( .A1(i_data_bus[209]), .A2(n10610), .B1(
        i_data_bus[145]), .B2(n10612), .ZN(n6977) );
  ND2D1BWP30P140LVT U10216 ( .A1(n6978), .A2(n6977), .ZN(N2678) );
  AOI22D1BWP30P140LVT U10217 ( .A1(i_data_bus[193]), .A2(n10610), .B1(
        i_data_bus[225]), .B2(n10611), .ZN(n6980) );
  AOI22D1BWP30P140LVT U10218 ( .A1(i_data_bus[161]), .A2(n10609), .B1(
        i_data_bus[129]), .B2(n10612), .ZN(n6979) );
  ND2D1BWP30P140LVT U10219 ( .A1(n6980), .A2(n6979), .ZN(N2662) );
  AOI22D1BWP30P140LVT U10220 ( .A1(i_data_bus[129]), .A2(n10513), .B1(
        i_data_bus[225]), .B2(n10516), .ZN(n6982) );
  AOI22D1BWP30P140LVT U10221 ( .A1(i_data_bus[161]), .A2(n10515), .B1(
        i_data_bus[193]), .B2(n10514), .ZN(n6981) );
  ND2D1BWP30P140LVT U10222 ( .A1(n6982), .A2(n6981), .ZN(N8284) );
  AOI22D1BWP30P140LVT U10223 ( .A1(i_data_bus[183]), .A2(n10515), .B1(
        i_data_bus[247]), .B2(n10516), .ZN(n6984) );
  AOI22D1BWP30P140LVT U10224 ( .A1(i_data_bus[151]), .A2(n10513), .B1(
        i_data_bus[215]), .B2(n10514), .ZN(n6983) );
  ND2D1BWP30P140LVT U10225 ( .A1(n6984), .A2(n6983), .ZN(N8306) );
  AOI22D1BWP30P140LVT U10226 ( .A1(i_data_bus[201]), .A2(n10514), .B1(
        i_data_bus[233]), .B2(n10516), .ZN(n6986) );
  AOI22D1BWP30P140LVT U10227 ( .A1(i_data_bus[137]), .A2(n10513), .B1(
        i_data_bus[169]), .B2(n10515), .ZN(n6985) );
  ND2D1BWP30P140LVT U10228 ( .A1(n6986), .A2(n6985), .ZN(N8292) );
  AOI22D1BWP30P140LVT U10229 ( .A1(i_data_bus[156]), .A2(n10513), .B1(
        i_data_bus[252]), .B2(n10516), .ZN(n6988) );
  AOI22D1BWP30P140LVT U10230 ( .A1(i_data_bus[220]), .A2(n10514), .B1(
        i_data_bus[188]), .B2(n10515), .ZN(n6987) );
  ND2D1BWP30P140LVT U10231 ( .A1(n6988), .A2(n6987), .ZN(N8311) );
  AOI22D1BWP30P140LVT U10232 ( .A1(i_data_bus[212]), .A2(n10514), .B1(
        i_data_bus[244]), .B2(n10516), .ZN(n6990) );
  AOI22D1BWP30P140LVT U10233 ( .A1(i_data_bus[148]), .A2(n10513), .B1(
        i_data_bus[180]), .B2(n10515), .ZN(n6989) );
  ND2D1BWP30P140LVT U10234 ( .A1(n6990), .A2(n6989), .ZN(N8303) );
  AOI22D1BWP30P140LVT U10235 ( .A1(i_data_bus[1008]), .A2(n10393), .B1(
        i_data_bus[912]), .B2(n10395), .ZN(n6992) );
  AOI22D1BWP30P140LVT U10236 ( .A1(i_data_bus[976]), .A2(n10396), .B1(
        i_data_bus[944]), .B2(n10394), .ZN(n6991) );
  ND2D1BWP30P140LVT U10237 ( .A1(n6992), .A2(n6991), .ZN(N15217) );
  AOI22D1BWP30P140LVT U10238 ( .A1(i_data_bus[925]), .A2(n10395), .B1(
        i_data_bus[1021]), .B2(n10393), .ZN(n6994) );
  AOI22D1BWP30P140LVT U10239 ( .A1(i_data_bus[989]), .A2(n10396), .B1(
        i_data_bus[957]), .B2(n10394), .ZN(n6993) );
  ND2D1BWP30P140LVT U10240 ( .A1(n6994), .A2(n6993), .ZN(N15230) );
  AOI22D1BWP30P140LVT U10241 ( .A1(i_data_bus[1000]), .A2(n10393), .B1(
        i_data_bus[904]), .B2(n10395), .ZN(n6996) );
  AOI22D1BWP30P140LVT U10242 ( .A1(i_data_bus[968]), .A2(n10396), .B1(
        i_data_bus[936]), .B2(n10394), .ZN(n6995) );
  ND2D1BWP30P140LVT U10243 ( .A1(n6996), .A2(n6995), .ZN(N15209) );
  AOI22D1BWP30P140LVT U10244 ( .A1(i_data_bus[898]), .A2(n10395), .B1(
        i_data_bus[994]), .B2(n10393), .ZN(n6998) );
  AOI22D1BWP30P140LVT U10245 ( .A1(i_data_bus[962]), .A2(n10396), .B1(
        i_data_bus[930]), .B2(n10394), .ZN(n6997) );
  ND2D1BWP30P140LVT U10246 ( .A1(n6998), .A2(n6997), .ZN(N15203) );
  AOI22D1BWP30P140LVT U10247 ( .A1(i_data_bus[997]), .A2(n10393), .B1(
        i_data_bus[901]), .B2(n10395), .ZN(n7000) );
  AOI22D1BWP30P140LVT U10248 ( .A1(i_data_bus[965]), .A2(n10396), .B1(
        i_data_bus[933]), .B2(n10394), .ZN(n6999) );
  ND2D1BWP30P140LVT U10249 ( .A1(n7000), .A2(n6999), .ZN(N15206) );
  AOI22D1BWP30P140LVT U10250 ( .A1(i_data_bus[973]), .A2(n10396), .B1(
        i_data_bus[909]), .B2(n10395), .ZN(n7002) );
  AOI22D1BWP30P140LVT U10251 ( .A1(i_data_bus[1005]), .A2(n10393), .B1(
        i_data_bus[941]), .B2(n10394), .ZN(n7001) );
  ND2D1BWP30P140LVT U10252 ( .A1(n7002), .A2(n7001), .ZN(N15214) );
  AOI22D1BWP30P140LVT U10253 ( .A1(i_data_bus[1001]), .A2(n10393), .B1(
        i_data_bus[905]), .B2(n10395), .ZN(n7004) );
  AOI22D1BWP30P140LVT U10254 ( .A1(i_data_bus[969]), .A2(n10396), .B1(
        i_data_bus[937]), .B2(n10394), .ZN(n7003) );
  ND2D1BWP30P140LVT U10255 ( .A1(n7004), .A2(n7003), .ZN(N15210) );
  AOI22D1BWP30P140LVT U10256 ( .A1(i_data_bus[820]), .A2(n10496), .B1(
        i_data_bus[884]), .B2(n10494), .ZN(n7006) );
  AOI22D1BWP30P140LVT U10257 ( .A1(i_data_bus[788]), .A2(n10493), .B1(
        i_data_bus[852]), .B2(n10495), .ZN(n7005) );
  ND2D1BWP30P140LVT U10258 ( .A1(n7006), .A2(n7005), .ZN(N9383) );
  AOI22D1BWP30P140LVT U10259 ( .A1(i_data_bus[822]), .A2(n10496), .B1(
        i_data_bus[886]), .B2(n10494), .ZN(n7008) );
  AOI22D1BWP30P140LVT U10260 ( .A1(i_data_bus[790]), .A2(n10493), .B1(
        i_data_bus[854]), .B2(n10495), .ZN(n7007) );
  ND2D1BWP30P140LVT U10261 ( .A1(n7008), .A2(n7007), .ZN(N9385) );
  AOI22D1BWP30P140LVT U10262 ( .A1(i_data_bus[865]), .A2(n10494), .B1(
        i_data_bus[769]), .B2(n10493), .ZN(n7010) );
  AOI22D1BWP30P140LVT U10263 ( .A1(i_data_bus[801]), .A2(n10496), .B1(
        i_data_bus[833]), .B2(n10495), .ZN(n7009) );
  ND2D1BWP30P140LVT U10264 ( .A1(n7010), .A2(n7009), .ZN(N9364) );
  AOI22D1BWP30P140LVT U10265 ( .A1(i_data_bus[827]), .A2(n10496), .B1(
        i_data_bus[891]), .B2(n10494), .ZN(n7012) );
  AOI22D1BWP30P140LVT U10266 ( .A1(i_data_bus[795]), .A2(n10493), .B1(
        i_data_bus[859]), .B2(n10495), .ZN(n7011) );
  ND2D1BWP30P140LVT U10267 ( .A1(n7012), .A2(n7011), .ZN(N9390) );
  AOI22D1BWP30P140LVT U10268 ( .A1(i_data_bus[878]), .A2(n10494), .B1(
        i_data_bus[782]), .B2(n10493), .ZN(n7014) );
  AOI22D1BWP30P140LVT U10269 ( .A1(i_data_bus[814]), .A2(n10496), .B1(
        i_data_bus[846]), .B2(n10495), .ZN(n7013) );
  ND2D1BWP30P140LVT U10270 ( .A1(n7014), .A2(n7013), .ZN(N9377) );
  AOI22D1BWP30P140LVT U10271 ( .A1(i_data_bus[805]), .A2(n10496), .B1(
        i_data_bus[773]), .B2(n10493), .ZN(n7016) );
  AOI22D1BWP30P140LVT U10272 ( .A1(i_data_bus[869]), .A2(n10494), .B1(
        i_data_bus[837]), .B2(n10495), .ZN(n7015) );
  ND2D1BWP30P140LVT U10273 ( .A1(n7016), .A2(n7015), .ZN(N9368) );
  AOI22D1BWP30P140LVT U10274 ( .A1(i_data_bus[198]), .A2(n10548), .B1(
        i_data_bus[134]), .B2(n10546), .ZN(n7018) );
  AOI22D1BWP30P140LVT U10275 ( .A1(i_data_bus[230]), .A2(n10547), .B1(
        i_data_bus[166]), .B2(n10545), .ZN(n7017) );
  ND2D1BWP30P140LVT U10276 ( .A1(n7018), .A2(n7017), .ZN(N6415) );
  AOI22D1BWP30P140LVT U10277 ( .A1(i_data_bus[870]), .A2(n10431), .B1(
        i_data_bus[806]), .B2(n10430), .ZN(n7020) );
  AOI22D1BWP30P140LVT U10278 ( .A1(i_data_bus[838]), .A2(n10432), .B1(
        i_data_bus[774]), .B2(n10429), .ZN(n7019) );
  ND2D1BWP30P140LVT U10279 ( .A1(n7020), .A2(n7019), .ZN(N13117) );
  AOI22D1BWP30P140LVT U10280 ( .A1(i_data_bus[872]), .A2(n10431), .B1(
        i_data_bus[808]), .B2(n10430), .ZN(n7022) );
  AOI22D1BWP30P140LVT U10281 ( .A1(i_data_bus[840]), .A2(n10432), .B1(
        i_data_bus[776]), .B2(n10429), .ZN(n7021) );
  ND2D1BWP30P140LVT U10282 ( .A1(n7022), .A2(n7021), .ZN(N13119) );
  AOI22D1BWP30P140LVT U10283 ( .A1(i_data_bus[801]), .A2(n10430), .B1(
        i_data_bus[833]), .B2(n10432), .ZN(n7024) );
  AOI22D1BWP30P140LVT U10284 ( .A1(i_data_bus[865]), .A2(n10431), .B1(
        i_data_bus[769]), .B2(n10429), .ZN(n7023) );
  ND2D1BWP30P140LVT U10285 ( .A1(n7024), .A2(n7023), .ZN(N13112) );
  AOI22D1BWP30P140LVT U10286 ( .A1(i_data_bus[884]), .A2(n10431), .B1(
        i_data_bus[852]), .B2(n10432), .ZN(n7026) );
  AOI22D1BWP30P140LVT U10287 ( .A1(i_data_bus[820]), .A2(n10430), .B1(
        i_data_bus[788]), .B2(n10429), .ZN(n7025) );
  ND2D1BWP30P140LVT U10288 ( .A1(n7026), .A2(n7025), .ZN(N13131) );
  AOI22D1BWP30P140LVT U10289 ( .A1(i_data_bus[886]), .A2(n10431), .B1(
        i_data_bus[854]), .B2(n10432), .ZN(n7028) );
  AOI22D1BWP30P140LVT U10290 ( .A1(i_data_bus[822]), .A2(n10430), .B1(
        i_data_bus[790]), .B2(n10429), .ZN(n7027) );
  ND2D1BWP30P140LVT U10291 ( .A1(n7028), .A2(n7027), .ZN(N13133) );
  AOI22D1BWP30P140LVT U10292 ( .A1(i_data_bus[871]), .A2(n10431), .B1(
        i_data_bus[839]), .B2(n10432), .ZN(n7030) );
  AOI22D1BWP30P140LVT U10293 ( .A1(i_data_bus[807]), .A2(n10430), .B1(
        i_data_bus[775]), .B2(n10429), .ZN(n7029) );
  ND2D1BWP30P140LVT U10294 ( .A1(n7030), .A2(n7029), .ZN(N13118) );
  AOI22D1BWP30P140LVT U10295 ( .A1(i_data_bus[894]), .A2(n10431), .B1(
        i_data_bus[830]), .B2(n10430), .ZN(n7032) );
  AOI22D1BWP30P140LVT U10296 ( .A1(i_data_bus[862]), .A2(n10432), .B1(
        i_data_bus[798]), .B2(n10429), .ZN(n7031) );
  ND2D1BWP30P140LVT U10297 ( .A1(n7032), .A2(n7031), .ZN(N13141) );
  AOI22D1BWP30P140LVT U10298 ( .A1(i_data_bus[878]), .A2(n10431), .B1(
        i_data_bus[846]), .B2(n10432), .ZN(n7034) );
  AOI22D1BWP30P140LVT U10299 ( .A1(i_data_bus[814]), .A2(n10430), .B1(
        i_data_bus[782]), .B2(n10429), .ZN(n7033) );
  ND2D1BWP30P140LVT U10300 ( .A1(n7034), .A2(n7033), .ZN(N13125) );
  AOI22D1BWP30P140LVT U10301 ( .A1(i_data_bus[819]), .A2(n10430), .B1(
        i_data_bus[851]), .B2(n10432), .ZN(n7036) );
  AOI22D1BWP30P140LVT U10302 ( .A1(i_data_bus[883]), .A2(n10431), .B1(
        i_data_bus[787]), .B2(n10429), .ZN(n7035) );
  ND2D1BWP30P140LVT U10303 ( .A1(n7036), .A2(n7035), .ZN(N13130) );
  NR4D1BWP30P140LVT U10304 ( .A1(i_cmd[142]), .A2(n7039), .A3(n9837), .A4(
        n7037), .ZN(n10440) );
  INR4D1BWP30P140LVT U10305 ( .A1(i_cmd[134]), .B1(i_cmd[150]), .B2(n9839), 
        .B3(n7040), .ZN(n10438) );
  AOI22D1BWP30P140LVT U10306 ( .A1(i_data_bus[630]), .A2(n10440), .B1(
        i_data_bus[534]), .B2(n10438), .ZN(n7042) );
  NR4D1BWP30P140LVT U10307 ( .A1(i_cmd[158]), .A2(n7039), .A3(n9833), .A4(
        n7038), .ZN(n10439) );
  INR4D1BWP30P140LVT U10308 ( .A1(i_cmd[150]), .B1(i_cmd[134]), .B2(n9834), 
        .B3(n7040), .ZN(n10437) );
  AOI22D1BWP30P140LVT U10309 ( .A1(i_data_bus[566]), .A2(n10439), .B1(
        i_data_bus[598]), .B2(n10437), .ZN(n7041) );
  ND2D1BWP30P140LVT U10310 ( .A1(n7042), .A2(n7041), .ZN(N12701) );
  AOI22D1BWP30P140LVT U10311 ( .A1(i_data_bus[617]), .A2(n10440), .B1(
        i_data_bus[553]), .B2(n10439), .ZN(n7044) );
  AOI22D1BWP30P140LVT U10312 ( .A1(i_data_bus[521]), .A2(n10438), .B1(
        i_data_bus[585]), .B2(n10437), .ZN(n7043) );
  ND2D1BWP30P140LVT U10313 ( .A1(n7044), .A2(n7043), .ZN(N12688) );
  AOI22D1BWP30P140LVT U10314 ( .A1(i_data_bus[635]), .A2(n10440), .B1(
        i_data_bus[539]), .B2(n10438), .ZN(n7046) );
  AOI22D1BWP30P140LVT U10315 ( .A1(i_data_bus[571]), .A2(n10439), .B1(
        i_data_bus[603]), .B2(n10437), .ZN(n7045) );
  ND2D1BWP30P140LVT U10316 ( .A1(n7046), .A2(n7045), .ZN(N12706) );
  AOI22D1BWP30P140LVT U10317 ( .A1(i_data_bus[638]), .A2(n10440), .B1(
        i_data_bus[574]), .B2(n10439), .ZN(n7048) );
  AOI22D1BWP30P140LVT U10318 ( .A1(i_data_bus[542]), .A2(n10438), .B1(
        i_data_bus[606]), .B2(n10437), .ZN(n7047) );
  ND2D1BWP30P140LVT U10319 ( .A1(n7048), .A2(n7047), .ZN(N12709) );
  AOI22D1BWP30P140LVT U10320 ( .A1(i_data_bus[618]), .A2(n10440), .B1(
        i_data_bus[522]), .B2(n10438), .ZN(n7050) );
  AOI22D1BWP30P140LVT U10321 ( .A1(i_data_bus[554]), .A2(n10439), .B1(
        i_data_bus[586]), .B2(n10437), .ZN(n7049) );
  ND2D1BWP30P140LVT U10322 ( .A1(n7050), .A2(n7049), .ZN(N12689) );
  AOI22D1BWP30P140LVT U10323 ( .A1(i_data_bus[292]), .A2(n10573), .B1(
        i_data_bus[356]), .B2(n10574), .ZN(n7052) );
  AOI22D1BWP30P140LVT U10324 ( .A1(i_data_bus[324]), .A2(n10576), .B1(
        i_data_bus[260]), .B2(n10575), .ZN(n7051) );
  ND2D1BWP30P140LVT U10325 ( .A1(n7052), .A2(n7051), .ZN(N4755) );
  AOI22D1BWP30P140LVT U10326 ( .A1(i_data_bus[298]), .A2(n10573), .B1(
        i_data_bus[362]), .B2(n10574), .ZN(n7054) );
  AOI22D1BWP30P140LVT U10327 ( .A1(i_data_bus[266]), .A2(n10575), .B1(
        i_data_bus[330]), .B2(n10576), .ZN(n7053) );
  ND2D1BWP30P140LVT U10328 ( .A1(n7054), .A2(n7053), .ZN(N4761) );
  AOI22D1BWP30P140LVT U10329 ( .A1(i_data_bus[349]), .A2(n10576), .B1(
        i_data_bus[381]), .B2(n10574), .ZN(n7056) );
  AOI22D1BWP30P140LVT U10330 ( .A1(i_data_bus[317]), .A2(n10573), .B1(
        i_data_bus[285]), .B2(n10575), .ZN(n7055) );
  ND2D1BWP30P140LVT U10331 ( .A1(n7056), .A2(n7055), .ZN(N4780) );
  AOI22D1BWP30P140LVT U10332 ( .A1(i_data_bus[327]), .A2(n10576), .B1(
        i_data_bus[359]), .B2(n10574), .ZN(n7058) );
  AOI22D1BWP30P140LVT U10333 ( .A1(i_data_bus[295]), .A2(n10573), .B1(
        i_data_bus[263]), .B2(n10575), .ZN(n7057) );
  ND2D1BWP30P140LVT U10334 ( .A1(n7058), .A2(n7057), .ZN(N4758) );
  AOI22D1BWP30P140LVT U10335 ( .A1(i_data_bus[436]), .A2(n10443), .B1(
        i_data_bus[500]), .B2(n10444), .ZN(n7060) );
  AOI22D1BWP30P140LVT U10336 ( .A1(i_data_bus[404]), .A2(n10441), .B1(
        i_data_bus[468]), .B2(n10442), .ZN(n7059) );
  ND2D1BWP30P140LVT U10337 ( .A1(n7060), .A2(n7059), .ZN(N12483) );
  AOI22D1BWP30P140LVT U10338 ( .A1(i_data_bus[397]), .A2(n10441), .B1(
        i_data_bus[493]), .B2(n10444), .ZN(n7062) );
  AOI22D1BWP30P140LVT U10339 ( .A1(i_data_bus[429]), .A2(n10443), .B1(
        i_data_bus[461]), .B2(n10442), .ZN(n7061) );
  ND2D1BWP30P140LVT U10340 ( .A1(n7062), .A2(n7061), .ZN(N12476) );
  AOI22D1BWP30P140LVT U10341 ( .A1(i_data_bus[495]), .A2(n10444), .B1(
        i_data_bus[399]), .B2(n10441), .ZN(n7064) );
  AOI22D1BWP30P140LVT U10342 ( .A1(i_data_bus[431]), .A2(n10443), .B1(
        i_data_bus[463]), .B2(n10442), .ZN(n7063) );
  ND2D1BWP30P140LVT U10343 ( .A1(n7064), .A2(n7063), .ZN(N12478) );
  AOI22D1BWP30P140LVT U10344 ( .A1(i_data_bus[434]), .A2(n10443), .B1(
        i_data_bus[402]), .B2(n10441), .ZN(n7066) );
  AOI22D1BWP30P140LVT U10345 ( .A1(i_data_bus[498]), .A2(n10444), .B1(
        i_data_bus[466]), .B2(n10442), .ZN(n7065) );
  ND2D1BWP30P140LVT U10346 ( .A1(n7066), .A2(n7065), .ZN(N12481) );
  AOI22D1BWP30P140LVT U10347 ( .A1(i_data_bus[508]), .A2(n10444), .B1(
        i_data_bus[412]), .B2(n10441), .ZN(n7068) );
  AOI22D1BWP30P140LVT U10348 ( .A1(i_data_bus[444]), .A2(n10443), .B1(
        i_data_bus[476]), .B2(n10442), .ZN(n7067) );
  ND2D1BWP30P140LVT U10349 ( .A1(n7068), .A2(n7067), .ZN(N12491) );
  AOI22D1BWP30P140LVT U10350 ( .A1(i_data_bus[414]), .A2(n10441), .B1(
        i_data_bus[510]), .B2(n10444), .ZN(n7070) );
  AOI22D1BWP30P140LVT U10351 ( .A1(i_data_bus[446]), .A2(n10443), .B1(
        i_data_bus[478]), .B2(n10442), .ZN(n7069) );
  ND2D1BWP30P140LVT U10352 ( .A1(n7070), .A2(n7069), .ZN(N12493) );
  AOI22D1BWP30P140LVT U10353 ( .A1(i_data_bus[509]), .A2(n10444), .B1(
        i_data_bus[445]), .B2(n10443), .ZN(n7072) );
  AOI22D1BWP30P140LVT U10354 ( .A1(i_data_bus[413]), .A2(n10441), .B1(
        i_data_bus[477]), .B2(n10442), .ZN(n7071) );
  ND2D1BWP30P140LVT U10355 ( .A1(n7072), .A2(n7071), .ZN(N12492) );
  AOI22D1BWP30P140LVT U10356 ( .A1(i_data_bus[437]), .A2(n10443), .B1(
        i_data_bus[501]), .B2(n10444), .ZN(n7074) );
  AOI22D1BWP30P140LVT U10357 ( .A1(i_data_bus[405]), .A2(n10441), .B1(
        i_data_bus[469]), .B2(n10442), .ZN(n7073) );
  ND2D1BWP30P140LVT U10358 ( .A1(n7074), .A2(n7073), .ZN(N12484) );
  AOI22D1BWP30P140LVT U10359 ( .A1(i_data_bus[410]), .A2(n10441), .B1(
        i_data_bus[442]), .B2(n10443), .ZN(n7076) );
  AOI22D1BWP30P140LVT U10360 ( .A1(i_data_bus[506]), .A2(n10444), .B1(
        i_data_bus[474]), .B2(n10442), .ZN(n7075) );
  ND2D1BWP30P140LVT U10361 ( .A1(n7076), .A2(n7075), .ZN(N12489) );
  AOI22D1BWP30P140LVT U10362 ( .A1(i_data_bus[315]), .A2(n10448), .B1(
        i_data_bus[347]), .B2(n10446), .ZN(n7078) );
  AOI22D1BWP30P140LVT U10363 ( .A1(i_data_bus[379]), .A2(n10445), .B1(
        i_data_bus[283]), .B2(n10447), .ZN(n7077) );
  ND2D1BWP30P140LVT U10364 ( .A1(n7078), .A2(n7077), .ZN(N12274) );
  AOI22D1BWP30P140LVT U10365 ( .A1(i_data_bus[357]), .A2(n10445), .B1(
        i_data_bus[293]), .B2(n10448), .ZN(n7080) );
  AOI22D1BWP30P140LVT U10366 ( .A1(i_data_bus[325]), .A2(n10446), .B1(
        i_data_bus[261]), .B2(n10447), .ZN(n7079) );
  ND2D1BWP30P140LVT U10367 ( .A1(n7080), .A2(n7079), .ZN(N12252) );
  AOI22D1BWP30P140LVT U10368 ( .A1(i_data_bus[352]), .A2(n10445), .B1(
        i_data_bus[320]), .B2(n10446), .ZN(n7082) );
  AOI22D1BWP30P140LVT U10369 ( .A1(i_data_bus[288]), .A2(n10448), .B1(
        i_data_bus[256]), .B2(n10447), .ZN(n7081) );
  ND2D1BWP30P140LVT U10370 ( .A1(n7082), .A2(n7081), .ZN(N12247) );
  AOI22D1BWP30P140LVT U10371 ( .A1(i_data_bus[368]), .A2(n10445), .B1(
        i_data_bus[336]), .B2(n10446), .ZN(n7084) );
  AOI22D1BWP30P140LVT U10372 ( .A1(i_data_bus[304]), .A2(n10448), .B1(
        i_data_bus[272]), .B2(n10447), .ZN(n7083) );
  ND2D1BWP30P140LVT U10373 ( .A1(n7084), .A2(n7083), .ZN(N12263) );
  AOI22D1BWP30P140LVT U10374 ( .A1(i_data_bus[295]), .A2(n10448), .B1(
        i_data_bus[327]), .B2(n10446), .ZN(n7086) );
  AOI22D1BWP30P140LVT U10375 ( .A1(i_data_bus[359]), .A2(n10445), .B1(
        i_data_bus[263]), .B2(n10447), .ZN(n7085) );
  ND2D1BWP30P140LVT U10376 ( .A1(n7086), .A2(n7085), .ZN(N12254) );
  AOI22D1BWP30P140LVT U10377 ( .A1(i_data_bus[118]), .A2(n10616), .B1(
        i_data_bus[22]), .B2(n10615), .ZN(n7088) );
  AOI22D1BWP30P140LVT U10378 ( .A1(i_data_bus[86]), .A2(n10613), .B1(
        i_data_bus[54]), .B2(n10614), .ZN(n7087) );
  ND2D1BWP30P140LVT U10379 ( .A1(n7088), .A2(n7087), .ZN(N2467) );
  AOI22D1BWP30P140LVT U10380 ( .A1(i_data_bus[66]), .A2(n10613), .B1(
        i_data_bus[2]), .B2(n10615), .ZN(n7090) );
  AOI22D1BWP30P140LVT U10381 ( .A1(i_data_bus[98]), .A2(n10616), .B1(
        i_data_bus[34]), .B2(n10614), .ZN(n7089) );
  ND2D1BWP30P140LVT U10382 ( .A1(n7090), .A2(n7089), .ZN(N2447) );
  AOI22D1BWP30P140LVT U10383 ( .A1(i_data_bus[99]), .A2(n10616), .B1(
        i_data_bus[3]), .B2(n10615), .ZN(n7092) );
  AOI22D1BWP30P140LVT U10384 ( .A1(i_data_bus[67]), .A2(n10613), .B1(
        i_data_bus[35]), .B2(n10614), .ZN(n7091) );
  ND2D1BWP30P140LVT U10385 ( .A1(n7092), .A2(n7091), .ZN(N2448) );
  AOI22D1BWP30P140LVT U10386 ( .A1(i_data_bus[82]), .A2(n10613), .B1(
        i_data_bus[18]), .B2(n10615), .ZN(n7094) );
  AOI22D1BWP30P140LVT U10387 ( .A1(i_data_bus[114]), .A2(n10616), .B1(
        i_data_bus[50]), .B2(n10614), .ZN(n7093) );
  ND2D1BWP30P140LVT U10388 ( .A1(n7094), .A2(n7093), .ZN(N2463) );
  AOI22D1BWP30P140LVT U10389 ( .A1(i_data_bus[94]), .A2(n10613), .B1(
        i_data_bus[30]), .B2(n10615), .ZN(n7096) );
  AOI22D1BWP30P140LVT U10390 ( .A1(i_data_bus[126]), .A2(n10616), .B1(
        i_data_bus[62]), .B2(n10614), .ZN(n7095) );
  ND2D1BWP30P140LVT U10391 ( .A1(n7096), .A2(n7095), .ZN(N2475) );
  AOI22D1BWP30P140LVT U10392 ( .A1(i_data_bus[266]), .A2(n10447), .B1(
        i_data_bus[362]), .B2(n10445), .ZN(n7098) );
  AOI22D1BWP30P140LVT U10393 ( .A1(i_data_bus[330]), .A2(n10446), .B1(
        i_data_bus[298]), .B2(n10448), .ZN(n7097) );
  ND2D1BWP30P140LVT U10394 ( .A1(n7098), .A2(n7097), .ZN(N12257) );
  AOI22D1BWP30P140LVT U10395 ( .A1(i_data_bus[317]), .A2(n10448), .B1(
        i_data_bus[381]), .B2(n10445), .ZN(n7100) );
  AOI22D1BWP30P140LVT U10396 ( .A1(i_data_bus[349]), .A2(n10446), .B1(
        i_data_bus[285]), .B2(n10447), .ZN(n7099) );
  ND2D1BWP30P140LVT U10397 ( .A1(n7100), .A2(n7099), .ZN(N12276) );
  AOI22D1BWP30P140LVT U10398 ( .A1(i_data_bus[296]), .A2(n10448), .B1(
        i_data_bus[360]), .B2(n10445), .ZN(n7102) );
  AOI22D1BWP30P140LVT U10399 ( .A1(i_data_bus[328]), .A2(n10446), .B1(
        i_data_bus[264]), .B2(n10447), .ZN(n7101) );
  ND2D1BWP30P140LVT U10400 ( .A1(n7102), .A2(n7101), .ZN(N12255) );
  AOI22D1BWP30P140LVT U10401 ( .A1(i_data_bus[10]), .A2(n10456), .B1(
        i_data_bus[106]), .B2(n10455), .ZN(n7104) );
  AOI22D1BWP30P140LVT U10402 ( .A1(i_data_bus[74]), .A2(n10454), .B1(
        i_data_bus[42]), .B2(n10453), .ZN(n7103) );
  ND2D1BWP30P140LVT U10403 ( .A1(n7104), .A2(n7103), .ZN(N11825) );
  AOI22D1BWP30P140LVT U10404 ( .A1(i_data_bus[370]), .A2(n10479), .B1(
        i_data_bus[306]), .B2(n10477), .ZN(n7106) );
  AOI22D1BWP30P140LVT U10405 ( .A1(i_data_bus[338]), .A2(n10478), .B1(
        i_data_bus[274]), .B2(n10480), .ZN(n7105) );
  ND2D1BWP30P140LVT U10406 ( .A1(n7106), .A2(n7105), .ZN(N10391) );
  AOI22D1BWP30P140LVT U10407 ( .A1(i_data_bus[368]), .A2(n10479), .B1(
        i_data_bus[304]), .B2(n10477), .ZN(n7108) );
  AOI22D1BWP30P140LVT U10408 ( .A1(i_data_bus[336]), .A2(n10478), .B1(
        i_data_bus[272]), .B2(n10480), .ZN(n7107) );
  ND2D1BWP30P140LVT U10409 ( .A1(n7108), .A2(n7107), .ZN(N10389) );
  AOI22D1BWP30P140LVT U10410 ( .A1(i_data_bus[288]), .A2(n10477), .B1(
        i_data_bus[320]), .B2(n10478), .ZN(n7110) );
  AOI22D1BWP30P140LVT U10411 ( .A1(i_data_bus[352]), .A2(n10479), .B1(
        i_data_bus[256]), .B2(n10480), .ZN(n7109) );
  ND2D1BWP30P140LVT U10412 ( .A1(n7110), .A2(n7109), .ZN(N10373) );
  AOI22D1BWP30P140LVT U10413 ( .A1(i_data_bus[100]), .A2(n10455), .B1(
        i_data_bus[68]), .B2(n10454), .ZN(n7112) );
  AOI22D1BWP30P140LVT U10414 ( .A1(i_data_bus[4]), .A2(n10456), .B1(
        i_data_bus[36]), .B2(n10453), .ZN(n7111) );
  ND2D1BWP30P140LVT U10415 ( .A1(n7112), .A2(n7111), .ZN(N11819) );
  AOI22D1BWP30P140LVT U10416 ( .A1(i_data_bus[95]), .A2(n10454), .B1(
        i_data_bus[127]), .B2(n10455), .ZN(n7114) );
  AOI22D1BWP30P140LVT U10417 ( .A1(i_data_bus[31]), .A2(n10456), .B1(
        i_data_bus[63]), .B2(n10453), .ZN(n7113) );
  ND2D1BWP30P140LVT U10418 ( .A1(n7114), .A2(n7113), .ZN(N11846) );
  AOI22D1BWP30P140LVT U10419 ( .A1(i_data_bus[73]), .A2(n10454), .B1(
        i_data_bus[105]), .B2(n10455), .ZN(n7116) );
  AOI22D1BWP30P140LVT U10420 ( .A1(i_data_bus[9]), .A2(n10456), .B1(
        i_data_bus[41]), .B2(n10453), .ZN(n7115) );
  ND2D1BWP30P140LVT U10421 ( .A1(n7116), .A2(n7115), .ZN(N11824) );
  AOI22D1BWP30P140LVT U10422 ( .A1(i_data_bus[136]), .A2(n10577), .B1(
        i_data_bus[232]), .B2(n10580), .ZN(n7118) );
  AOI22D1BWP30P140LVT U10423 ( .A1(i_data_bus[200]), .A2(n10578), .B1(
        i_data_bus[168]), .B2(n10579), .ZN(n7117) );
  ND2D1BWP30P140LVT U10424 ( .A1(n7118), .A2(n7117), .ZN(N4543) );
  AOI22D1BWP30P140LVT U10425 ( .A1(i_data_bus[212]), .A2(n10578), .B1(
        i_data_bus[244]), .B2(n10580), .ZN(n7120) );
  AOI22D1BWP30P140LVT U10426 ( .A1(i_data_bus[148]), .A2(n10577), .B1(
        i_data_bus[180]), .B2(n10579), .ZN(n7119) );
  ND2D1BWP30P140LVT U10427 ( .A1(n7120), .A2(n7119), .ZN(N4555) );
  AOI22D1BWP30P140LVT U10428 ( .A1(i_data_bus[132]), .A2(n10577), .B1(
        i_data_bus[196]), .B2(n10578), .ZN(n7122) );
  AOI22D1BWP30P140LVT U10429 ( .A1(i_data_bus[228]), .A2(n10580), .B1(
        i_data_bus[164]), .B2(n10579), .ZN(n7121) );
  ND2D1BWP30P140LVT U10430 ( .A1(n7122), .A2(n7121), .ZN(N4539) );
  AOI22D1BWP30P140LVT U10431 ( .A1(i_data_bus[128]), .A2(n10577), .B1(
        i_data_bus[192]), .B2(n10578), .ZN(n7124) );
  AOI22D1BWP30P140LVT U10432 ( .A1(i_data_bus[224]), .A2(n10580), .B1(
        i_data_bus[160]), .B2(n10579), .ZN(n7123) );
  ND2D1BWP30P140LVT U10433 ( .A1(n7124), .A2(n7123), .ZN(N4535) );
  NR4D1BWP30P140LVT U10434 ( .A1(i_cmd[234]), .A2(n7128), .A3(n10030), .A4(
        n7125), .ZN(n10556) );
  INR4D1BWP30P140LVT U10435 ( .A1(i_cmd[226]), .B1(i_cmd[242]), .B2(n10028), 
        .B3(n7126), .ZN(n10554) );
  AOI22D1BWP30P140LVT U10436 ( .A1(i_data_bus[1012]), .A2(n10556), .B1(
        i_data_bus[916]), .B2(n10554), .ZN(n7130) );
  INR4D1BWP30P140LVT U10437 ( .A1(i_cmd[242]), .B1(i_cmd[226]), .B2(n10024), 
        .B3(n7126), .ZN(n10555) );
  NR4D1BWP30P140LVT U10438 ( .A1(i_cmd[250]), .A2(n7128), .A3(n10023), .A4(
        n7127), .ZN(n10553) );
  AOI22D1BWP30P140LVT U10439 ( .A1(i_data_bus[980]), .A2(n10555), .B1(
        i_data_bus[948]), .B2(n10553), .ZN(n7129) );
  ND2D1BWP30P140LVT U10440 ( .A1(n7130), .A2(n7129), .ZN(N5851) );
  AOI22D1BWP30P140LVT U10441 ( .A1(i_data_bus[906]), .A2(n10554), .B1(
        i_data_bus[1002]), .B2(n10556), .ZN(n7132) );
  AOI22D1BWP30P140LVT U10442 ( .A1(i_data_bus[970]), .A2(n10555), .B1(
        i_data_bus[938]), .B2(n10553), .ZN(n7131) );
  ND2D1BWP30P140LVT U10443 ( .A1(n7132), .A2(n7131), .ZN(N5841) );
  AOI22D1BWP30P140LVT U10444 ( .A1(i_data_bus[917]), .A2(n10554), .B1(
        i_data_bus[1013]), .B2(n10556), .ZN(n7134) );
  AOI22D1BWP30P140LVT U10445 ( .A1(i_data_bus[981]), .A2(n10555), .B1(
        i_data_bus[949]), .B2(n10553), .ZN(n7133) );
  ND2D1BWP30P140LVT U10446 ( .A1(n7134), .A2(n7133), .ZN(N5852) );
  AOI22D1BWP30P140LVT U10447 ( .A1(i_data_bus[899]), .A2(n10554), .B1(
        i_data_bus[963]), .B2(n10555), .ZN(n7136) );
  AOI22D1BWP30P140LVT U10448 ( .A1(i_data_bus[995]), .A2(n10556), .B1(
        i_data_bus[931]), .B2(n10553), .ZN(n7135) );
  ND2D1BWP30P140LVT U10449 ( .A1(n7136), .A2(n7135), .ZN(N5834) );
  AOI22D1BWP30P140LVT U10450 ( .A1(i_data_bus[927]), .A2(n10554), .B1(
        i_data_bus[991]), .B2(n10555), .ZN(n7138) );
  AOI22D1BWP30P140LVT U10451 ( .A1(i_data_bus[1023]), .A2(n10556), .B1(
        i_data_bus[959]), .B2(n10553), .ZN(n7137) );
  ND2D1BWP30P140LVT U10452 ( .A1(n7138), .A2(n7137), .ZN(N5862) );
  AOI22D1BWP30P140LVT U10453 ( .A1(i_data_bus[967]), .A2(n10555), .B1(
        i_data_bus[999]), .B2(n10556), .ZN(n7140) );
  AOI22D1BWP30P140LVT U10454 ( .A1(i_data_bus[903]), .A2(n10554), .B1(
        i_data_bus[935]), .B2(n10553), .ZN(n7139) );
  ND2D1BWP30P140LVT U10455 ( .A1(n7140), .A2(n7139), .ZN(N5838) );
  AOI22D1BWP30P140LVT U10456 ( .A1(i_data_bus[982]), .A2(n10555), .B1(
        i_data_bus[918]), .B2(n10554), .ZN(n7142) );
  AOI22D1BWP30P140LVT U10457 ( .A1(i_data_bus[1014]), .A2(n10556), .B1(
        i_data_bus[950]), .B2(n10553), .ZN(n7141) );
  ND2D1BWP30P140LVT U10458 ( .A1(n7142), .A2(n7141), .ZN(N5853) );
  AOI22D1BWP30P140LVT U10459 ( .A1(i_data_bus[1008]), .A2(n10556), .B1(
        i_data_bus[976]), .B2(n10555), .ZN(n7144) );
  AOI22D1BWP30P140LVT U10460 ( .A1(i_data_bus[912]), .A2(n10554), .B1(
        i_data_bus[944]), .B2(n10553), .ZN(n7143) );
  ND2D1BWP30P140LVT U10461 ( .A1(n7144), .A2(n7143), .ZN(N5847) );
  AOI22D1BWP30P140LVT U10462 ( .A1(i_data_bus[913]), .A2(n10554), .B1(
        i_data_bus[977]), .B2(n10555), .ZN(n7146) );
  AOI22D1BWP30P140LVT U10463 ( .A1(i_data_bus[1009]), .A2(n10556), .B1(
        i_data_bus[945]), .B2(n10553), .ZN(n7145) );
  ND2D1BWP30P140LVT U10464 ( .A1(n7146), .A2(n7145), .ZN(N5848) );
  AOI22D1BWP30P140LVT U10465 ( .A1(i_data_bus[405]), .A2(n10473), .B1(
        i_data_bus[437]), .B2(n10474), .ZN(n7148) );
  AOI22D1BWP30P140LVT U10466 ( .A1(i_data_bus[469]), .A2(n10476), .B1(
        i_data_bus[501]), .B2(n10475), .ZN(n7147) );
  ND2D1BWP30P140LVT U10467 ( .A1(n7148), .A2(n7147), .ZN(N10610) );
  AOI22D1BWP30P140LVT U10468 ( .A1(i_data_bus[384]), .A2(n10473), .B1(
        i_data_bus[416]), .B2(n10474), .ZN(n7150) );
  AOI22D1BWP30P140LVT U10469 ( .A1(i_data_bus[448]), .A2(n10476), .B1(
        i_data_bus[480]), .B2(n10475), .ZN(n7149) );
  ND2D1BWP30P140LVT U10470 ( .A1(n7150), .A2(n7149), .ZN(N10589) );
  AOI22D1BWP30P140LVT U10471 ( .A1(i_data_bus[473]), .A2(n10476), .B1(
        i_data_bus[441]), .B2(n10474), .ZN(n7152) );
  AOI22D1BWP30P140LVT U10472 ( .A1(i_data_bus[409]), .A2(n10473), .B1(
        i_data_bus[505]), .B2(n10475), .ZN(n7151) );
  ND2D1BWP30P140LVT U10473 ( .A1(n7152), .A2(n7151), .ZN(N10614) );
  AOI22D1BWP30P140LVT U10474 ( .A1(i_data_bus[401]), .A2(n10473), .B1(
        i_data_bus[433]), .B2(n10474), .ZN(n7154) );
  AOI22D1BWP30P140LVT U10475 ( .A1(i_data_bus[465]), .A2(n10476), .B1(
        i_data_bus[497]), .B2(n10475), .ZN(n7153) );
  ND2D1BWP30P140LVT U10476 ( .A1(n7154), .A2(n7153), .ZN(N10606) );
  NR4D1BWP30P140LVT U10477 ( .A1(i_cmd[154]), .A2(n7157), .A3(n9833), .A4(
        n7155), .ZN(n10567) );
  INR4D1BWP30P140LVT U10478 ( .A1(i_cmd[130]), .B1(i_cmd[146]), .B2(n9839), 
        .B3(n7158), .ZN(n10566) );
  AOI22D1BWP30P140LVT U10479 ( .A1(i_data_bus[566]), .A2(n10567), .B1(
        i_data_bus[534]), .B2(n10566), .ZN(n7160) );
  NR4D1BWP30P140LVT U10480 ( .A1(i_cmd[138]), .A2(n7157), .A3(n9837), .A4(
        n7156), .ZN(n10568) );
  INR4D1BWP30P140LVT U10481 ( .A1(i_cmd[146]), .B1(i_cmd[130]), .B2(n9834), 
        .B3(n7158), .ZN(n10565) );
  AOI22D1BWP30P140LVT U10482 ( .A1(i_data_bus[630]), .A2(n10568), .B1(
        i_data_bus[598]), .B2(n10565), .ZN(n7159) );
  ND2D1BWP30P140LVT U10483 ( .A1(n7160), .A2(n7159), .ZN(N5205) );
  NR4D1BWP30P140LVT U10484 ( .A1(i_cmd[141]), .A2(n7161), .A3(n9837), .A4(
        n7163), .ZN(n10470) );
  NR4D1BWP30P140LVT U10485 ( .A1(i_cmd[157]), .A2(n7161), .A3(n9833), .A4(
        n7162), .ZN(n10472) );
  AOI22D1BWP30P140LVT U10486 ( .A1(i_data_bus[615]), .A2(n10470), .B1(
        i_data_bus[551]), .B2(n10472), .ZN(n7166) );
  INR4D1BWP30P140LVT U10487 ( .A1(i_cmd[133]), .B1(i_cmd[149]), .B2(n9839), 
        .B3(n7164), .ZN(n10471) );
  INR4D1BWP30P140LVT U10488 ( .A1(i_cmd[149]), .B1(i_cmd[133]), .B2(n9834), 
        .B3(n7164), .ZN(n10469) );
  AOI22D1BWP30P140LVT U10489 ( .A1(i_data_bus[519]), .A2(n10471), .B1(
        i_data_bus[583]), .B2(n10469), .ZN(n7165) );
  ND2D1BWP30P140LVT U10490 ( .A1(n7166), .A2(n7165), .ZN(N10812) );
  AOI22D1BWP30P140LVT U10491 ( .A1(i_data_bus[531]), .A2(n10566), .B1(
        i_data_bus[563]), .B2(n10567), .ZN(n7168) );
  AOI22D1BWP30P140LVT U10492 ( .A1(i_data_bus[627]), .A2(n10568), .B1(
        i_data_bus[595]), .B2(n10565), .ZN(n7167) );
  ND2D1BWP30P140LVT U10493 ( .A1(n7168), .A2(n7167), .ZN(N5202) );
  AOI22D1BWP30P140LVT U10494 ( .A1(i_data_bus[516]), .A2(n10566), .B1(
        i_data_bus[548]), .B2(n10567), .ZN(n7170) );
  AOI22D1BWP30P140LVT U10495 ( .A1(i_data_bus[612]), .A2(n10568), .B1(
        i_data_bus[580]), .B2(n10565), .ZN(n7169) );
  ND2D1BWP30P140LVT U10496 ( .A1(n7170), .A2(n7169), .ZN(N5187) );
  AOI22D1BWP30P140LVT U10497 ( .A1(i_data_bus[625]), .A2(n10470), .B1(
        i_data_bus[529]), .B2(n10471), .ZN(n7172) );
  AOI22D1BWP30P140LVT U10498 ( .A1(i_data_bus[561]), .A2(n10472), .B1(
        i_data_bus[593]), .B2(n10469), .ZN(n7171) );
  ND2D1BWP30P140LVT U10499 ( .A1(n7172), .A2(n7171), .ZN(N10822) );
  AOI22D1BWP30P140LVT U10500 ( .A1(i_data_bus[517]), .A2(n10566), .B1(
        i_data_bus[549]), .B2(n10567), .ZN(n7174) );
  AOI22D1BWP30P140LVT U10501 ( .A1(i_data_bus[613]), .A2(n10568), .B1(
        i_data_bus[581]), .B2(n10565), .ZN(n7173) );
  ND2D1BWP30P140LVT U10502 ( .A1(n7174), .A2(n7173), .ZN(N5188) );
  AOI22D1BWP30P140LVT U10503 ( .A1(i_data_bus[614]), .A2(n10470), .B1(
        i_data_bus[518]), .B2(n10471), .ZN(n7176) );
  AOI22D1BWP30P140LVT U10504 ( .A1(i_data_bus[550]), .A2(n10472), .B1(
        i_data_bus[582]), .B2(n10469), .ZN(n7175) );
  ND2D1BWP30P140LVT U10505 ( .A1(n7176), .A2(n7175), .ZN(N10811) );
  AOI22D1BWP30P140LVT U10506 ( .A1(i_data_bus[550]), .A2(n10567), .B1(
        i_data_bus[518]), .B2(n10566), .ZN(n7178) );
  AOI22D1BWP30P140LVT U10507 ( .A1(i_data_bus[614]), .A2(n10568), .B1(
        i_data_bus[582]), .B2(n10565), .ZN(n7177) );
  ND2D1BWP30P140LVT U10508 ( .A1(n7178), .A2(n7177), .ZN(N5189) );
  AOI22D1BWP30P140LVT U10509 ( .A1(i_data_bus[541]), .A2(n10471), .B1(
        i_data_bus[573]), .B2(n10472), .ZN(n7180) );
  AOI22D1BWP30P140LVT U10510 ( .A1(i_data_bus[637]), .A2(n10470), .B1(
        i_data_bus[605]), .B2(n10469), .ZN(n7179) );
  ND2D1BWP30P140LVT U10511 ( .A1(n7180), .A2(n7179), .ZN(N10834) );
  AOI22D1BWP30P140LVT U10512 ( .A1(i_data_bus[628]), .A2(n10568), .B1(
        i_data_bus[532]), .B2(n10566), .ZN(n7182) );
  AOI22D1BWP30P140LVT U10513 ( .A1(i_data_bus[564]), .A2(n10567), .B1(
        i_data_bus[596]), .B2(n10565), .ZN(n7181) );
  ND2D1BWP30P140LVT U10514 ( .A1(n7182), .A2(n7181), .ZN(N5203) );
  AOI22D1BWP30P140LVT U10515 ( .A1(i_data_bus[319]), .A2(n10606), .B1(
        i_data_bus[383]), .B2(n10608), .ZN(n7184) );
  AOI22D1BWP30P140LVT U10516 ( .A1(i_data_bus[351]), .A2(n10607), .B1(
        i_data_bus[287]), .B2(n10605), .ZN(n7183) );
  ND2D1BWP30P140LVT U10517 ( .A1(n7184), .A2(n7183), .ZN(N2908) );
  AOI22D1BWP30P140LVT U10518 ( .A1(i_data_bus[317]), .A2(n10606), .B1(
        i_data_bus[381]), .B2(n10608), .ZN(n7186) );
  AOI22D1BWP30P140LVT U10519 ( .A1(i_data_bus[349]), .A2(n10607), .B1(
        i_data_bus[285]), .B2(n10605), .ZN(n7185) );
  ND2D1BWP30P140LVT U10520 ( .A1(n7186), .A2(n7185), .ZN(N2906) );
  AOI22D1BWP30P140LVT U10521 ( .A1(i_data_bus[341]), .A2(n10607), .B1(
        i_data_bus[373]), .B2(n10608), .ZN(n7188) );
  AOI22D1BWP30P140LVT U10522 ( .A1(i_data_bus[309]), .A2(n10606), .B1(
        i_data_bus[277]), .B2(n10605), .ZN(n7187) );
  ND2D1BWP30P140LVT U10523 ( .A1(n7188), .A2(n7187), .ZN(N2898) );
  AOI22D1BWP30P140LVT U10524 ( .A1(i_data_bus[342]), .A2(n10607), .B1(
        i_data_bus[374]), .B2(n10608), .ZN(n7190) );
  AOI22D1BWP30P140LVT U10525 ( .A1(i_data_bus[310]), .A2(n10606), .B1(
        i_data_bus[278]), .B2(n10605), .ZN(n7189) );
  ND2D1BWP30P140LVT U10526 ( .A1(n7190), .A2(n7189), .ZN(N2899) );
  INR4D1BWP30P140LVT U10527 ( .A1(i_cmd[195]), .B1(i_cmd[211]), .B2(n9744), 
        .B3(n7192), .ZN(n10528) );
  NR4D1BWP30P140LVT U10528 ( .A1(i_cmd[219]), .A2(n7191), .A3(n9743), .A4(
        n7193), .ZN(n10525) );
  AOI22D1BWP30P140LVT U10529 ( .A1(i_data_bus[798]), .A2(n10528), .B1(
        i_data_bus[830]), .B2(n10525), .ZN(n7196) );
  INR4D1BWP30P140LVT U10530 ( .A1(i_cmd[211]), .B1(i_cmd[195]), .B2(n9741), 
        .B3(n7192), .ZN(n10527) );
  NR4D1BWP30P140LVT U10531 ( .A1(i_cmd[203]), .A2(n9747), .A3(n7194), .A4(
        n7193), .ZN(n10526) );
  AOI22D1BWP30P140LVT U10532 ( .A1(i_data_bus[862]), .A2(n10527), .B1(
        i_data_bus[894]), .B2(n10526), .ZN(n7195) );
  ND2D1BWP30P140LVT U10533 ( .A1(n7196), .A2(n7195), .ZN(N7519) );
  NR4D1BWP30P140LVT U10534 ( .A1(i_cmd[177]), .A2(n7199), .A3(n9843), .A4(
        n7197), .ZN(n10596) );
  INR4D1BWP30P140LVT U10535 ( .A1(i_cmd[185]), .B1(i_cmd[169]), .B2(n9844), 
        .B3(n7200), .ZN(n10595) );
  AOI22D1BWP30P140LVT U10536 ( .A1(i_data_bus[643]), .A2(n10596), .B1(
        i_data_bus[739]), .B2(n10595), .ZN(n7202) );
  NR4D1BWP30P140LVT U10537 ( .A1(i_cmd[161]), .A2(n7199), .A3(n9850), .A4(
        n7198), .ZN(n10594) );
  INR4D1BWP30P140LVT U10538 ( .A1(i_cmd[169]), .B1(i_cmd[185]), .B2(n9847), 
        .B3(n7200), .ZN(n10593) );
  AOI22D1BWP30P140LVT U10539 ( .A1(i_data_bus[707]), .A2(n10594), .B1(
        i_data_bus[675]), .B2(n10593), .ZN(n7201) );
  ND2D1BWP30P140LVT U10540 ( .A1(n7202), .A2(n7201), .ZN(N3528) );
  AOI22D1BWP30P140LVT U10541 ( .A1(i_data_bus[755]), .A2(n10595), .B1(
        i_data_bus[723]), .B2(n10594), .ZN(n7204) );
  AOI22D1BWP30P140LVT U10542 ( .A1(i_data_bus[659]), .A2(n10596), .B1(
        i_data_bus[691]), .B2(n10593), .ZN(n7203) );
  ND2D1BWP30P140LVT U10543 ( .A1(n7204), .A2(n7203), .ZN(N3544) );
  AOI22D1BWP30P140LVT U10544 ( .A1(i_data_bus[722]), .A2(n10594), .B1(
        i_data_bus[658]), .B2(n10596), .ZN(n7206) );
  AOI22D1BWP30P140LVT U10545 ( .A1(i_data_bus[754]), .A2(n10595), .B1(
        i_data_bus[690]), .B2(n10593), .ZN(n7205) );
  ND2D1BWP30P140LVT U10546 ( .A1(n7206), .A2(n7205), .ZN(N3543) );
  AOI22D1BWP30P140LVT U10547 ( .A1(i_data_bus[667]), .A2(n10596), .B1(
        i_data_bus[731]), .B2(n10594), .ZN(n7208) );
  AOI22D1BWP30P140LVT U10548 ( .A1(i_data_bus[763]), .A2(n10595), .B1(
        i_data_bus[699]), .B2(n10593), .ZN(n7207) );
  ND2D1BWP30P140LVT U10549 ( .A1(n7208), .A2(n7207), .ZN(N3552) );
  AOI22D1BWP30P140LVT U10550 ( .A1(i_data_bus[924]), .A2(n10395), .B1(
        i_data_bus[956]), .B2(n10394), .ZN(n7210) );
  AOI22D1BWP30P140LVT U10551 ( .A1(i_data_bus[988]), .A2(n10396), .B1(
        i_data_bus[1020]), .B2(n10393), .ZN(n7209) );
  ND2D1BWP30P140LVT U10552 ( .A1(n7210), .A2(n7209), .ZN(N15229) );
  AOI22D1BWP30P140LVT U10553 ( .A1(i_data_bus[961]), .A2(n10396), .B1(
        i_data_bus[897]), .B2(n10395), .ZN(n7212) );
  AOI22D1BWP30P140LVT U10554 ( .A1(i_data_bus[929]), .A2(n10394), .B1(
        i_data_bus[993]), .B2(n10393), .ZN(n7211) );
  ND2D1BWP30P140LVT U10555 ( .A1(n7212), .A2(n7211), .ZN(N15202) );
  AOI22D1BWP30P140LVT U10556 ( .A1(i_data_bus[970]), .A2(n10396), .B1(
        i_data_bus[938]), .B2(n10394), .ZN(n7214) );
  AOI22D1BWP30P140LVT U10557 ( .A1(i_data_bus[906]), .A2(n10395), .B1(
        i_data_bus[1002]), .B2(n10393), .ZN(n7213) );
  ND2D1BWP30P140LVT U10558 ( .A1(n7214), .A2(n7213), .ZN(N15211) );
  AOI22D1BWP30P140LVT U10559 ( .A1(i_data_bus[715]), .A2(n10594), .B1(
        i_data_bus[651]), .B2(n10596), .ZN(n7216) );
  AOI22D1BWP30P140LVT U10560 ( .A1(i_data_bus[747]), .A2(n10595), .B1(
        i_data_bus[683]), .B2(n10593), .ZN(n7215) );
  ND2D1BWP30P140LVT U10561 ( .A1(n7216), .A2(n7215), .ZN(N3536) );
  AOI22D1BWP30P140LVT U10562 ( .A1(i_data_bus[257]), .A2(n10605), .B1(
        i_data_bus[353]), .B2(n10608), .ZN(n7218) );
  AOI22D1BWP30P140LVT U10563 ( .A1(i_data_bus[321]), .A2(n10607), .B1(
        i_data_bus[289]), .B2(n10606), .ZN(n7217) );
  ND2D1BWP30P140LVT U10564 ( .A1(n7218), .A2(n7217), .ZN(N2878) );
  AOI22D1BWP30P140LVT U10565 ( .A1(i_data_bus[266]), .A2(n10605), .B1(
        i_data_bus[362]), .B2(n10608), .ZN(n7220) );
  AOI22D1BWP30P140LVT U10566 ( .A1(i_data_bus[330]), .A2(n10607), .B1(
        i_data_bus[298]), .B2(n10606), .ZN(n7219) );
  ND2D1BWP30P140LVT U10567 ( .A1(n7220), .A2(n7219), .ZN(N2887) );
  AOI22D1BWP30P140LVT U10568 ( .A1(i_data_bus[141]), .A2(n10481), .B1(
        i_data_bus[237]), .B2(n10484), .ZN(n7222) );
  AOI22D1BWP30P140LVT U10569 ( .A1(i_data_bus[205]), .A2(n10482), .B1(
        i_data_bus[173]), .B2(n10483), .ZN(n7221) );
  ND2D1BWP30P140LVT U10570 ( .A1(n7222), .A2(n7221), .ZN(N10170) );
  AOI22D1BWP30P140LVT U10571 ( .A1(i_data_bus[203]), .A2(n10482), .B1(
        i_data_bus[235]), .B2(n10484), .ZN(n7224) );
  AOI22D1BWP30P140LVT U10572 ( .A1(i_data_bus[139]), .A2(n10481), .B1(
        i_data_bus[171]), .B2(n10483), .ZN(n7223) );
  ND2D1BWP30P140LVT U10573 ( .A1(n7224), .A2(n7223), .ZN(N10168) );
  AOI22D1BWP30P140LVT U10574 ( .A1(i_data_bus[895]), .A2(n10398), .B1(
        i_data_bus[831]), .B2(n10400), .ZN(n7226) );
  AOI22D1BWP30P140LVT U10575 ( .A1(i_data_bus[863]), .A2(n10399), .B1(
        i_data_bus[799]), .B2(n10397), .ZN(n7225) );
  ND2D1BWP30P140LVT U10576 ( .A1(n7226), .A2(n7225), .ZN(N15016) );
  AOI22D1BWP30P140LVT U10577 ( .A1(i_data_bus[870]), .A2(n10398), .B1(
        i_data_bus[806]), .B2(n10400), .ZN(n7228) );
  AOI22D1BWP30P140LVT U10578 ( .A1(i_data_bus[838]), .A2(n10399), .B1(
        i_data_bus[774]), .B2(n10397), .ZN(n7227) );
  ND2D1BWP30P140LVT U10579 ( .A1(n7228), .A2(n7227), .ZN(N14991) );
  AOI22D1BWP30P140LVT U10580 ( .A1(i_data_bus[856]), .A2(n10399), .B1(
        i_data_bus[824]), .B2(n10400), .ZN(n7230) );
  AOI22D1BWP30P140LVT U10581 ( .A1(i_data_bus[888]), .A2(n10398), .B1(
        i_data_bus[792]), .B2(n10397), .ZN(n7229) );
  ND2D1BWP30P140LVT U10582 ( .A1(n7230), .A2(n7229), .ZN(N15009) );
  AOI22D1BWP30P140LVT U10583 ( .A1(i_data_bus[850]), .A2(n10399), .B1(
        i_data_bus[818]), .B2(n10400), .ZN(n7232) );
  AOI22D1BWP30P140LVT U10584 ( .A1(i_data_bus[882]), .A2(n10398), .B1(
        i_data_bus[786]), .B2(n10397), .ZN(n7231) );
  ND2D1BWP30P140LVT U10585 ( .A1(n7232), .A2(n7231), .ZN(N15003) );
  AOI22D1BWP30P140LVT U10586 ( .A1(i_data_bus[890]), .A2(n10398), .B1(
        i_data_bus[826]), .B2(n10400), .ZN(n7234) );
  AOI22D1BWP30P140LVT U10587 ( .A1(i_data_bus[858]), .A2(n10399), .B1(
        i_data_bus[794]), .B2(n10397), .ZN(n7233) );
  ND2D1BWP30P140LVT U10588 ( .A1(n7234), .A2(n7233), .ZN(N15011) );
  AOI22D1BWP30P140LVT U10589 ( .A1(i_data_bus[847]), .A2(n10399), .B1(
        i_data_bus[815]), .B2(n10400), .ZN(n7236) );
  AOI22D1BWP30P140LVT U10590 ( .A1(i_data_bus[783]), .A2(n10397), .B1(
        i_data_bus[879]), .B2(n10398), .ZN(n7235) );
  ND2D1BWP30P140LVT U10591 ( .A1(n7236), .A2(n7235), .ZN(N15000) );
  AOI22D1BWP30P140LVT U10592 ( .A1(i_data_bus[776]), .A2(n10397), .B1(
        i_data_bus[808]), .B2(n10400), .ZN(n7238) );
  AOI22D1BWP30P140LVT U10593 ( .A1(i_data_bus[840]), .A2(n10399), .B1(
        i_data_bus[872]), .B2(n10398), .ZN(n7237) );
  ND2D1BWP30P140LVT U10594 ( .A1(n7238), .A2(n7237), .ZN(N14993) );
  AOI22D1BWP30P140LVT U10595 ( .A1(i_data_bus[778]), .A2(n10397), .B1(
        i_data_bus[810]), .B2(n10400), .ZN(n7240) );
  AOI22D1BWP30P140LVT U10596 ( .A1(i_data_bus[842]), .A2(n10399), .B1(
        i_data_bus[874]), .B2(n10398), .ZN(n7239) );
  ND2D1BWP30P140LVT U10597 ( .A1(n7240), .A2(n7239), .ZN(N14995) );
  AOI22D1BWP30P140LVT U10598 ( .A1(i_data_bus[772]), .A2(n10397), .B1(
        i_data_bus[804]), .B2(n10400), .ZN(n7242) );
  AOI22D1BWP30P140LVT U10599 ( .A1(i_data_bus[836]), .A2(n10399), .B1(
        i_data_bus[868]), .B2(n10398), .ZN(n7241) );
  ND2D1BWP30P140LVT U10600 ( .A1(n7242), .A2(n7241), .ZN(N14989) );
  AOI22D1BWP30P140LVT U10601 ( .A1(i_data_bus[848]), .A2(n10399), .B1(
        i_data_bus[816]), .B2(n10400), .ZN(n7244) );
  AOI22D1BWP30P140LVT U10602 ( .A1(i_data_bus[784]), .A2(n10397), .B1(
        i_data_bus[880]), .B2(n10398), .ZN(n7243) );
  ND2D1BWP30P140LVT U10603 ( .A1(n7244), .A2(n7243), .ZN(N15001) );
  AOI22D1BWP30P140LVT U10604 ( .A1(i_data_bus[60]), .A2(n10583), .B1(
        i_data_bus[28]), .B2(n10581), .ZN(n7246) );
  AOI22D1BWP30P140LVT U10605 ( .A1(i_data_bus[124]), .A2(n10584), .B1(
        i_data_bus[92]), .B2(n10582), .ZN(n7245) );
  ND2D1BWP30P140LVT U10606 ( .A1(n7246), .A2(n7245), .ZN(N4347) );
  AOI22D1BWP30P140LVT U10607 ( .A1(i_data_bus[322]), .A2(n10509), .B1(
        i_data_bus[354]), .B2(n10511), .ZN(n7248) );
  AOI22D1BWP30P140LVT U10608 ( .A1(i_data_bus[258]), .A2(n10510), .B1(
        i_data_bus[290]), .B2(n10512), .ZN(n7247) );
  ND2D1BWP30P140LVT U10609 ( .A1(n7248), .A2(n7247), .ZN(N8501) );
  AOI22D1BWP30P140LVT U10610 ( .A1(i_data_bus[317]), .A2(n10512), .B1(
        i_data_bus[381]), .B2(n10511), .ZN(n7250) );
  AOI22D1BWP30P140LVT U10611 ( .A1(i_data_bus[349]), .A2(n10509), .B1(
        i_data_bus[285]), .B2(n10510), .ZN(n7249) );
  ND2D1BWP30P140LVT U10612 ( .A1(n7250), .A2(n7249), .ZN(N8528) );
  AOI22D1BWP30P140LVT U10613 ( .A1(i_data_bus[341]), .A2(n10509), .B1(
        i_data_bus[373]), .B2(n10511), .ZN(n7252) );
  AOI22D1BWP30P140LVT U10614 ( .A1(i_data_bus[309]), .A2(n10512), .B1(
        i_data_bus[277]), .B2(n10510), .ZN(n7251) );
  ND2D1BWP30P140LVT U10615 ( .A1(n7252), .A2(n7251), .ZN(N8520) );
  NR4D1BWP30P140LVT U10616 ( .A1(i_cmd[140]), .A2(n7255), .A3(n9837), .A4(
        n7253), .ZN(n10501) );
  INR4D1BWP30P140LVT U10617 ( .A1(i_cmd[132]), .B1(i_cmd[148]), .B2(n9839), 
        .B3(n7256), .ZN(n10503) );
  AOI22D1BWP30P140LVT U10618 ( .A1(i_data_bus[621]), .A2(n10501), .B1(
        i_data_bus[525]), .B2(n10503), .ZN(n7258) );
  NR4D1BWP30P140LVT U10619 ( .A1(i_cmd[156]), .A2(n7255), .A3(n9833), .A4(
        n7254), .ZN(n10504) );
  INR4D1BWP30P140LVT U10620 ( .A1(i_cmd[148]), .B1(i_cmd[132]), .B2(n9834), 
        .B3(n7256), .ZN(n10502) );
  AOI22D1BWP30P140LVT U10621 ( .A1(i_data_bus[557]), .A2(n10504), .B1(
        i_data_bus[589]), .B2(n10502), .ZN(n7257) );
  ND2D1BWP30P140LVT U10622 ( .A1(n7258), .A2(n7257), .ZN(N8944) );
  AOI22D1BWP30P140LVT U10623 ( .A1(i_data_bus[521]), .A2(n10503), .B1(
        i_data_bus[553]), .B2(n10504), .ZN(n7260) );
  AOI22D1BWP30P140LVT U10624 ( .A1(i_data_bus[617]), .A2(n10501), .B1(
        i_data_bus[585]), .B2(n10502), .ZN(n7259) );
  ND2D1BWP30P140LVT U10625 ( .A1(n7260), .A2(n7259), .ZN(N8940) );
  AOI22D1BWP30P140LVT U10626 ( .A1(i_data_bus[560]), .A2(n10504), .B1(
        i_data_bus[528]), .B2(n10503), .ZN(n7262) );
  AOI22D1BWP30P140LVT U10627 ( .A1(i_data_bus[624]), .A2(n10501), .B1(
        i_data_bus[592]), .B2(n10502), .ZN(n7261) );
  ND2D1BWP30P140LVT U10628 ( .A1(n7262), .A2(n7261), .ZN(N8947) );
  AOI22D1BWP30P140LVT U10629 ( .A1(i_data_bus[635]), .A2(n10501), .B1(
        i_data_bus[539]), .B2(n10503), .ZN(n7264) );
  AOI22D1BWP30P140LVT U10630 ( .A1(i_data_bus[571]), .A2(n10504), .B1(
        i_data_bus[603]), .B2(n10502), .ZN(n7263) );
  ND2D1BWP30P140LVT U10631 ( .A1(n7264), .A2(n7263), .ZN(N8958) );
  AOI22D1BWP30P140LVT U10632 ( .A1(i_data_bus[542]), .A2(n10503), .B1(
        i_data_bus[574]), .B2(n10504), .ZN(n7266) );
  AOI22D1BWP30P140LVT U10633 ( .A1(i_data_bus[638]), .A2(n10501), .B1(
        i_data_bus[606]), .B2(n10502), .ZN(n7265) );
  ND2D1BWP30P140LVT U10634 ( .A1(n7266), .A2(n7265), .ZN(N8961) );
  AOI22D1BWP30P140LVT U10635 ( .A1(i_data_bus[536]), .A2(n10405), .B1(
        i_data_bus[632]), .B2(n10407), .ZN(n7268) );
  AOI22D1BWP30P140LVT U10636 ( .A1(i_data_bus[600]), .A2(n10408), .B1(
        i_data_bus[568]), .B2(n10406), .ZN(n7267) );
  ND2D1BWP30P140LVT U10637 ( .A1(n7268), .A2(n7267), .ZN(N14577) );
  INR4D1BWP30P140LVT U10638 ( .A1(i_cmd[13]), .B1(i_cmd[29]), .B2(n10018), 
        .B3(n7269), .ZN(n10485) );
  INR4D1BWP30P140LVT U10639 ( .A1(i_cmd[29]), .B1(i_cmd[13]), .B2(n10019), 
        .B3(n7269), .ZN(n10488) );
  AOI22D1BWP30P140LVT U10640 ( .A1(i_data_bus[35]), .A2(n10485), .B1(
        i_data_bus[99]), .B2(n10488), .ZN(n7274) );
  NR4D1BWP30P140LVT U10641 ( .A1(i_cmd[5]), .A2(n7270), .A3(n10014), .A4(n7271), .ZN(n10487) );
  NR4D1BWP30P140LVT U10642 ( .A1(i_cmd[21]), .A2(n10013), .A3(n7272), .A4(
        n7271), .ZN(n10486) );
  AOI22D1BWP30P140LVT U10643 ( .A1(i_data_bus[67]), .A2(n10487), .B1(
        i_data_bus[3]), .B2(n10486), .ZN(n7273) );
  ND2D1BWP30P140LVT U10644 ( .A1(n7274), .A2(n7273), .ZN(N9944) );
  AOI22D1BWP30P140LVT U10645 ( .A1(i_data_bus[48]), .A2(n10485), .B1(
        i_data_bus[112]), .B2(n10488), .ZN(n7276) );
  AOI22D1BWP30P140LVT U10646 ( .A1(i_data_bus[80]), .A2(n10487), .B1(
        i_data_bus[16]), .B2(n10486), .ZN(n7275) );
  ND2D1BWP30P140LVT U10647 ( .A1(n7276), .A2(n7275), .ZN(N9957) );
  AOI22D1BWP30P140LVT U10648 ( .A1(i_data_bus[105]), .A2(n10488), .B1(
        i_data_bus[41]), .B2(n10485), .ZN(n7278) );
  AOI22D1BWP30P140LVT U10649 ( .A1(i_data_bus[73]), .A2(n10487), .B1(
        i_data_bus[9]), .B2(n10486), .ZN(n7277) );
  ND2D1BWP30P140LVT U10650 ( .A1(n7278), .A2(n7277), .ZN(N9950) );
  AOI22D1BWP30P140LVT U10651 ( .A1(i_data_bus[33]), .A2(n10485), .B1(
        i_data_bus[97]), .B2(n10488), .ZN(n7280) );
  AOI22D1BWP30P140LVT U10652 ( .A1(i_data_bus[65]), .A2(n10487), .B1(
        i_data_bus[1]), .B2(n10486), .ZN(n7279) );
  ND2D1BWP30P140LVT U10653 ( .A1(n7280), .A2(n7279), .ZN(N9942) );
  AOI22D1BWP30P140LVT U10654 ( .A1(i_data_bus[127]), .A2(n10488), .B1(
        i_data_bus[63]), .B2(n10485), .ZN(n7282) );
  AOI22D1BWP30P140LVT U10655 ( .A1(i_data_bus[95]), .A2(n10487), .B1(
        i_data_bus[31]), .B2(n10486), .ZN(n7281) );
  ND2D1BWP30P140LVT U10656 ( .A1(n7282), .A2(n7281), .ZN(N9972) );
  AOI22D1BWP30P140LVT U10657 ( .A1(i_data_bus[75]), .A2(n10487), .B1(
        i_data_bus[107]), .B2(n10488), .ZN(n7284) );
  AOI22D1BWP30P140LVT U10658 ( .A1(i_data_bus[43]), .A2(n10485), .B1(
        i_data_bus[11]), .B2(n10486), .ZN(n7283) );
  ND2D1BWP30P140LVT U10659 ( .A1(n7284), .A2(n7283), .ZN(N9952) );
  AOI22D1BWP30P140LVT U10660 ( .A1(i_data_bus[114]), .A2(n10488), .B1(
        i_data_bus[50]), .B2(n10485), .ZN(n7286) );
  AOI22D1BWP30P140LVT U10661 ( .A1(i_data_bus[82]), .A2(n10487), .B1(
        i_data_bus[18]), .B2(n10486), .ZN(n7285) );
  ND2D1BWP30P140LVT U10662 ( .A1(n7286), .A2(n7285), .ZN(N9959) );
  AOI22D1BWP30P140LVT U10663 ( .A1(i_data_bus[122]), .A2(n10488), .B1(
        i_data_bus[58]), .B2(n10485), .ZN(n7288) );
  AOI22D1BWP30P140LVT U10664 ( .A1(i_data_bus[90]), .A2(n10487), .B1(
        i_data_bus[26]), .B2(n10486), .ZN(n7287) );
  ND2D1BWP30P140LVT U10665 ( .A1(n7288), .A2(n7287), .ZN(N9967) );
  INR4D1BWP30P140LVT U10666 ( .A1(i_cmd[180]), .B1(i_cmd[164]), .B2(n9850), 
        .B3(n7292), .ZN(n10497) );
  NR4D1BWP30P140LVT U10667 ( .A1(i_cmd[172]), .A2(n7291), .A3(n9844), .A4(
        n7289), .ZN(n10500) );
  AOI22D1BWP30P140LVT U10668 ( .A1(i_data_bus[734]), .A2(n10497), .B1(
        i_data_bus[766]), .B2(n10500), .ZN(n7294) );
  NR4D1BWP30P140LVT U10669 ( .A1(i_cmd[188]), .A2(n7291), .A3(n9847), .A4(
        n7290), .ZN(n10499) );
  INR4D1BWP30P140LVT U10670 ( .A1(i_cmd[164]), .B1(i_cmd[180]), .B2(n9843), 
        .B3(n7292), .ZN(n10498) );
  AOI22D1BWP30P140LVT U10671 ( .A1(i_data_bus[702]), .A2(n10499), .B1(
        i_data_bus[670]), .B2(n10498), .ZN(n7293) );
  ND2D1BWP30P140LVT U10672 ( .A1(n7294), .A2(n7293), .ZN(N9177) );
  AOI22D1BWP30P140LVT U10673 ( .A1(i_data_bus[719]), .A2(n10497), .B1(
        i_data_bus[751]), .B2(n10500), .ZN(n7296) );
  AOI22D1BWP30P140LVT U10674 ( .A1(i_data_bus[687]), .A2(n10499), .B1(
        i_data_bus[655]), .B2(n10498), .ZN(n7295) );
  ND2D1BWP30P140LVT U10675 ( .A1(n7296), .A2(n7295), .ZN(N9162) );
  AOI22D1BWP30P140LVT U10676 ( .A1(i_data_bus[735]), .A2(n10497), .B1(
        i_data_bus[767]), .B2(n10500), .ZN(n7298) );
  AOI22D1BWP30P140LVT U10677 ( .A1(i_data_bus[703]), .A2(n10499), .B1(
        i_data_bus[671]), .B2(n10498), .ZN(n7297) );
  ND2D1BWP30P140LVT U10678 ( .A1(n7298), .A2(n7297), .ZN(N9178) );
  AOI22D1BWP30P140LVT U10679 ( .A1(i_data_bus[561]), .A2(n10406), .B1(
        i_data_bus[625]), .B2(n10407), .ZN(n7300) );
  AOI22D1BWP30P140LVT U10680 ( .A1(i_data_bus[593]), .A2(n10408), .B1(
        i_data_bus[529]), .B2(n10405), .ZN(n7299) );
  ND2D1BWP30P140LVT U10681 ( .A1(n7300), .A2(n7299), .ZN(N14570) );
  AOI22D1BWP30P140LVT U10682 ( .A1(i_data_bus[559]), .A2(n10406), .B1(
        i_data_bus[623]), .B2(n10407), .ZN(n7302) );
  AOI22D1BWP30P140LVT U10683 ( .A1(i_data_bus[591]), .A2(n10408), .B1(
        i_data_bus[527]), .B2(n10405), .ZN(n7301) );
  ND2D1BWP30P140LVT U10684 ( .A1(n7302), .A2(n7301), .ZN(N14568) );
  AOI22D1BWP30P140LVT U10685 ( .A1(i_data_bus[566]), .A2(n10406), .B1(
        i_data_bus[630]), .B2(n10407), .ZN(n7304) );
  AOI22D1BWP30P140LVT U10686 ( .A1(i_data_bus[598]), .A2(n10408), .B1(
        i_data_bus[534]), .B2(n10405), .ZN(n7303) );
  ND2D1BWP30P140LVT U10687 ( .A1(n7304), .A2(n7303), .ZN(N14575) );
  AOI22D1BWP30P140LVT U10688 ( .A1(i_data_bus[526]), .A2(n10405), .B1(
        i_data_bus[622]), .B2(n10407), .ZN(n7306) );
  AOI22D1BWP30P140LVT U10689 ( .A1(i_data_bus[558]), .A2(n10406), .B1(
        i_data_bus[590]), .B2(n10408), .ZN(n7305) );
  ND2D1BWP30P140LVT U10690 ( .A1(n7306), .A2(n7305), .ZN(N14567) );
  AOI22D1BWP30P140LVT U10691 ( .A1(i_data_bus[571]), .A2(n10406), .B1(
        i_data_bus[635]), .B2(n10407), .ZN(n7308) );
  AOI22D1BWP30P140LVT U10692 ( .A1(i_data_bus[539]), .A2(n10405), .B1(
        i_data_bus[603]), .B2(n10408), .ZN(n7307) );
  ND2D1BWP30P140LVT U10693 ( .A1(n7308), .A2(n7307), .ZN(N14580) );
  AOI22D1BWP30P140LVT U10694 ( .A1(i_data_bus[556]), .A2(n10406), .B1(
        i_data_bus[620]), .B2(n10407), .ZN(n7310) );
  AOI22D1BWP30P140LVT U10695 ( .A1(i_data_bus[524]), .A2(n10405), .B1(
        i_data_bus[588]), .B2(n10408), .ZN(n7309) );
  ND2D1BWP30P140LVT U10696 ( .A1(n7310), .A2(n7309), .ZN(N14565) );
  INR4D1BWP30P140LVT U10697 ( .A1(i_cmd[11]), .B1(i_cmd[27]), .B2(n10018), 
        .B3(n7314), .ZN(n10550) );
  NR4D1BWP30P140LVT U10698 ( .A1(i_cmd[3]), .A2(n7313), .A3(n10014), .A4(n7311), .ZN(n10551) );
  AOI22D1BWP30P140LVT U10699 ( .A1(i_data_bus[61]), .A2(n10550), .B1(
        i_data_bus[93]), .B2(n10551), .ZN(n7316) );
  NR4D1BWP30P140LVT U10700 ( .A1(i_cmd[19]), .A2(n7313), .A3(n10013), .A4(
        n7312), .ZN(n10552) );
  INR4D1BWP30P140LVT U10701 ( .A1(i_cmd[27]), .B1(i_cmd[11]), .B2(n10019), 
        .B3(n7314), .ZN(n10549) );
  AOI22D1BWP30P140LVT U10702 ( .A1(i_data_bus[29]), .A2(n10552), .B1(
        i_data_bus[125]), .B2(n10549), .ZN(n7315) );
  ND2D1BWP30P140LVT U10703 ( .A1(n7316), .A2(n7315), .ZN(N6222) );
  AOI22D1BWP30P140LVT U10704 ( .A1(i_data_bus[47]), .A2(n10550), .B1(
        i_data_bus[79]), .B2(n10551), .ZN(n7318) );
  AOI22D1BWP30P140LVT U10705 ( .A1(i_data_bus[15]), .A2(n10552), .B1(
        i_data_bus[111]), .B2(n10549), .ZN(n7317) );
  ND2D1BWP30P140LVT U10706 ( .A1(n7318), .A2(n7317), .ZN(N6208) );
  AOI22D1BWP30P140LVT U10707 ( .A1(i_data_bus[989]), .A2(n10490), .B1(
        i_data_bus[957]), .B2(n10491), .ZN(n7320) );
  AOI22D1BWP30P140LVT U10708 ( .A1(i_data_bus[925]), .A2(n10492), .B1(
        i_data_bus[1021]), .B2(n10489), .ZN(n7319) );
  ND2D1BWP30P140LVT U10709 ( .A1(n7320), .A2(n7319), .ZN(N9608) );
  AOI22D1BWP30P140LVT U10710 ( .A1(i_data_bus[966]), .A2(n10490), .B1(
        i_data_bus[902]), .B2(n10492), .ZN(n7322) );
  AOI22D1BWP30P140LVT U10711 ( .A1(i_data_bus[934]), .A2(n10491), .B1(
        i_data_bus[998]), .B2(n10489), .ZN(n7321) );
  ND2D1BWP30P140LVT U10712 ( .A1(n7322), .A2(n7321), .ZN(N9585) );
  AOI22D1BWP30P140LVT U10713 ( .A1(i_data_bus[921]), .A2(n10492), .B1(
        i_data_bus[953]), .B2(n10491), .ZN(n7324) );
  AOI22D1BWP30P140LVT U10714 ( .A1(i_data_bus[985]), .A2(n10490), .B1(
        i_data_bus[1017]), .B2(n10489), .ZN(n7323) );
  ND2D1BWP30P140LVT U10715 ( .A1(n7324), .A2(n7323), .ZN(N9604) );
  AOI22D1BWP30P140LVT U10716 ( .A1(i_data_bus[974]), .A2(n10490), .B1(
        i_data_bus[942]), .B2(n10491), .ZN(n7326) );
  AOI22D1BWP30P140LVT U10717 ( .A1(i_data_bus[910]), .A2(n10492), .B1(
        i_data_bus[1006]), .B2(n10489), .ZN(n7325) );
  ND2D1BWP30P140LVT U10718 ( .A1(n7326), .A2(n7325), .ZN(N9593) );
  AOI22D1BWP30P140LVT U10719 ( .A1(i_data_bus[968]), .A2(n10490), .B1(
        i_data_bus[904]), .B2(n10492), .ZN(n7328) );
  AOI22D1BWP30P140LVT U10720 ( .A1(i_data_bus[936]), .A2(n10491), .B1(
        i_data_bus[1000]), .B2(n10489), .ZN(n7327) );
  ND2D1BWP30P140LVT U10721 ( .A1(n7328), .A2(n7327), .ZN(N9587) );
  AOI22D1BWP30P140LVT U10722 ( .A1(i_data_bus[777]), .A2(n10462), .B1(
        i_data_bus[873]), .B2(n10461), .ZN(n7330) );
  AOI22D1BWP30P140LVT U10723 ( .A1(i_data_bus[841]), .A2(n10463), .B1(
        i_data_bus[809]), .B2(n10464), .ZN(n7329) );
  ND2D1BWP30P140LVT U10724 ( .A1(n7330), .A2(n7329), .ZN(N11246) );
  AOI22D1BWP30P140LVT U10725 ( .A1(i_data_bus[887]), .A2(n10461), .B1(
        i_data_bus[791]), .B2(n10462), .ZN(n7332) );
  AOI22D1BWP30P140LVT U10726 ( .A1(i_data_bus[855]), .A2(n10463), .B1(
        i_data_bus[823]), .B2(n10464), .ZN(n7331) );
  ND2D1BWP30P140LVT U10727 ( .A1(n7332), .A2(n7331), .ZN(N11260) );
  AOI22D1BWP30P140LVT U10728 ( .A1(i_data_bus[768]), .A2(n10462), .B1(
        i_data_bus[864]), .B2(n10461), .ZN(n7334) );
  AOI22D1BWP30P140LVT U10729 ( .A1(i_data_bus[832]), .A2(n10463), .B1(
        i_data_bus[800]), .B2(n10464), .ZN(n7333) );
  ND2D1BWP30P140LVT U10730 ( .A1(n7334), .A2(n7333), .ZN(N11237) );
  AOI22D1BWP30P140LVT U10731 ( .A1(i_data_bus[836]), .A2(n10463), .B1(
        i_data_bus[772]), .B2(n10462), .ZN(n7336) );
  AOI22D1BWP30P140LVT U10732 ( .A1(i_data_bus[868]), .A2(n10461), .B1(
        i_data_bus[804]), .B2(n10464), .ZN(n7335) );
  ND2D1BWP30P140LVT U10733 ( .A1(n7336), .A2(n7335), .ZN(N11241) );
  AOI22D1BWP30P140LVT U10734 ( .A1(i_data_bus[834]), .A2(n10463), .B1(
        i_data_bus[770]), .B2(n10462), .ZN(n7338) );
  AOI22D1BWP30P140LVT U10735 ( .A1(i_data_bus[866]), .A2(n10461), .B1(
        i_data_bus[802]), .B2(n10464), .ZN(n7337) );
  ND2D1BWP30P140LVT U10736 ( .A1(n7338), .A2(n7337), .ZN(N11239) );
  AOI22D1BWP30P140LVT U10737 ( .A1(i_data_bus[840]), .A2(n10463), .B1(
        i_data_bus[872]), .B2(n10461), .ZN(n7340) );
  AOI22D1BWP30P140LVT U10738 ( .A1(i_data_bus[776]), .A2(n10462), .B1(
        i_data_bus[808]), .B2(n10464), .ZN(n7339) );
  ND2D1BWP30P140LVT U10739 ( .A1(n7340), .A2(n7339), .ZN(N11245) );
  AOI22D1BWP30P140LVT U10740 ( .A1(i_data_bus[848]), .A2(n10463), .B1(
        i_data_bus[880]), .B2(n10461), .ZN(n7342) );
  AOI22D1BWP30P140LVT U10741 ( .A1(i_data_bus[784]), .A2(n10462), .B1(
        i_data_bus[816]), .B2(n10464), .ZN(n7341) );
  ND2D1BWP30P140LVT U10742 ( .A1(n7342), .A2(n7341), .ZN(N11253) );
  AOI22D1BWP30P140LVT U10743 ( .A1(i_data_bus[858]), .A2(n10463), .B1(
        i_data_bus[890]), .B2(n10461), .ZN(n7344) );
  AOI22D1BWP30P140LVT U10744 ( .A1(i_data_bus[794]), .A2(n10462), .B1(
        i_data_bus[826]), .B2(n10464), .ZN(n7343) );
  ND2D1BWP30P140LVT U10745 ( .A1(n7344), .A2(n7343), .ZN(N11263) );
  AOI22D1BWP30P140LVT U10746 ( .A1(i_data_bus[444]), .A2(n10474), .B1(
        i_data_bus[508]), .B2(n10475), .ZN(n7346) );
  AOI22D1BWP30P140LVT U10747 ( .A1(i_data_bus[476]), .A2(n10476), .B1(
        i_data_bus[412]), .B2(n10473), .ZN(n7345) );
  ND2D1BWP30P140LVT U10748 ( .A1(n7346), .A2(n7345), .ZN(N10617) );
  AOI22D1BWP30P140LVT U10749 ( .A1(i_data_bus[249]), .A2(n10580), .B1(
        i_data_bus[153]), .B2(n10577), .ZN(n7348) );
  AOI22D1BWP30P140LVT U10750 ( .A1(i_data_bus[185]), .A2(n10579), .B1(
        i_data_bus[217]), .B2(n10578), .ZN(n7347) );
  ND2D1BWP30P140LVT U10751 ( .A1(n7348), .A2(n7347), .ZN(N4560) );
  AOI22D1BWP30P140LVT U10752 ( .A1(i_data_bus[431]), .A2(n10474), .B1(
        i_data_bus[463]), .B2(n10476), .ZN(n7350) );
  AOI22D1BWP30P140LVT U10753 ( .A1(i_data_bus[495]), .A2(n10475), .B1(
        i_data_bus[399]), .B2(n10473), .ZN(n7349) );
  ND2D1BWP30P140LVT U10754 ( .A1(n7350), .A2(n7349), .ZN(N10604) );
  AOI22D1BWP30P140LVT U10755 ( .A1(i_data_bus[491]), .A2(n10475), .B1(
        i_data_bus[459]), .B2(n10476), .ZN(n7352) );
  AOI22D1BWP30P140LVT U10756 ( .A1(i_data_bus[427]), .A2(n10474), .B1(
        i_data_bus[395]), .B2(n10473), .ZN(n7351) );
  ND2D1BWP30P140LVT U10757 ( .A1(n7352), .A2(n7351), .ZN(N10600) );
  AOI22D1BWP30P140LVT U10758 ( .A1(i_data_bus[471]), .A2(n10476), .B1(
        i_data_bus[439]), .B2(n10474), .ZN(n7354) );
  AOI22D1BWP30P140LVT U10759 ( .A1(i_data_bus[503]), .A2(n10475), .B1(
        i_data_bus[407]), .B2(n10473), .ZN(n7353) );
  ND2D1BWP30P140LVT U10760 ( .A1(n7354), .A2(n7353), .ZN(N10612) );
  AOI22D1BWP30P140LVT U10761 ( .A1(i_data_bus[496]), .A2(n10475), .B1(
        i_data_bus[432]), .B2(n10474), .ZN(n7356) );
  AOI22D1BWP30P140LVT U10762 ( .A1(i_data_bus[464]), .A2(n10476), .B1(
        i_data_bus[400]), .B2(n10473), .ZN(n7355) );
  ND2D1BWP30P140LVT U10763 ( .A1(n7356), .A2(n7355), .ZN(N10605) );
  AOI22D1BWP30P140LVT U10764 ( .A1(i_data_bus[172]), .A2(n10515), .B1(
        i_data_bus[140]), .B2(n10513), .ZN(n7358) );
  AOI22D1BWP30P140LVT U10765 ( .A1(i_data_bus[236]), .A2(n10516), .B1(
        i_data_bus[204]), .B2(n10514), .ZN(n7357) );
  ND2D1BWP30P140LVT U10766 ( .A1(n7358), .A2(n7357), .ZN(N8295) );
  AOI22D1BWP30P140LVT U10767 ( .A1(i_data_bus[167]), .A2(n10515), .B1(
        i_data_bus[135]), .B2(n10513), .ZN(n7360) );
  AOI22D1BWP30P140LVT U10768 ( .A1(i_data_bus[231]), .A2(n10516), .B1(
        i_data_bus[199]), .B2(n10514), .ZN(n7359) );
  ND2D1BWP30P140LVT U10769 ( .A1(n7360), .A2(n7359), .ZN(N8290) );
  AOI22D1BWP30P140LVT U10770 ( .A1(i_data_bus[238]), .A2(n10516), .B1(
        i_data_bus[142]), .B2(n10513), .ZN(n7362) );
  AOI22D1BWP30P140LVT U10771 ( .A1(i_data_bus[174]), .A2(n10515), .B1(
        i_data_bus[206]), .B2(n10514), .ZN(n7361) );
  ND2D1BWP30P140LVT U10772 ( .A1(n7362), .A2(n7361), .ZN(N8297) );
  AOI22D1BWP30P140LVT U10773 ( .A1(i_data_bus[372]), .A2(n10416), .B1(
        i_data_bus[276]), .B2(n10415), .ZN(n7364) );
  AOI22D1BWP30P140LVT U10774 ( .A1(i_data_bus[308]), .A2(n10414), .B1(
        i_data_bus[340]), .B2(n10413), .ZN(n7363) );
  ND2D1BWP30P140LVT U10775 ( .A1(n7364), .A2(n7363), .ZN(N14141) );
  AOI22D1BWP30P140LVT U10776 ( .A1(i_data_bus[355]), .A2(n10416), .B1(
        i_data_bus[259]), .B2(n10415), .ZN(n7366) );
  AOI22D1BWP30P140LVT U10777 ( .A1(i_data_bus[291]), .A2(n10414), .B1(
        i_data_bus[323]), .B2(n10413), .ZN(n7365) );
  ND2D1BWP30P140LVT U10778 ( .A1(n7366), .A2(n7365), .ZN(N14124) );
  AOI22D1BWP30P140LVT U10779 ( .A1(i_data_bus[284]), .A2(n10415), .B1(
        i_data_bus[316]), .B2(n10414), .ZN(n7368) );
  AOI22D1BWP30P140LVT U10780 ( .A1(i_data_bus[380]), .A2(n10416), .B1(
        i_data_bus[348]), .B2(n10413), .ZN(n7367) );
  ND2D1BWP30P140LVT U10781 ( .A1(n7368), .A2(n7367), .ZN(N14149) );
  AOI22D1BWP30P140LVT U10782 ( .A1(i_data_bus[353]), .A2(n10416), .B1(
        i_data_bus[289]), .B2(n10414), .ZN(n7370) );
  AOI22D1BWP30P140LVT U10783 ( .A1(i_data_bus[257]), .A2(n10415), .B1(
        i_data_bus[321]), .B2(n10413), .ZN(n7369) );
  ND2D1BWP30P140LVT U10784 ( .A1(n7370), .A2(n7369), .ZN(N14122) );
  AOI22D1BWP30P140LVT U10785 ( .A1(i_data_bus[217]), .A2(n10514), .B1(
        i_data_bus[153]), .B2(n10513), .ZN(n7372) );
  AOI22D1BWP30P140LVT U10786 ( .A1(i_data_bus[249]), .A2(n10516), .B1(
        i_data_bus[185]), .B2(n10515), .ZN(n7371) );
  ND2D1BWP30P140LVT U10787 ( .A1(n7372), .A2(n7371), .ZN(N8308) );
  AOI22D1BWP30P140LVT U10788 ( .A1(i_data_bus[958]), .A2(n10521), .B1(
        i_data_bus[926]), .B2(n10524), .ZN(n7374) );
  AOI22D1BWP30P140LVT U10789 ( .A1(i_data_bus[990]), .A2(n10522), .B1(
        i_data_bus[1022]), .B2(n10523), .ZN(n7373) );
  ND2D1BWP30P140LVT U10790 ( .A1(n7374), .A2(n7373), .ZN(N7735) );
  AOI22D1BWP30P140LVT U10791 ( .A1(i_data_bus[216]), .A2(n10578), .B1(
        i_data_bus[152]), .B2(n10577), .ZN(n7376) );
  AOI22D1BWP30P140LVT U10792 ( .A1(i_data_bus[248]), .A2(n10580), .B1(
        i_data_bus[184]), .B2(n10579), .ZN(n7375) );
  ND2D1BWP30P140LVT U10793 ( .A1(n7376), .A2(n7375), .ZN(N4559) );
  AOI22D1BWP30P140LVT U10794 ( .A1(i_data_bus[979]), .A2(n10522), .B1(
        i_data_bus[915]), .B2(n10524), .ZN(n7378) );
  AOI22D1BWP30P140LVT U10795 ( .A1(i_data_bus[947]), .A2(n10521), .B1(
        i_data_bus[1011]), .B2(n10523), .ZN(n7377) );
  ND2D1BWP30P140LVT U10796 ( .A1(n7378), .A2(n7377), .ZN(N7724) );
  AOI22D1BWP30P140LVT U10797 ( .A1(i_data_bus[253]), .A2(n10580), .B1(
        i_data_bus[157]), .B2(n10577), .ZN(n7380) );
  AOI22D1BWP30P140LVT U10798 ( .A1(i_data_bus[221]), .A2(n10578), .B1(
        i_data_bus[189]), .B2(n10579), .ZN(n7379) );
  ND2D1BWP30P140LVT U10799 ( .A1(n7380), .A2(n7379), .ZN(N4564) );
  AOI22D1BWP30P140LVT U10800 ( .A1(i_data_bus[954]), .A2(n10521), .B1(
        i_data_bus[922]), .B2(n10524), .ZN(n7382) );
  AOI22D1BWP30P140LVT U10801 ( .A1(i_data_bus[986]), .A2(n10522), .B1(
        i_data_bus[1018]), .B2(n10523), .ZN(n7381) );
  ND2D1BWP30P140LVT U10802 ( .A1(n7382), .A2(n7381), .ZN(N7731) );
  AOI22D1BWP30P140LVT U10803 ( .A1(i_data_bus[921]), .A2(n10524), .B1(
        i_data_bus[953]), .B2(n10521), .ZN(n7384) );
  AOI22D1BWP30P140LVT U10804 ( .A1(i_data_bus[985]), .A2(n10522), .B1(
        i_data_bus[1017]), .B2(n10523), .ZN(n7383) );
  ND2D1BWP30P140LVT U10805 ( .A1(n7384), .A2(n7383), .ZN(N7730) );
  AOI22D1BWP30P140LVT U10806 ( .A1(i_data_bus[199]), .A2(n10578), .B1(
        i_data_bus[135]), .B2(n10577), .ZN(n7386) );
  AOI22D1BWP30P140LVT U10807 ( .A1(i_data_bus[231]), .A2(n10580), .B1(
        i_data_bus[167]), .B2(n10579), .ZN(n7385) );
  ND2D1BWP30P140LVT U10808 ( .A1(n7386), .A2(n7385), .ZN(N4542) );
  AOI22D1BWP30P140LVT U10809 ( .A1(i_data_bus[235]), .A2(n10580), .B1(
        i_data_bus[139]), .B2(n10577), .ZN(n7388) );
  AOI22D1BWP30P140LVT U10810 ( .A1(i_data_bus[203]), .A2(n10578), .B1(
        i_data_bus[171]), .B2(n10579), .ZN(n7387) );
  ND2D1BWP30P140LVT U10811 ( .A1(n7388), .A2(n7387), .ZN(N4546) );
  AOI22D1BWP30P140LVT U10812 ( .A1(i_data_bus[288]), .A2(n10414), .B1(
        i_data_bus[320]), .B2(n10413), .ZN(n7390) );
  AOI22D1BWP30P140LVT U10813 ( .A1(i_data_bus[352]), .A2(n10416), .B1(
        i_data_bus[256]), .B2(n10415), .ZN(n7389) );
  ND2D1BWP30P140LVT U10814 ( .A1(n7390), .A2(n7389), .ZN(N14121) );
  AOI22D1BWP30P140LVT U10815 ( .A1(i_data_bus[325]), .A2(n10413), .B1(
        i_data_bus[293]), .B2(n10414), .ZN(n7392) );
  AOI22D1BWP30P140LVT U10816 ( .A1(i_data_bus[357]), .A2(n10416), .B1(
        i_data_bus[261]), .B2(n10415), .ZN(n7391) );
  ND2D1BWP30P140LVT U10817 ( .A1(n7392), .A2(n7391), .ZN(N14126) );
  AOI22D1BWP30P140LVT U10818 ( .A1(i_data_bus[1003]), .A2(n10427), .B1(
        i_data_bus[971]), .B2(n10426), .ZN(n7394) );
  AOI22D1BWP30P140LVT U10819 ( .A1(i_data_bus[939]), .A2(n10428), .B1(
        i_data_bus[907]), .B2(n10425), .ZN(n7393) );
  ND2D1BWP30P140LVT U10820 ( .A1(n7394), .A2(n7393), .ZN(N13338) );
  AOI22D1BWP30P140LVT U10821 ( .A1(i_data_bus[350]), .A2(n10413), .B1(
        i_data_bus[318]), .B2(n10414), .ZN(n7396) );
  AOI22D1BWP30P140LVT U10822 ( .A1(i_data_bus[382]), .A2(n10416), .B1(
        i_data_bus[286]), .B2(n10415), .ZN(n7395) );
  ND2D1BWP30P140LVT U10823 ( .A1(n7396), .A2(n7395), .ZN(N14151) );
  AOI22D1BWP30P140LVT U10824 ( .A1(i_data_bus[338]), .A2(n10413), .B1(
        i_data_bus[306]), .B2(n10414), .ZN(n7398) );
  AOI22D1BWP30P140LVT U10825 ( .A1(i_data_bus[370]), .A2(n10416), .B1(
        i_data_bus[274]), .B2(n10415), .ZN(n7397) );
  ND2D1BWP30P140LVT U10826 ( .A1(n7398), .A2(n7397), .ZN(N14139) );
  AOI22D1BWP30P140LVT U10827 ( .A1(i_data_bus[932]), .A2(n10428), .B1(
        i_data_bus[964]), .B2(n10426), .ZN(n7400) );
  AOI22D1BWP30P140LVT U10828 ( .A1(i_data_bus[996]), .A2(n10427), .B1(
        i_data_bus[900]), .B2(n10425), .ZN(n7399) );
  ND2D1BWP30P140LVT U10829 ( .A1(n7400), .A2(n7399), .ZN(N13331) );
  AOI22D1BWP30P140LVT U10830 ( .A1(i_data_bus[294]), .A2(n10414), .B1(
        i_data_bus[326]), .B2(n10413), .ZN(n7402) );
  AOI22D1BWP30P140LVT U10831 ( .A1(i_data_bus[358]), .A2(n10416), .B1(
        i_data_bus[262]), .B2(n10415), .ZN(n7401) );
  ND2D1BWP30P140LVT U10832 ( .A1(n7402), .A2(n7401), .ZN(N14127) );
  AOI22D1BWP30P140LVT U10833 ( .A1(i_data_bus[945]), .A2(n10428), .B1(
        i_data_bus[977]), .B2(n10426), .ZN(n7404) );
  AOI22D1BWP30P140LVT U10834 ( .A1(i_data_bus[1009]), .A2(n10427), .B1(
        i_data_bus[913]), .B2(n10425), .ZN(n7403) );
  ND2D1BWP30P140LVT U10835 ( .A1(n7404), .A2(n7403), .ZN(N13344) );
  AOI22D1BWP30P140LVT U10836 ( .A1(i_data_bus[1014]), .A2(n10427), .B1(
        i_data_bus[982]), .B2(n10426), .ZN(n7406) );
  AOI22D1BWP30P140LVT U10837 ( .A1(i_data_bus[950]), .A2(n10428), .B1(
        i_data_bus[918]), .B2(n10425), .ZN(n7405) );
  ND2D1BWP30P140LVT U10838 ( .A1(n7406), .A2(n7405), .ZN(N13349) );
  AOI22D1BWP30P140LVT U10839 ( .A1(i_data_bus[1023]), .A2(n10427), .B1(
        i_data_bus[991]), .B2(n10426), .ZN(n7408) );
  AOI22D1BWP30P140LVT U10840 ( .A1(i_data_bus[927]), .A2(n10425), .B1(
        i_data_bus[959]), .B2(n10428), .ZN(n7407) );
  ND2D1BWP30P140LVT U10841 ( .A1(n7408), .A2(n7407), .ZN(N13358) );
  AOI22D1BWP30P140LVT U10842 ( .A1(i_data_bus[898]), .A2(n10425), .B1(
        i_data_bus[962]), .B2(n10426), .ZN(n7410) );
  AOI22D1BWP30P140LVT U10843 ( .A1(i_data_bus[994]), .A2(n10427), .B1(
        i_data_bus[930]), .B2(n10428), .ZN(n7409) );
  ND2D1BWP30P140LVT U10844 ( .A1(n7410), .A2(n7409), .ZN(N13329) );
  AOI22D1BWP30P140LVT U10845 ( .A1(i_data_bus[908]), .A2(n10425), .B1(
        i_data_bus[972]), .B2(n10426), .ZN(n7412) );
  AOI22D1BWP30P140LVT U10846 ( .A1(i_data_bus[940]), .A2(n10428), .B1(
        i_data_bus[1004]), .B2(n10427), .ZN(n7411) );
  ND2D1BWP30P140LVT U10847 ( .A1(n7412), .A2(n7411), .ZN(N13339) );
  AOI22D1BWP30P140LVT U10848 ( .A1(i_data_bus[899]), .A2(n10425), .B1(
        i_data_bus[963]), .B2(n10426), .ZN(n7414) );
  AOI22D1BWP30P140LVT U10849 ( .A1(i_data_bus[995]), .A2(n10427), .B1(
        i_data_bus[931]), .B2(n10428), .ZN(n7413) );
  ND2D1BWP30P140LVT U10850 ( .A1(n7414), .A2(n7413), .ZN(N13330) );
  AOI22D1BWP30P140LVT U10851 ( .A1(i_data_bus[911]), .A2(n10425), .B1(
        i_data_bus[975]), .B2(n10426), .ZN(n7416) );
  AOI22D1BWP30P140LVT U10852 ( .A1(i_data_bus[943]), .A2(n10428), .B1(
        i_data_bus[1007]), .B2(n10427), .ZN(n7415) );
  ND2D1BWP30P140LVT U10853 ( .A1(n7416), .A2(n7415), .ZN(N13342) );
  AOI22D1BWP30P140LVT U10854 ( .A1(i_data_bus[1006]), .A2(n10427), .B1(
        i_data_bus[974]), .B2(n10426), .ZN(n7418) );
  AOI22D1BWP30P140LVT U10855 ( .A1(i_data_bus[910]), .A2(n10425), .B1(
        i_data_bus[942]), .B2(n10428), .ZN(n7417) );
  ND2D1BWP30P140LVT U10856 ( .A1(n7418), .A2(n7417), .ZN(N13341) );
  AOI22D1BWP30P140LVT U10857 ( .A1(i_data_bus[896]), .A2(n10425), .B1(
        i_data_bus[960]), .B2(n10426), .ZN(n7420) );
  AOI22D1BWP30P140LVT U10858 ( .A1(i_data_bus[992]), .A2(n10427), .B1(
        i_data_bus[928]), .B2(n10428), .ZN(n7419) );
  ND2D1BWP30P140LVT U10859 ( .A1(n7420), .A2(n7419), .ZN(N13327) );
  AOI22D1BWP30P140LVT U10860 ( .A1(i_data_bus[903]), .A2(n10425), .B1(
        i_data_bus[967]), .B2(n10426), .ZN(n7422) );
  AOI22D1BWP30P140LVT U10861 ( .A1(i_data_bus[935]), .A2(n10428), .B1(
        i_data_bus[999]), .B2(n10427), .ZN(n7421) );
  ND2D1BWP30P140LVT U10862 ( .A1(n7422), .A2(n7421), .ZN(N13334) );
  AOI22D1BWP30P140LVT U10863 ( .A1(i_data_bus[787]), .A2(n10493), .B1(
        i_data_bus[819]), .B2(n10496), .ZN(n7424) );
  AOI22D1BWP30P140LVT U10864 ( .A1(i_data_bus[883]), .A2(n10494), .B1(
        i_data_bus[851]), .B2(n10495), .ZN(n7423) );
  ND2D1BWP30P140LVT U10865 ( .A1(n7424), .A2(n7423), .ZN(N9382) );
  AOI22D1BWP30P140LVT U10866 ( .A1(i_data_bus[777]), .A2(n10493), .B1(
        i_data_bus[809]), .B2(n10496), .ZN(n7426) );
  AOI22D1BWP30P140LVT U10867 ( .A1(i_data_bus[841]), .A2(n10495), .B1(
        i_data_bus[873]), .B2(n10494), .ZN(n7425) );
  ND2D1BWP30P140LVT U10868 ( .A1(n7426), .A2(n7425), .ZN(N9372) );
  AOI22D1BWP30P140LVT U10869 ( .A1(i_data_bus[778]), .A2(n10493), .B1(
        i_data_bus[810]), .B2(n10496), .ZN(n7428) );
  AOI22D1BWP30P140LVT U10870 ( .A1(i_data_bus[842]), .A2(n10495), .B1(
        i_data_bus[874]), .B2(n10494), .ZN(n7427) );
  ND2D1BWP30P140LVT U10871 ( .A1(n7428), .A2(n7427), .ZN(N9373) );
  AOI22D1BWP30P140LVT U10872 ( .A1(i_data_bus[245]), .A2(n10449), .B1(
        i_data_bus[181]), .B2(n10450), .ZN(n7430) );
  AOI22D1BWP30P140LVT U10873 ( .A1(i_data_bus[149]), .A2(n10452), .B1(
        i_data_bus[213]), .B2(n10451), .ZN(n7429) );
  ND2D1BWP30P140LVT U10874 ( .A1(n7430), .A2(n7429), .ZN(N12052) );
  AOI22D1BWP30P140LVT U10875 ( .A1(i_data_bus[178]), .A2(n10450), .B1(
        i_data_bus[242]), .B2(n10449), .ZN(n7432) );
  AOI22D1BWP30P140LVT U10876 ( .A1(i_data_bus[146]), .A2(n10452), .B1(
        i_data_bus[210]), .B2(n10451), .ZN(n7431) );
  ND2D1BWP30P140LVT U10877 ( .A1(n7432), .A2(n7431), .ZN(N12049) );
  AOI22D1BWP30P140LVT U10878 ( .A1(i_data_bus[224]), .A2(n10449), .B1(
        i_data_bus[160]), .B2(n10450), .ZN(n7434) );
  AOI22D1BWP30P140LVT U10879 ( .A1(i_data_bus[128]), .A2(n10452), .B1(
        i_data_bus[192]), .B2(n10451), .ZN(n7433) );
  ND2D1BWP30P140LVT U10880 ( .A1(n7434), .A2(n7433), .ZN(N12031) );
  AOI22D1BWP30P140LVT U10881 ( .A1(i_data_bus[926]), .A2(n10492), .B1(
        i_data_bus[990]), .B2(n10490), .ZN(n7436) );
  AOI22D1BWP30P140LVT U10882 ( .A1(i_data_bus[958]), .A2(n10491), .B1(
        i_data_bus[1022]), .B2(n10489), .ZN(n7435) );
  ND2D1BWP30P140LVT U10883 ( .A1(n7436), .A2(n7435), .ZN(N9609) );
  AOI22D1BWP30P140LVT U10884 ( .A1(i_data_bus[848]), .A2(n10590), .B1(
        i_data_bus[816]), .B2(n10592), .ZN(n7438) );
  AOI22D1BWP30P140LVT U10885 ( .A1(i_data_bus[784]), .A2(n10589), .B1(
        i_data_bus[880]), .B2(n10591), .ZN(n7437) );
  ND2D1BWP30P140LVT U10886 ( .A1(n7438), .A2(n7437), .ZN(N3757) );
  AOI22D1BWP30P140LVT U10887 ( .A1(i_data_bus[784]), .A2(n10558), .B1(
        i_data_bus[816]), .B2(n10560), .ZN(n7440) );
  AOI22D1BWP30P140LVT U10888 ( .A1(i_data_bus[848]), .A2(n10557), .B1(
        i_data_bus[880]), .B2(n10559), .ZN(n7439) );
  ND2D1BWP30P140LVT U10889 ( .A1(n7440), .A2(n7439), .ZN(N5631) );
  AOI22D1BWP30P140LVT U10890 ( .A1(i_data_bus[955]), .A2(n10491), .B1(
        i_data_bus[987]), .B2(n10490), .ZN(n7442) );
  AOI22D1BWP30P140LVT U10891 ( .A1(i_data_bus[923]), .A2(n10492), .B1(
        i_data_bus[1019]), .B2(n10489), .ZN(n7441) );
  ND2D1BWP30P140LVT U10892 ( .A1(n7442), .A2(n7441), .ZN(N9606) );
  AOI22D1BWP30P140LVT U10893 ( .A1(i_data_bus[796]), .A2(n10558), .B1(
        i_data_bus[828]), .B2(n10560), .ZN(n7444) );
  AOI22D1BWP30P140LVT U10894 ( .A1(i_data_bus[860]), .A2(n10557), .B1(
        i_data_bus[892]), .B2(n10559), .ZN(n7443) );
  ND2D1BWP30P140LVT U10895 ( .A1(n7444), .A2(n7443), .ZN(N5643) );
  AOI22D1BWP30P140LVT U10896 ( .A1(i_data_bus[920]), .A2(n10492), .B1(
        i_data_bus[984]), .B2(n10490), .ZN(n7446) );
  AOI22D1BWP30P140LVT U10897 ( .A1(i_data_bus[952]), .A2(n10491), .B1(
        i_data_bus[1016]), .B2(n10489), .ZN(n7445) );
  ND2D1BWP30P140LVT U10898 ( .A1(n7446), .A2(n7445), .ZN(N9603) );
  AOI22D1BWP30P140LVT U10899 ( .A1(i_data_bus[908]), .A2(n10492), .B1(
        i_data_bus[972]), .B2(n10490), .ZN(n7448) );
  AOI22D1BWP30P140LVT U10900 ( .A1(i_data_bus[940]), .A2(n10491), .B1(
        i_data_bus[1004]), .B2(n10489), .ZN(n7447) );
  ND2D1BWP30P140LVT U10901 ( .A1(n7448), .A2(n7447), .ZN(N9591) );
  AOI22D1BWP30P140LVT U10902 ( .A1(i_data_bus[779]), .A2(n10558), .B1(
        i_data_bus[811]), .B2(n10560), .ZN(n7450) );
  AOI22D1BWP30P140LVT U10903 ( .A1(i_data_bus[843]), .A2(n10557), .B1(
        i_data_bus[875]), .B2(n10559), .ZN(n7449) );
  ND2D1BWP30P140LVT U10904 ( .A1(n7450), .A2(n7449), .ZN(N5626) );
  AOI22D1BWP30P140LVT U10905 ( .A1(i_data_bus[104]), .A2(n10488), .B1(
        i_data_bus[72]), .B2(n10487), .ZN(n7452) );
  AOI22D1BWP30P140LVT U10906 ( .A1(i_data_bus[40]), .A2(n10485), .B1(
        i_data_bus[8]), .B2(n10486), .ZN(n7451) );
  ND2D1BWP30P140LVT U10907 ( .A1(n7452), .A2(n7451), .ZN(N9949) );
  AOI22D1BWP30P140LVT U10908 ( .A1(i_data_bus[798]), .A2(n10589), .B1(
        i_data_bus[830]), .B2(n10592), .ZN(n7454) );
  AOI22D1BWP30P140LVT U10909 ( .A1(i_data_bus[862]), .A2(n10590), .B1(
        i_data_bus[894]), .B2(n10591), .ZN(n7453) );
  ND2D1BWP30P140LVT U10910 ( .A1(n7454), .A2(n7453), .ZN(N3771) );
  AOI22D1BWP30P140LVT U10911 ( .A1(i_data_bus[780]), .A2(n10589), .B1(
        i_data_bus[812]), .B2(n10592), .ZN(n7456) );
  AOI22D1BWP30P140LVT U10912 ( .A1(i_data_bus[844]), .A2(n10590), .B1(
        i_data_bus[876]), .B2(n10591), .ZN(n7455) );
  ND2D1BWP30P140LVT U10913 ( .A1(n7456), .A2(n7455), .ZN(N3753) );
  AOI22D1BWP30P140LVT U10914 ( .A1(i_data_bus[772]), .A2(n10558), .B1(
        i_data_bus[804]), .B2(n10560), .ZN(n7458) );
  AOI22D1BWP30P140LVT U10915 ( .A1(i_data_bus[836]), .A2(n10557), .B1(
        i_data_bus[868]), .B2(n10559), .ZN(n7457) );
  ND2D1BWP30P140LVT U10916 ( .A1(n7458), .A2(n7457), .ZN(N5619) );
  AOI22D1BWP30P140LVT U10917 ( .A1(i_data_bus[995]), .A2(n10489), .B1(
        i_data_bus[963]), .B2(n10490), .ZN(n7460) );
  AOI22D1BWP30P140LVT U10918 ( .A1(i_data_bus[899]), .A2(n10492), .B1(
        i_data_bus[931]), .B2(n10491), .ZN(n7459) );
  ND2D1BWP30P140LVT U10919 ( .A1(n7460), .A2(n7459), .ZN(N9582) );
  AOI22D1BWP30P140LVT U10920 ( .A1(i_data_bus[992]), .A2(n10489), .B1(
        i_data_bus[960]), .B2(n10490), .ZN(n7462) );
  AOI22D1BWP30P140LVT U10921 ( .A1(i_data_bus[896]), .A2(n10492), .B1(
        i_data_bus[928]), .B2(n10491), .ZN(n7461) );
  ND2D1BWP30P140LVT U10922 ( .A1(n7462), .A2(n7461), .ZN(N9579) );
  AOI22D1BWP30P140LVT U10923 ( .A1(i_data_bus[1015]), .A2(n10489), .B1(
        i_data_bus[983]), .B2(n10490), .ZN(n7464) );
  AOI22D1BWP30P140LVT U10924 ( .A1(i_data_bus[919]), .A2(n10492), .B1(
        i_data_bus[951]), .B2(n10491), .ZN(n7463) );
  ND2D1BWP30P140LVT U10925 ( .A1(n7464), .A2(n7463), .ZN(N9602) );
  AOI22D1BWP30P140LVT U10926 ( .A1(i_data_bus[927]), .A2(n10492), .B1(
        i_data_bus[991]), .B2(n10490), .ZN(n7466) );
  AOI22D1BWP30P140LVT U10927 ( .A1(i_data_bus[1023]), .A2(n10489), .B1(
        i_data_bus[959]), .B2(n10491), .ZN(n7465) );
  ND2D1BWP30P140LVT U10928 ( .A1(n7466), .A2(n7465), .ZN(N9610) );
  AOI22D1BWP30P140LVT U10929 ( .A1(i_data_bus[82]), .A2(n10454), .B1(
        i_data_bus[18]), .B2(n10456), .ZN(n7468) );
  AOI22D1BWP30P140LVT U10930 ( .A1(i_data_bus[114]), .A2(n10455), .B1(
        i_data_bus[50]), .B2(n10453), .ZN(n7467) );
  ND2D1BWP30P140LVT U10931 ( .A1(n7468), .A2(n7467), .ZN(N11833) );
  AOI22D1BWP30P140LVT U10932 ( .A1(i_data_bus[65]), .A2(n10454), .B1(
        i_data_bus[1]), .B2(n10456), .ZN(n7470) );
  AOI22D1BWP30P140LVT U10933 ( .A1(i_data_bus[33]), .A2(n10453), .B1(
        i_data_bus[97]), .B2(n10455), .ZN(n7469) );
  ND2D1BWP30P140LVT U10934 ( .A1(n7470), .A2(n7469), .ZN(N11816) );
  AOI22D1BWP30P140LVT U10935 ( .A1(i_data_bus[69]), .A2(n10454), .B1(
        i_data_bus[5]), .B2(n10456), .ZN(n7472) );
  AOI22D1BWP30P140LVT U10936 ( .A1(i_data_bus[37]), .A2(n10453), .B1(
        i_data_bus[101]), .B2(n10455), .ZN(n7471) );
  ND2D1BWP30P140LVT U10937 ( .A1(n7472), .A2(n7471), .ZN(N11820) );
  AOI22D1BWP30P140LVT U10938 ( .A1(i_data_bus[39]), .A2(n10453), .B1(
        i_data_bus[7]), .B2(n10456), .ZN(n7474) );
  AOI22D1BWP30P140LVT U10939 ( .A1(i_data_bus[71]), .A2(n10454), .B1(
        i_data_bus[103]), .B2(n10455), .ZN(n7473) );
  ND2D1BWP30P140LVT U10940 ( .A1(n7474), .A2(n7473), .ZN(N11822) );
  AOI22D1BWP30P140LVT U10941 ( .A1(i_data_bus[75]), .A2(n10454), .B1(
        i_data_bus[11]), .B2(n10456), .ZN(n7476) );
  AOI22D1BWP30P140LVT U10942 ( .A1(i_data_bus[43]), .A2(n10453), .B1(
        i_data_bus[107]), .B2(n10455), .ZN(n7475) );
  ND2D1BWP30P140LVT U10943 ( .A1(n7476), .A2(n7475), .ZN(N11826) );
  AOI22D1BWP30P140LVT U10944 ( .A1(i_data_bus[120]), .A2(n10549), .B1(
        i_data_bus[88]), .B2(n10551), .ZN(n7478) );
  AOI22D1BWP30P140LVT U10945 ( .A1(i_data_bus[24]), .A2(n10552), .B1(
        i_data_bus[56]), .B2(n10550), .ZN(n7477) );
  ND2D1BWP30P140LVT U10946 ( .A1(n7478), .A2(n7477), .ZN(N6217) );
  AOI22D1BWP30P140LVT U10947 ( .A1(i_data_bus[73]), .A2(n10551), .B1(
        i_data_bus[105]), .B2(n10549), .ZN(n7480) );
  AOI22D1BWP30P140LVT U10948 ( .A1(i_data_bus[9]), .A2(n10552), .B1(
        i_data_bus[41]), .B2(n10550), .ZN(n7479) );
  ND2D1BWP30P140LVT U10949 ( .A1(n7480), .A2(n7479), .ZN(N6202) );
  AOI22D1BWP30P140LVT U10950 ( .A1(i_data_bus[23]), .A2(n10552), .B1(
        i_data_bus[119]), .B2(n10549), .ZN(n7482) );
  AOI22D1BWP30P140LVT U10951 ( .A1(i_data_bus[87]), .A2(n10551), .B1(
        i_data_bus[55]), .B2(n10550), .ZN(n7481) );
  ND2D1BWP30P140LVT U10952 ( .A1(n7482), .A2(n7481), .ZN(N6216) );
  AOI22D1BWP30P140LVT U10953 ( .A1(i_data_bus[571]), .A2(n10598), .B1(
        i_data_bus[603]), .B2(n10600), .ZN(n7484) );
  AOI22D1BWP30P140LVT U10954 ( .A1(i_data_bus[635]), .A2(n10599), .B1(
        i_data_bus[539]), .B2(n10597), .ZN(n7483) );
  ND2D1BWP30P140LVT U10955 ( .A1(n7484), .A2(n7483), .ZN(N3336) );
  AOI22D1BWP30P140LVT U10956 ( .A1(i_data_bus[564]), .A2(n10598), .B1(
        i_data_bus[596]), .B2(n10600), .ZN(n7486) );
  AOI22D1BWP30P140LVT U10957 ( .A1(i_data_bus[628]), .A2(n10599), .B1(
        i_data_bus[532]), .B2(n10597), .ZN(n7485) );
  ND2D1BWP30P140LVT U10958 ( .A1(n7486), .A2(n7485), .ZN(N3329) );
  AOI22D1BWP30P140LVT U10959 ( .A1(i_data_bus[626]), .A2(n10599), .B1(
        i_data_bus[562]), .B2(n10598), .ZN(n7488) );
  AOI22D1BWP30P140LVT U10960 ( .A1(i_data_bus[594]), .A2(n10600), .B1(
        i_data_bus[530]), .B2(n10597), .ZN(n7487) );
  ND2D1BWP30P140LVT U10961 ( .A1(n7488), .A2(n7487), .ZN(N3327) );
  AOI22D1BWP30P140LVT U10962 ( .A1(i_data_bus[616]), .A2(n10599), .B1(
        i_data_bus[584]), .B2(n10600), .ZN(n7490) );
  AOI22D1BWP30P140LVT U10963 ( .A1(i_data_bus[552]), .A2(n10598), .B1(
        i_data_bus[520]), .B2(n10597), .ZN(n7489) );
  ND2D1BWP30P140LVT U10964 ( .A1(n7490), .A2(n7489), .ZN(N3317) );
  AOI22D1BWP30P140LVT U10965 ( .A1(i_data_bus[631]), .A2(n10599), .B1(
        i_data_bus[567]), .B2(n10598), .ZN(n7492) );
  AOI22D1BWP30P140LVT U10966 ( .A1(i_data_bus[599]), .A2(n10600), .B1(
        i_data_bus[535]), .B2(n10597), .ZN(n7491) );
  ND2D1BWP30P140LVT U10967 ( .A1(n7492), .A2(n7491), .ZN(N3332) );
  AOI22D1BWP30P140LVT U10968 ( .A1(i_data_bus[179]), .A2(n10483), .B1(
        i_data_bus[243]), .B2(n10484), .ZN(n7494) );
  AOI22D1BWP30P140LVT U10969 ( .A1(i_data_bus[147]), .A2(n10481), .B1(
        i_data_bus[211]), .B2(n10482), .ZN(n7493) );
  ND2D1BWP30P140LVT U10970 ( .A1(n7494), .A2(n7493), .ZN(N10176) );
  AOI22D1BWP30P140LVT U10971 ( .A1(i_data_bus[172]), .A2(n10483), .B1(
        i_data_bus[140]), .B2(n10481), .ZN(n7496) );
  AOI22D1BWP30P140LVT U10972 ( .A1(i_data_bus[236]), .A2(n10484), .B1(
        i_data_bus[204]), .B2(n10482), .ZN(n7495) );
  ND2D1BWP30P140LVT U10973 ( .A1(n7496), .A2(n7495), .ZN(N10169) );
  AOI22D1BWP30P140LVT U10974 ( .A1(i_data_bus[149]), .A2(n10481), .B1(
        i_data_bus[181]), .B2(n10483), .ZN(n7498) );
  AOI22D1BWP30P140LVT U10975 ( .A1(i_data_bus[245]), .A2(n10484), .B1(
        i_data_bus[213]), .B2(n10482), .ZN(n7497) );
  ND2D1BWP30P140LVT U10976 ( .A1(n7498), .A2(n7497), .ZN(N10178) );
  AOI22D1BWP30P140LVT U10977 ( .A1(i_data_bus[44]), .A2(n10485), .B1(
        i_data_bus[12]), .B2(n10486), .ZN(n7500) );
  AOI22D1BWP30P140LVT U10978 ( .A1(i_data_bus[76]), .A2(n10487), .B1(
        i_data_bus[108]), .B2(n10488), .ZN(n7499) );
  ND2D1BWP30P140LVT U10979 ( .A1(n7500), .A2(n7499), .ZN(N9953) );
  AOI22D1BWP30P140LVT U10980 ( .A1(i_data_bus[154]), .A2(n10481), .B1(
        i_data_bus[250]), .B2(n10484), .ZN(n7502) );
  AOI22D1BWP30P140LVT U10981 ( .A1(i_data_bus[186]), .A2(n10483), .B1(
        i_data_bus[218]), .B2(n10482), .ZN(n7501) );
  ND2D1BWP30P140LVT U10982 ( .A1(n7502), .A2(n7501), .ZN(N10183) );
  AOI22D1BWP30P140LVT U10983 ( .A1(i_data_bus[37]), .A2(n10485), .B1(
        i_data_bus[69]), .B2(n10487), .ZN(n7504) );
  AOI22D1BWP30P140LVT U10984 ( .A1(i_data_bus[5]), .A2(n10486), .B1(
        i_data_bus[101]), .B2(n10488), .ZN(n7503) );
  ND2D1BWP30P140LVT U10985 ( .A1(n7504), .A2(n7503), .ZN(N9946) );
  AOI22D1BWP30P140LVT U10986 ( .A1(i_data_bus[132]), .A2(n10481), .B1(
        i_data_bus[164]), .B2(n10483), .ZN(n7506) );
  AOI22D1BWP30P140LVT U10987 ( .A1(i_data_bus[228]), .A2(n10484), .B1(
        i_data_bus[196]), .B2(n10482), .ZN(n7505) );
  ND2D1BWP30P140LVT U10988 ( .A1(n7506), .A2(n7505), .ZN(N10161) );
  AOI22D1BWP30P140LVT U10989 ( .A1(i_data_bus[71]), .A2(n10487), .B1(
        i_data_bus[7]), .B2(n10486), .ZN(n7508) );
  AOI22D1BWP30P140LVT U10990 ( .A1(i_data_bus[39]), .A2(n10485), .B1(
        i_data_bus[103]), .B2(n10488), .ZN(n7507) );
  ND2D1BWP30P140LVT U10991 ( .A1(n7508), .A2(n7507), .ZN(N9948) );
  AOI22D1BWP30P140LVT U10992 ( .A1(i_data_bus[61]), .A2(n10485), .B1(
        i_data_bus[29]), .B2(n10486), .ZN(n7510) );
  AOI22D1BWP30P140LVT U10993 ( .A1(i_data_bus[93]), .A2(n10487), .B1(
        i_data_bus[125]), .B2(n10488), .ZN(n7509) );
  ND2D1BWP30P140LVT U10994 ( .A1(n7510), .A2(n7509), .ZN(N9970) );
  AOI22D1BWP30P140LVT U10995 ( .A1(i_data_bus[133]), .A2(n10481), .B1(
        i_data_bus[229]), .B2(n10484), .ZN(n7512) );
  AOI22D1BWP30P140LVT U10996 ( .A1(i_data_bus[165]), .A2(n10483), .B1(
        i_data_bus[197]), .B2(n10482), .ZN(n7511) );
  ND2D1BWP30P140LVT U10997 ( .A1(n7512), .A2(n7511), .ZN(N10162) );
  AOI22D1BWP30P140LVT U10998 ( .A1(i_data_bus[163]), .A2(n10483), .B1(
        i_data_bus[131]), .B2(n10481), .ZN(n7514) );
  AOI22D1BWP30P140LVT U10999 ( .A1(i_data_bus[227]), .A2(n10484), .B1(
        i_data_bus[195]), .B2(n10482), .ZN(n7513) );
  ND2D1BWP30P140LVT U11000 ( .A1(n7514), .A2(n7513), .ZN(N10160) );
  AOI22D1BWP30P140LVT U11001 ( .A1(i_data_bus[183]), .A2(n10483), .B1(
        i_data_bus[247]), .B2(n10484), .ZN(n7516) );
  AOI22D1BWP30P140LVT U11002 ( .A1(i_data_bus[151]), .A2(n10481), .B1(
        i_data_bus[215]), .B2(n10482), .ZN(n7515) );
  ND2D1BWP30P140LVT U11003 ( .A1(n7516), .A2(n7515), .ZN(N10180) );
  AOI22D1BWP30P140LVT U11004 ( .A1(i_data_bus[86]), .A2(n10487), .B1(
        i_data_bus[22]), .B2(n10486), .ZN(n7518) );
  AOI22D1BWP30P140LVT U11005 ( .A1(i_data_bus[118]), .A2(n10488), .B1(
        i_data_bus[54]), .B2(n10485), .ZN(n7517) );
  ND2D1BWP30P140LVT U11006 ( .A1(n7518), .A2(n7517), .ZN(N9963) );
  AOI22D1BWP30P140LVT U11007 ( .A1(i_data_bus[117]), .A2(n10488), .B1(
        i_data_bus[85]), .B2(n10487), .ZN(n7520) );
  AOI22D1BWP30P140LVT U11008 ( .A1(i_data_bus[21]), .A2(n10486), .B1(
        i_data_bus[53]), .B2(n10485), .ZN(n7519) );
  ND2D1BWP30P140LVT U11009 ( .A1(n7520), .A2(n7519), .ZN(N9962) );
  AOI22D1BWP30P140LVT U11010 ( .A1(i_data_bus[24]), .A2(n10486), .B1(
        i_data_bus[88]), .B2(n10487), .ZN(n7522) );
  AOI22D1BWP30P140LVT U11011 ( .A1(i_data_bus[120]), .A2(n10488), .B1(
        i_data_bus[56]), .B2(n10485), .ZN(n7521) );
  ND2D1BWP30P140LVT U11012 ( .A1(n7522), .A2(n7521), .ZN(N9965) );
  AOI22D1BWP30P140LVT U11013 ( .A1(i_data_bus[119]), .A2(n10488), .B1(
        i_data_bus[87]), .B2(n10487), .ZN(n7524) );
  AOI22D1BWP30P140LVT U11014 ( .A1(i_data_bus[23]), .A2(n10486), .B1(
        i_data_bus[55]), .B2(n10485), .ZN(n7523) );
  ND2D1BWP30P140LVT U11015 ( .A1(n7524), .A2(n7523), .ZN(N9964) );
  AOI22D1BWP30P140LVT U11016 ( .A1(i_data_bus[89]), .A2(n10487), .B1(
        i_data_bus[25]), .B2(n10486), .ZN(n7526) );
  AOI22D1BWP30P140LVT U11017 ( .A1(i_data_bus[121]), .A2(n10488), .B1(
        i_data_bus[57]), .B2(n10485), .ZN(n7525) );
  ND2D1BWP30P140LVT U11018 ( .A1(n7526), .A2(n7525), .ZN(N9966) );
  AOI22D1BWP30P140LVT U11019 ( .A1(i_data_bus[98]), .A2(n10488), .B1(
        i_data_bus[2]), .B2(n10486), .ZN(n7528) );
  AOI22D1BWP30P140LVT U11020 ( .A1(i_data_bus[66]), .A2(n10487), .B1(
        i_data_bus[34]), .B2(n10485), .ZN(n7527) );
  ND2D1BWP30P140LVT U11021 ( .A1(n7528), .A2(n7527), .ZN(N9943) );
  AOI22D1BWP30P140LVT U11022 ( .A1(i_data_bus[111]), .A2(n10488), .B1(
        i_data_bus[79]), .B2(n10487), .ZN(n7530) );
  AOI22D1BWP30P140LVT U11023 ( .A1(i_data_bus[15]), .A2(n10486), .B1(
        i_data_bus[47]), .B2(n10485), .ZN(n7529) );
  ND2D1BWP30P140LVT U11024 ( .A1(n7530), .A2(n7529), .ZN(N9956) );
  AOI22D1BWP30P140LVT U11025 ( .A1(i_data_bus[74]), .A2(n10487), .B1(
        i_data_bus[106]), .B2(n10488), .ZN(n7532) );
  AOI22D1BWP30P140LVT U11026 ( .A1(i_data_bus[10]), .A2(n10486), .B1(
        i_data_bus[42]), .B2(n10485), .ZN(n7531) );
  ND2D1BWP30P140LVT U11027 ( .A1(n7532), .A2(n7531), .ZN(N9951) );
  AOI22D1BWP30P140LVT U11028 ( .A1(i_data_bus[496]), .A2(n10602), .B1(
        i_data_bus[432]), .B2(n10601), .ZN(n7534) );
  AOI22D1BWP30P140LVT U11029 ( .A1(i_data_bus[464]), .A2(n10604), .B1(
        i_data_bus[400]), .B2(n10603), .ZN(n7533) );
  ND2D1BWP30P140LVT U11030 ( .A1(n7534), .A2(n7533), .ZN(N3109) );
  AOI22D1BWP30P140LVT U11031 ( .A1(i_data_bus[482]), .A2(n10602), .B1(
        i_data_bus[418]), .B2(n10601), .ZN(n7536) );
  AOI22D1BWP30P140LVT U11032 ( .A1(i_data_bus[450]), .A2(n10604), .B1(
        i_data_bus[386]), .B2(n10603), .ZN(n7535) );
  ND2D1BWP30P140LVT U11033 ( .A1(n7536), .A2(n7535), .ZN(N3095) );
  AOI22D1BWP30P140LVT U11034 ( .A1(i_data_bus[474]), .A2(n10604), .B1(
        i_data_bus[442]), .B2(n10601), .ZN(n7538) );
  AOI22D1BWP30P140LVT U11035 ( .A1(i_data_bus[506]), .A2(n10602), .B1(
        i_data_bus[410]), .B2(n10603), .ZN(n7537) );
  ND2D1BWP30P140LVT U11036 ( .A1(n7538), .A2(n7537), .ZN(N3119) );
  AOI22D1BWP30P140LVT U11037 ( .A1(i_data_bus[457]), .A2(n10604), .B1(
        i_data_bus[425]), .B2(n10601), .ZN(n7540) );
  AOI22D1BWP30P140LVT U11038 ( .A1(i_data_bus[489]), .A2(n10602), .B1(
        i_data_bus[393]), .B2(n10603), .ZN(n7539) );
  ND2D1BWP30P140LVT U11039 ( .A1(n7540), .A2(n7539), .ZN(N3102) );
  AOI22D1BWP30P140LVT U11040 ( .A1(i_data_bus[444]), .A2(n10601), .B1(
        i_data_bus[508]), .B2(n10602), .ZN(n7542) );
  AOI22D1BWP30P140LVT U11041 ( .A1(i_data_bus[476]), .A2(n10604), .B1(
        i_data_bus[412]), .B2(n10603), .ZN(n7541) );
  ND2D1BWP30P140LVT U11042 ( .A1(n7542), .A2(n7541), .ZN(N3121) );
  AOI22D1BWP30P140LVT U11043 ( .A1(i_data_bus[460]), .A2(n10604), .B1(
        i_data_bus[428]), .B2(n10601), .ZN(n7544) );
  AOI22D1BWP30P140LVT U11044 ( .A1(i_data_bus[492]), .A2(n10602), .B1(
        i_data_bus[396]), .B2(n10603), .ZN(n7543) );
  ND2D1BWP30P140LVT U11045 ( .A1(n7544), .A2(n7543), .ZN(N3105) );
  AOI22D1BWP30P140LVT U11046 ( .A1(i_data_bus[174]), .A2(n10420), .B1(
        i_data_bus[142]), .B2(n10417), .ZN(n7546) );
  AOI22D1BWP30P140LVT U11047 ( .A1(i_data_bus[238]), .A2(n10418), .B1(
        i_data_bus[206]), .B2(n10419), .ZN(n7545) );
  ND2D1BWP30P140LVT U11048 ( .A1(n7546), .A2(n7545), .ZN(N13919) );
  AOI22D1BWP30P140LVT U11049 ( .A1(i_data_bus[187]), .A2(n10420), .B1(
        i_data_bus[155]), .B2(n10417), .ZN(n7548) );
  AOI22D1BWP30P140LVT U11050 ( .A1(i_data_bus[251]), .A2(n10418), .B1(
        i_data_bus[219]), .B2(n10419), .ZN(n7547) );
  ND2D1BWP30P140LVT U11051 ( .A1(n7548), .A2(n7547), .ZN(N13932) );
  AOI22D1BWP30P140LVT U11052 ( .A1(i_data_bus[186]), .A2(n10420), .B1(
        i_data_bus[154]), .B2(n10417), .ZN(n7550) );
  AOI22D1BWP30P140LVT U11053 ( .A1(i_data_bus[250]), .A2(n10418), .B1(
        i_data_bus[218]), .B2(n10419), .ZN(n7549) );
  ND2D1BWP30P140LVT U11054 ( .A1(n7550), .A2(n7549), .ZN(N13931) );
  AOI22D1BWP30P140LVT U11055 ( .A1(i_data_bus[531]), .A2(n10533), .B1(
        i_data_bus[627]), .B2(n10534), .ZN(n7552) );
  AOI22D1BWP30P140LVT U11056 ( .A1(i_data_bus[595]), .A2(n10536), .B1(
        i_data_bus[563]), .B2(n10535), .ZN(n7551) );
  ND2D1BWP30P140LVT U11057 ( .A1(n7552), .A2(n7551), .ZN(N7076) );
  AOI22D1BWP30P140LVT U11058 ( .A1(i_data_bus[928]), .A2(n10521), .B1(
        i_data_bus[960]), .B2(n10522), .ZN(n7554) );
  AOI22D1BWP30P140LVT U11059 ( .A1(i_data_bus[896]), .A2(n10524), .B1(
        i_data_bus[992]), .B2(n10523), .ZN(n7553) );
  ND2D1BWP30P140LVT U11060 ( .A1(n7554), .A2(n7553), .ZN(N7705) );
  AOI22D1BWP30P140LVT U11061 ( .A1(i_data_bus[1004]), .A2(n10523), .B1(
        i_data_bus[972]), .B2(n10522), .ZN(n7556) );
  AOI22D1BWP30P140LVT U11062 ( .A1(i_data_bus[908]), .A2(n10524), .B1(
        i_data_bus[940]), .B2(n10521), .ZN(n7555) );
  ND2D1BWP30P140LVT U11063 ( .A1(n7556), .A2(n7555), .ZN(N7717) );
  AOI22D1BWP30P140LVT U11064 ( .A1(i_data_bus[899]), .A2(n10524), .B1(
        i_data_bus[963]), .B2(n10522), .ZN(n7558) );
  AOI22D1BWP30P140LVT U11065 ( .A1(i_data_bus[995]), .A2(n10523), .B1(
        i_data_bus[931]), .B2(n10521), .ZN(n7557) );
  ND2D1BWP30P140LVT U11066 ( .A1(n7558), .A2(n7557), .ZN(N7708) );
  AOI22D1BWP30P140LVT U11067 ( .A1(i_data_bus[955]), .A2(n10521), .B1(
        i_data_bus[987]), .B2(n10522), .ZN(n7560) );
  AOI22D1BWP30P140LVT U11068 ( .A1(i_data_bus[923]), .A2(n10524), .B1(
        i_data_bus[1019]), .B2(n10523), .ZN(n7559) );
  ND2D1BWP30P140LVT U11069 ( .A1(n7560), .A2(n7559), .ZN(N7732) );
  AOI22D1BWP30P140LVT U11070 ( .A1(i_data_bus[549]), .A2(n10472), .B1(
        i_data_bus[613]), .B2(n10470), .ZN(n7562) );
  AOI22D1BWP30P140LVT U11071 ( .A1(i_data_bus[517]), .A2(n10471), .B1(
        i_data_bus[581]), .B2(n10469), .ZN(n7561) );
  ND2D1BWP30P140LVT U11072 ( .A1(n7562), .A2(n7561), .ZN(N10810) );
  AOI22D1BWP30P140LVT U11073 ( .A1(i_data_bus[552]), .A2(n10535), .B1(
        i_data_bus[616]), .B2(n10534), .ZN(n7564) );
  AOI22D1BWP30P140LVT U11074 ( .A1(i_data_bus[584]), .A2(n10536), .B1(
        i_data_bus[520]), .B2(n10533), .ZN(n7563) );
  ND2D1BWP30P140LVT U11075 ( .A1(n7564), .A2(n7563), .ZN(N7065) );
  AOI22D1BWP30P140LVT U11076 ( .A1(i_data_bus[602]), .A2(n10536), .B1(
        i_data_bus[634]), .B2(n10534), .ZN(n7566) );
  AOI22D1BWP30P140LVT U11077 ( .A1(i_data_bus[570]), .A2(n10535), .B1(
        i_data_bus[538]), .B2(n10533), .ZN(n7565) );
  ND2D1BWP30P140LVT U11078 ( .A1(n7566), .A2(n7565), .ZN(N7083) );
  AOI22D1BWP30P140LVT U11079 ( .A1(i_data_bus[558]), .A2(n10535), .B1(
        i_data_bus[622]), .B2(n10534), .ZN(n7568) );
  AOI22D1BWP30P140LVT U11080 ( .A1(i_data_bus[526]), .A2(n10533), .B1(
        i_data_bus[590]), .B2(n10536), .ZN(n7567) );
  ND2D1BWP30P140LVT U11081 ( .A1(n7568), .A2(n7567), .ZN(N7071) );
  AOI22D1BWP30P140LVT U11082 ( .A1(i_data_bus[527]), .A2(n10533), .B1(
        i_data_bus[623]), .B2(n10534), .ZN(n7570) );
  AOI22D1BWP30P140LVT U11083 ( .A1(i_data_bus[559]), .A2(n10535), .B1(
        i_data_bus[591]), .B2(n10536), .ZN(n7569) );
  ND2D1BWP30P140LVT U11084 ( .A1(n7570), .A2(n7569), .ZN(N7072) );
  AOI22D1BWP30P140LVT U11085 ( .A1(i_data_bus[549]), .A2(n10535), .B1(
        i_data_bus[613]), .B2(n10534), .ZN(n7572) );
  AOI22D1BWP30P140LVT U11086 ( .A1(i_data_bus[517]), .A2(n10533), .B1(
        i_data_bus[581]), .B2(n10536), .ZN(n7571) );
  ND2D1BWP30P140LVT U11087 ( .A1(n7572), .A2(n7571), .ZN(N7062) );
  AOI22D1BWP30P140LVT U11088 ( .A1(i_data_bus[695]), .A2(n10532), .B1(
        i_data_bus[727]), .B2(n10531), .ZN(n7574) );
  AOI22D1BWP30P140LVT U11089 ( .A1(i_data_bus[663]), .A2(n10529), .B1(
        i_data_bus[759]), .B2(n10530), .ZN(n7573) );
  ND2D1BWP30P140LVT U11090 ( .A1(n7574), .A2(n7573), .ZN(N7296) );
  AOI22D1BWP30P140LVT U11091 ( .A1(i_data_bus[681]), .A2(n10532), .B1(
        i_data_bus[649]), .B2(n10529), .ZN(n7576) );
  AOI22D1BWP30P140LVT U11092 ( .A1(i_data_bus[713]), .A2(n10531), .B1(
        i_data_bus[745]), .B2(n10530), .ZN(n7575) );
  ND2D1BWP30P140LVT U11093 ( .A1(n7576), .A2(n7575), .ZN(N7282) );
  AOI22D1BWP30P140LVT U11094 ( .A1(i_data_bus[700]), .A2(n10532), .B1(
        i_data_bus[668]), .B2(n10529), .ZN(n7578) );
  AOI22D1BWP30P140LVT U11095 ( .A1(i_data_bus[732]), .A2(n10531), .B1(
        i_data_bus[764]), .B2(n10530), .ZN(n7577) );
  ND2D1BWP30P140LVT U11096 ( .A1(n7578), .A2(n7577), .ZN(N7301) );
  AOI22D1BWP30P140LVT U11097 ( .A1(i_data_bus[660]), .A2(n10529), .B1(
        i_data_bus[724]), .B2(n10531), .ZN(n7580) );
  AOI22D1BWP30P140LVT U11098 ( .A1(i_data_bus[692]), .A2(n10532), .B1(
        i_data_bus[756]), .B2(n10530), .ZN(n7579) );
  ND2D1BWP30P140LVT U11099 ( .A1(n7580), .A2(n7579), .ZN(N7293) );
  AOI22D1BWP30P140LVT U11100 ( .A1(i_data_bus[696]), .A2(n10532), .B1(
        i_data_bus[664]), .B2(n10529), .ZN(n7582) );
  AOI22D1BWP30P140LVT U11101 ( .A1(i_data_bus[728]), .A2(n10531), .B1(
        i_data_bus[760]), .B2(n10530), .ZN(n7581) );
  ND2D1BWP30P140LVT U11102 ( .A1(n7582), .A2(n7581), .ZN(N7297) );
  AOI22D1BWP30P140LVT U11103 ( .A1(i_data_bus[710]), .A2(n10531), .B1(
        i_data_bus[678]), .B2(n10532), .ZN(n7584) );
  AOI22D1BWP30P140LVT U11104 ( .A1(i_data_bus[646]), .A2(n10529), .B1(
        i_data_bus[742]), .B2(n10530), .ZN(n7583) );
  ND2D1BWP30P140LVT U11105 ( .A1(n7584), .A2(n7583), .ZN(N7279) );
  AOI22D1BWP30P140LVT U11106 ( .A1(i_data_bus[121]), .A2(n10549), .B1(
        i_data_bus[25]), .B2(n10552), .ZN(n7586) );
  AOI22D1BWP30P140LVT U11107 ( .A1(i_data_bus[89]), .A2(n10551), .B1(
        i_data_bus[57]), .B2(n10550), .ZN(n7585) );
  ND2D1BWP30P140LVT U11108 ( .A1(n7586), .A2(n7585), .ZN(N6218) );
  AOI22D1BWP30P140LVT U11109 ( .A1(i_data_bus[39]), .A2(n10550), .B1(
        i_data_bus[7]), .B2(n10552), .ZN(n7588) );
  AOI22D1BWP30P140LVT U11110 ( .A1(i_data_bus[71]), .A2(n10551), .B1(
        i_data_bus[103]), .B2(n10549), .ZN(n7587) );
  ND2D1BWP30P140LVT U11111 ( .A1(n7588), .A2(n7587), .ZN(N6200) );
  AOI22D1BWP30P140LVT U11112 ( .A1(i_data_bus[75]), .A2(n10551), .B1(
        i_data_bus[11]), .B2(n10552), .ZN(n7590) );
  AOI22D1BWP30P140LVT U11113 ( .A1(i_data_bus[43]), .A2(n10550), .B1(
        i_data_bus[107]), .B2(n10549), .ZN(n7589) );
  ND2D1BWP30P140LVT U11114 ( .A1(n7590), .A2(n7589), .ZN(N6204) );
  AOI22D1BWP30P140LVT U11115 ( .A1(i_data_bus[98]), .A2(n10549), .B1(
        i_data_bus[2]), .B2(n10552), .ZN(n7592) );
  AOI22D1BWP30P140LVT U11116 ( .A1(i_data_bus[66]), .A2(n10551), .B1(
        i_data_bus[34]), .B2(n10550), .ZN(n7591) );
  ND2D1BWP30P140LVT U11117 ( .A1(n7592), .A2(n7591), .ZN(N6195) );
  AOI22D1BWP30P140LVT U11118 ( .A1(i_data_bus[127]), .A2(n10549), .B1(
        i_data_bus[31]), .B2(n10552), .ZN(n7594) );
  AOI22D1BWP30P140LVT U11119 ( .A1(i_data_bus[95]), .A2(n10551), .B1(
        i_data_bus[63]), .B2(n10550), .ZN(n7593) );
  ND2D1BWP30P140LVT U11120 ( .A1(n7594), .A2(n7593), .ZN(N6224) );
  AOI22D1BWP30P140LVT U11121 ( .A1(i_data_bus[1007]), .A2(n10393), .B1(
        i_data_bus[975]), .B2(n10396), .ZN(n7596) );
  AOI22D1BWP30P140LVT U11122 ( .A1(i_data_bus[943]), .A2(n10394), .B1(
        i_data_bus[911]), .B2(n10395), .ZN(n7595) );
  ND2D1BWP30P140LVT U11123 ( .A1(n7596), .A2(n7595), .ZN(N15216) );
  AOI22D1BWP30P140LVT U11124 ( .A1(i_data_bus[947]), .A2(n10394), .B1(
        i_data_bus[979]), .B2(n10396), .ZN(n7598) );
  AOI22D1BWP30P140LVT U11125 ( .A1(i_data_bus[1011]), .A2(n10393), .B1(
        i_data_bus[915]), .B2(n10395), .ZN(n7597) );
  ND2D1BWP30P140LVT U11126 ( .A1(n7598), .A2(n7597), .ZN(N15220) );
  AOI22D1BWP30P140LVT U11127 ( .A1(i_data_bus[903]), .A2(n10395), .B1(
        i_data_bus[967]), .B2(n10396), .ZN(n7600) );
  AOI22D1BWP30P140LVT U11128 ( .A1(i_data_bus[935]), .A2(n10394), .B1(
        i_data_bus[999]), .B2(n10393), .ZN(n7599) );
  ND2D1BWP30P140LVT U11129 ( .A1(n7600), .A2(n7599), .ZN(N15208) );
  AOI22D1BWP30P140LVT U11130 ( .A1(i_data_bus[958]), .A2(n10588), .B1(
        i_data_bus[1022]), .B2(n10585), .ZN(n7602) );
  AOI22D1BWP30P140LVT U11131 ( .A1(i_data_bus[926]), .A2(n10587), .B1(
        i_data_bus[990]), .B2(n10586), .ZN(n7601) );
  ND2D1BWP30P140LVT U11132 ( .A1(n7602), .A2(n7601), .ZN(N3987) );
  AOI22D1BWP30P140LVT U11133 ( .A1(i_data_bus[939]), .A2(n10588), .B1(
        i_data_bus[907]), .B2(n10587), .ZN(n7604) );
  AOI22D1BWP30P140LVT U11134 ( .A1(i_data_bus[1003]), .A2(n10585), .B1(
        i_data_bus[971]), .B2(n10586), .ZN(n7603) );
  ND2D1BWP30P140LVT U11135 ( .A1(n7604), .A2(n7603), .ZN(N3968) );
  AOI22D1BWP30P140LVT U11136 ( .A1(i_data_bus[1008]), .A2(n10585), .B1(
        i_data_bus[944]), .B2(n10588), .ZN(n7606) );
  AOI22D1BWP30P140LVT U11137 ( .A1(i_data_bus[912]), .A2(n10587), .B1(
        i_data_bus[976]), .B2(n10586), .ZN(n7605) );
  ND2D1BWP30P140LVT U11138 ( .A1(n7606), .A2(n7605), .ZN(N3973) );
  AOI22D1BWP30P140LVT U11139 ( .A1(i_data_bus[1014]), .A2(n10585), .B1(
        i_data_bus[918]), .B2(n10587), .ZN(n7608) );
  AOI22D1BWP30P140LVT U11140 ( .A1(i_data_bus[950]), .A2(n10588), .B1(
        i_data_bus[982]), .B2(n10586), .ZN(n7607) );
  ND2D1BWP30P140LVT U11141 ( .A1(n7608), .A2(n7607), .ZN(N3979) );
  AOI22D1BWP30P140LVT U11142 ( .A1(i_data_bus[934]), .A2(n10588), .B1(
        i_data_bus[902]), .B2(n10587), .ZN(n7610) );
  AOI22D1BWP30P140LVT U11143 ( .A1(i_data_bus[998]), .A2(n10585), .B1(
        i_data_bus[966]), .B2(n10586), .ZN(n7609) );
  ND2D1BWP30P140LVT U11144 ( .A1(n7610), .A2(n7609), .ZN(N3963) );
  AOI22D1BWP30P140LVT U11145 ( .A1(i_data_bus[1023]), .A2(n10585), .B1(
        i_data_bus[959]), .B2(n10588), .ZN(n7612) );
  AOI22D1BWP30P140LVT U11146 ( .A1(i_data_bus[927]), .A2(n10587), .B1(
        i_data_bus[991]), .B2(n10586), .ZN(n7611) );
  ND2D1BWP30P140LVT U11147 ( .A1(n7612), .A2(n7611), .ZN(N3988) );
  AOI22D1BWP30P140LVT U11148 ( .A1(i_data_bus[1023]), .A2(n10393), .B1(
        i_data_bus[991]), .B2(n10396), .ZN(n7614) );
  AOI22D1BWP30P140LVT U11149 ( .A1(i_data_bus[927]), .A2(n10395), .B1(
        i_data_bus[959]), .B2(n10394), .ZN(n7613) );
  ND2D1BWP30P140LVT U11150 ( .A1(n7614), .A2(n7613), .ZN(N15232) );
  AOI22D1BWP30P140LVT U11151 ( .A1(i_data_bus[943]), .A2(n10588), .B1(
        i_data_bus[1007]), .B2(n10585), .ZN(n7616) );
  AOI22D1BWP30P140LVT U11152 ( .A1(i_data_bus[911]), .A2(n10587), .B1(
        i_data_bus[975]), .B2(n10586), .ZN(n7615) );
  ND2D1BWP30P140LVT U11153 ( .A1(n7616), .A2(n7615), .ZN(N3972) );
  AOI22D1BWP30P140LVT U11154 ( .A1(i_data_bus[932]), .A2(n10588), .B1(
        i_data_bus[900]), .B2(n10587), .ZN(n7618) );
  AOI22D1BWP30P140LVT U11155 ( .A1(i_data_bus[996]), .A2(n10585), .B1(
        i_data_bus[964]), .B2(n10586), .ZN(n7617) );
  ND2D1BWP30P140LVT U11156 ( .A1(n7618), .A2(n7617), .ZN(N3961) );
  AOI22D1BWP30P140LVT U11157 ( .A1(i_data_bus[558]), .A2(n10567), .B1(
        i_data_bus[622]), .B2(n10568), .ZN(n7620) );
  AOI22D1BWP30P140LVT U11158 ( .A1(i_data_bus[526]), .A2(n10566), .B1(
        i_data_bus[590]), .B2(n10565), .ZN(n7619) );
  ND2D1BWP30P140LVT U11159 ( .A1(n7620), .A2(n7619), .ZN(N5197) );
  AOI22D1BWP30P140LVT U11160 ( .A1(i_data_bus[524]), .A2(n10566), .B1(
        i_data_bus[620]), .B2(n10568), .ZN(n7622) );
  AOI22D1BWP30P140LVT U11161 ( .A1(i_data_bus[556]), .A2(n10567), .B1(
        i_data_bus[588]), .B2(n10565), .ZN(n7621) );
  ND2D1BWP30P140LVT U11162 ( .A1(n7622), .A2(n7621), .ZN(N5195) );
  AOI22D1BWP30P140LVT U11163 ( .A1(i_data_bus[439]), .A2(n10507), .B1(
        i_data_bus[503]), .B2(n10506), .ZN(n7624) );
  AOI22D1BWP30P140LVT U11164 ( .A1(i_data_bus[471]), .A2(n10508), .B1(
        i_data_bus[407]), .B2(n10505), .ZN(n7623) );
  ND2D1BWP30P140LVT U11165 ( .A1(n7624), .A2(n7623), .ZN(N8738) );
  AOI22D1BWP30P140LVT U11166 ( .A1(i_data_bus[457]), .A2(n10508), .B1(
        i_data_bus[425]), .B2(n10507), .ZN(n7626) );
  AOI22D1BWP30P140LVT U11167 ( .A1(i_data_bus[489]), .A2(n10506), .B1(
        i_data_bus[393]), .B2(n10505), .ZN(n7625) );
  ND2D1BWP30P140LVT U11168 ( .A1(n7626), .A2(n7625), .ZN(N8724) );
  AOI22D1BWP30P140LVT U11169 ( .A1(i_data_bus[432]), .A2(n10507), .B1(
        i_data_bus[464]), .B2(n10508), .ZN(n7628) );
  AOI22D1BWP30P140LVT U11170 ( .A1(i_data_bus[496]), .A2(n10506), .B1(
        i_data_bus[400]), .B2(n10505), .ZN(n7627) );
  ND2D1BWP30P140LVT U11171 ( .A1(n7628), .A2(n7627), .ZN(N8731) );
  AOI22D1BWP30P140LVT U11172 ( .A1(i_data_bus[434]), .A2(n10507), .B1(
        i_data_bus[466]), .B2(n10508), .ZN(n7630) );
  AOI22D1BWP30P140LVT U11173 ( .A1(i_data_bus[498]), .A2(n10506), .B1(
        i_data_bus[402]), .B2(n10505), .ZN(n7629) );
  ND2D1BWP30P140LVT U11174 ( .A1(n7630), .A2(n7629), .ZN(N8733) );
  AOI22D1BWP30P140LVT U11175 ( .A1(i_data_bus[493]), .A2(n10506), .B1(
        i_data_bus[461]), .B2(n10508), .ZN(n7632) );
  AOI22D1BWP30P140LVT U11176 ( .A1(i_data_bus[429]), .A2(n10507), .B1(
        i_data_bus[397]), .B2(n10505), .ZN(n7631) );
  ND2D1BWP30P140LVT U11177 ( .A1(n7632), .A2(n7631), .ZN(N8728) );
  AOI22D1BWP30P140LVT U11178 ( .A1(i_data_bus[445]), .A2(n10507), .B1(
        i_data_bus[477]), .B2(n10508), .ZN(n7634) );
  AOI22D1BWP30P140LVT U11179 ( .A1(i_data_bus[509]), .A2(n10506), .B1(
        i_data_bus[413]), .B2(n10505), .ZN(n7633) );
  ND2D1BWP30P140LVT U11180 ( .A1(n7634), .A2(n7633), .ZN(N8744) );
  AOI22D1BWP30P140LVT U11181 ( .A1(i_data_bus[418]), .A2(n10507), .B1(
        i_data_bus[450]), .B2(n10508), .ZN(n7636) );
  AOI22D1BWP30P140LVT U11182 ( .A1(i_data_bus[482]), .A2(n10506), .B1(
        i_data_bus[386]), .B2(n10505), .ZN(n7635) );
  ND2D1BWP30P140LVT U11183 ( .A1(n7636), .A2(n7635), .ZN(N8717) );
  AOI22D1BWP30P140LVT U11184 ( .A1(i_data_bus[458]), .A2(n10508), .B1(
        i_data_bus[426]), .B2(n10507), .ZN(n7638) );
  AOI22D1BWP30P140LVT U11185 ( .A1(i_data_bus[490]), .A2(n10506), .B1(
        i_data_bus[394]), .B2(n10505), .ZN(n7637) );
  ND2D1BWP30P140LVT U11186 ( .A1(n7638), .A2(n7637), .ZN(N8725) );
  AOI22D1BWP30P140LVT U11187 ( .A1(i_data_bus[455]), .A2(n10508), .B1(
        i_data_bus[423]), .B2(n10507), .ZN(n7640) );
  AOI22D1BWP30P140LVT U11188 ( .A1(i_data_bus[487]), .A2(n10506), .B1(
        i_data_bus[391]), .B2(n10505), .ZN(n7639) );
  ND2D1BWP30P140LVT U11189 ( .A1(n7640), .A2(n7639), .ZN(N8722) );
  AOI22D1BWP30P140LVT U11190 ( .A1(i_data_bus[952]), .A2(n10588), .B1(
        i_data_bus[984]), .B2(n10586), .ZN(n7642) );
  AOI22D1BWP30P140LVT U11191 ( .A1(i_data_bus[920]), .A2(n10587), .B1(
        i_data_bus[1016]), .B2(n10585), .ZN(n7641) );
  ND2D1BWP30P140LVT U11192 ( .A1(n7642), .A2(n7641), .ZN(N3981) );
  AOI22D1BWP30P140LVT U11193 ( .A1(i_data_bus[919]), .A2(n10587), .B1(
        i_data_bus[983]), .B2(n10586), .ZN(n7644) );
  AOI22D1BWP30P140LVT U11194 ( .A1(i_data_bus[951]), .A2(n10588), .B1(
        i_data_bus[1015]), .B2(n10585), .ZN(n7643) );
  ND2D1BWP30P140LVT U11195 ( .A1(n7644), .A2(n7643), .ZN(N3980) );
  AOI22D1BWP30P140LVT U11196 ( .A1(i_data_bus[978]), .A2(n10586), .B1(
        i_data_bus[914]), .B2(n10587), .ZN(n7646) );
  AOI22D1BWP30P140LVT U11197 ( .A1(i_data_bus[946]), .A2(n10588), .B1(
        i_data_bus[1010]), .B2(n10585), .ZN(n7645) );
  ND2D1BWP30P140LVT U11198 ( .A1(n7646), .A2(n7645), .ZN(N3975) );
  AOI22D1BWP30P140LVT U11199 ( .A1(i_data_bus[925]), .A2(n10587), .B1(
        i_data_bus[989]), .B2(n10586), .ZN(n7648) );
  AOI22D1BWP30P140LVT U11200 ( .A1(i_data_bus[957]), .A2(n10588), .B1(
        i_data_bus[1021]), .B2(n10585), .ZN(n7647) );
  ND2D1BWP30P140LVT U11201 ( .A1(n7648), .A2(n7647), .ZN(N3986) );
  AOI22D1BWP30P140LVT U11202 ( .A1(i_data_bus[903]), .A2(n10587), .B1(
        i_data_bus[935]), .B2(n10588), .ZN(n7650) );
  AOI22D1BWP30P140LVT U11203 ( .A1(i_data_bus[967]), .A2(n10586), .B1(
        i_data_bus[999]), .B2(n10585), .ZN(n7649) );
  ND2D1BWP30P140LVT U11204 ( .A1(n7650), .A2(n7649), .ZN(N3964) );
  AOI22D1BWP30P140LVT U11205 ( .A1(i_data_bus[924]), .A2(n10587), .B1(
        i_data_bus[956]), .B2(n10588), .ZN(n7652) );
  AOI22D1BWP30P140LVT U11206 ( .A1(i_data_bus[988]), .A2(n10586), .B1(
        i_data_bus[1020]), .B2(n10585), .ZN(n7651) );
  ND2D1BWP30P140LVT U11207 ( .A1(n7652), .A2(n7651), .ZN(N3985) );
  AOI22D1BWP30P140LVT U11208 ( .A1(i_data_bus[940]), .A2(n10588), .B1(
        i_data_bus[972]), .B2(n10586), .ZN(n7654) );
  AOI22D1BWP30P140LVT U11209 ( .A1(i_data_bus[908]), .A2(n10587), .B1(
        i_data_bus[1004]), .B2(n10585), .ZN(n7653) );
  ND2D1BWP30P140LVT U11210 ( .A1(n7654), .A2(n7653), .ZN(N3969) );
  AOI22D1BWP30P140LVT U11211 ( .A1(i_data_bus[961]), .A2(n10586), .B1(
        i_data_bus[897]), .B2(n10587), .ZN(n7656) );
  AOI22D1BWP30P140LVT U11212 ( .A1(i_data_bus[929]), .A2(n10588), .B1(
        i_data_bus[993]), .B2(n10585), .ZN(n7655) );
  ND2D1BWP30P140LVT U11213 ( .A1(n7656), .A2(n7655), .ZN(N3958) );
  AOI22D1BWP30P140LVT U11214 ( .A1(i_data_bus[923]), .A2(n10587), .B1(
        i_data_bus[987]), .B2(n10586), .ZN(n7658) );
  AOI22D1BWP30P140LVT U11215 ( .A1(i_data_bus[955]), .A2(n10588), .B1(
        i_data_bus[1019]), .B2(n10585), .ZN(n7657) );
  ND2D1BWP30P140LVT U11216 ( .A1(n7658), .A2(n7657), .ZN(N3984) );
  AOI22D1BWP30P140LVT U11217 ( .A1(i_data_bus[550]), .A2(n10598), .B1(
        i_data_bus[518]), .B2(n10597), .ZN(n7660) );
  AOI22D1BWP30P140LVT U11218 ( .A1(i_data_bus[614]), .A2(n10599), .B1(
        i_data_bus[582]), .B2(n10600), .ZN(n7659) );
  ND2D1BWP30P140LVT U11219 ( .A1(n7660), .A2(n7659), .ZN(N3315) );
  AOI22D1BWP30P140LVT U11220 ( .A1(i_data_bus[512]), .A2(n10597), .B1(
        i_data_bus[544]), .B2(n10598), .ZN(n7662) );
  AOI22D1BWP30P140LVT U11221 ( .A1(i_data_bus[608]), .A2(n10599), .B1(
        i_data_bus[576]), .B2(n10600), .ZN(n7661) );
  ND2D1BWP30P140LVT U11222 ( .A1(n7662), .A2(n7661), .ZN(N3309) );
  AOI22D1BWP30P140LVT U11223 ( .A1(i_data_bus[615]), .A2(n10599), .B1(
        i_data_bus[551]), .B2(n10598), .ZN(n7664) );
  AOI22D1BWP30P140LVT U11224 ( .A1(i_data_bus[519]), .A2(n10597), .B1(
        i_data_bus[583]), .B2(n10600), .ZN(n7663) );
  ND2D1BWP30P140LVT U11225 ( .A1(n7664), .A2(n7663), .ZN(N3316) );
  AOI22D1BWP30P140LVT U11226 ( .A1(i_data_bus[638]), .A2(n10599), .B1(
        i_data_bus[542]), .B2(n10597), .ZN(n7666) );
  AOI22D1BWP30P140LVT U11227 ( .A1(i_data_bus[574]), .A2(n10598), .B1(
        i_data_bus[606]), .B2(n10600), .ZN(n7665) );
  ND2D1BWP30P140LVT U11228 ( .A1(n7666), .A2(n7665), .ZN(N3339) );
  AOI22D1BWP30P140LVT U11229 ( .A1(i_data_bus[609]), .A2(n10599), .B1(
        i_data_bus[545]), .B2(n10598), .ZN(n7668) );
  AOI22D1BWP30P140LVT U11230 ( .A1(i_data_bus[513]), .A2(n10597), .B1(
        i_data_bus[577]), .B2(n10600), .ZN(n7667) );
  ND2D1BWP30P140LVT U11231 ( .A1(n7668), .A2(n7667), .ZN(N3310) );
  AOI22D1BWP30P140LVT U11232 ( .A1(i_data_bus[648]), .A2(n10563), .B1(
        i_data_bus[712]), .B2(n10561), .ZN(n7670) );
  AOI22D1BWP30P140LVT U11233 ( .A1(i_data_bus[744]), .A2(n10562), .B1(
        i_data_bus[680]), .B2(n10564), .ZN(n7669) );
  ND2D1BWP30P140LVT U11234 ( .A1(n7670), .A2(n7669), .ZN(N5407) );
  AOI22D1BWP30P140LVT U11235 ( .A1(i_data_bus[715]), .A2(n10561), .B1(
        i_data_bus[747]), .B2(n10562), .ZN(n7672) );
  AOI22D1BWP30P140LVT U11236 ( .A1(i_data_bus[651]), .A2(n10563), .B1(
        i_data_bus[683]), .B2(n10564), .ZN(n7671) );
  ND2D1BWP30P140LVT U11237 ( .A1(n7672), .A2(n7671), .ZN(N5410) );
  AOI22D1BWP30P140LVT U11238 ( .A1(i_data_bus[657]), .A2(n10563), .B1(
        i_data_bus[721]), .B2(n10561), .ZN(n7674) );
  AOI22D1BWP30P140LVT U11239 ( .A1(i_data_bus[753]), .A2(n10562), .B1(
        i_data_bus[689]), .B2(n10564), .ZN(n7673) );
  ND2D1BWP30P140LVT U11240 ( .A1(n7674), .A2(n7673), .ZN(N5416) );
  AOI22D1BWP30P140LVT U11241 ( .A1(i_data_bus[764]), .A2(n10562), .B1(
        i_data_bus[668]), .B2(n10563), .ZN(n7676) );
  AOI22D1BWP30P140LVT U11242 ( .A1(i_data_bus[732]), .A2(n10561), .B1(
        i_data_bus[700]), .B2(n10564), .ZN(n7675) );
  ND2D1BWP30P140LVT U11243 ( .A1(n7676), .A2(n7675), .ZN(N5427) );
  AOI22D1BWP30P140LVT U11244 ( .A1(i_data_bus[734]), .A2(n10561), .B1(
        i_data_bus[670]), .B2(n10563), .ZN(n7678) );
  AOI22D1BWP30P140LVT U11245 ( .A1(i_data_bus[766]), .A2(n10562), .B1(
        i_data_bus[702]), .B2(n10564), .ZN(n7677) );
  ND2D1BWP30P140LVT U11246 ( .A1(n7678), .A2(n7677), .ZN(N5429) );
  AOI22D1BWP30P140LVT U11247 ( .A1(i_data_bus[710]), .A2(n10561), .B1(
        i_data_bus[742]), .B2(n10562), .ZN(n7680) );
  AOI22D1BWP30P140LVT U11248 ( .A1(i_data_bus[646]), .A2(n10563), .B1(
        i_data_bus[678]), .B2(n10564), .ZN(n7679) );
  ND2D1BWP30P140LVT U11249 ( .A1(n7680), .A2(n7679), .ZN(N5405) );
  AOI22D1BWP30P140LVT U11250 ( .A1(i_data_bus[733]), .A2(n10561), .B1(
        i_data_bus[765]), .B2(n10562), .ZN(n7682) );
  AOI22D1BWP30P140LVT U11251 ( .A1(i_data_bus[669]), .A2(n10563), .B1(
        i_data_bus[701]), .B2(n10564), .ZN(n7681) );
  ND2D1BWP30P140LVT U11252 ( .A1(n7682), .A2(n7681), .ZN(N5428) );
  AOI22D1BWP30P140LVT U11253 ( .A1(i_data_bus[604]), .A2(n10437), .B1(
        i_data_bus[572]), .B2(n10439), .ZN(n7684) );
  AOI22D1BWP30P140LVT U11254 ( .A1(i_data_bus[636]), .A2(n10440), .B1(
        i_data_bus[540]), .B2(n10438), .ZN(n7683) );
  ND2D1BWP30P140LVT U11255 ( .A1(n7684), .A2(n7683), .ZN(N12707) );
  AOI22D1BWP30P140LVT U11256 ( .A1(i_data_bus[557]), .A2(n10439), .B1(
        i_data_bus[589]), .B2(n10437), .ZN(n7686) );
  AOI22D1BWP30P140LVT U11257 ( .A1(i_data_bus[621]), .A2(n10440), .B1(
        i_data_bus[525]), .B2(n10438), .ZN(n7685) );
  ND2D1BWP30P140LVT U11258 ( .A1(n7686), .A2(n7685), .ZN(N12692) );
  AOI22D1BWP30P140LVT U11259 ( .A1(i_data_bus[579]), .A2(n10437), .B1(
        i_data_bus[547]), .B2(n10439), .ZN(n7688) );
  AOI22D1BWP30P140LVT U11260 ( .A1(i_data_bus[611]), .A2(n10440), .B1(
        i_data_bus[515]), .B2(n10438), .ZN(n7687) );
  ND2D1BWP30P140LVT U11261 ( .A1(n7688), .A2(n7687), .ZN(N12682) );
  AOI22D1BWP30P140LVT U11262 ( .A1(i_data_bus[550]), .A2(n10439), .B1(
        i_data_bus[582]), .B2(n10437), .ZN(n7690) );
  AOI22D1BWP30P140LVT U11263 ( .A1(i_data_bus[614]), .A2(n10440), .B1(
        i_data_bus[518]), .B2(n10438), .ZN(n7689) );
  ND2D1BWP30P140LVT U11264 ( .A1(n7690), .A2(n7689), .ZN(N12685) );
  AOI22D1BWP30P140LVT U11265 ( .A1(i_data_bus[552]), .A2(n10439), .B1(
        i_data_bus[584]), .B2(n10437), .ZN(n7692) );
  AOI22D1BWP30P140LVT U11266 ( .A1(i_data_bus[616]), .A2(n10440), .B1(
        i_data_bus[520]), .B2(n10438), .ZN(n7691) );
  ND2D1BWP30P140LVT U11267 ( .A1(n7692), .A2(n7691), .ZN(N12687) );
  AOI22D1BWP30P140LVT U11268 ( .A1(i_data_bus[805]), .A2(n10560), .B1(
        i_data_bus[773]), .B2(n10558), .ZN(n7694) );
  AOI22D1BWP30P140LVT U11269 ( .A1(i_data_bus[869]), .A2(n10559), .B1(
        i_data_bus[837]), .B2(n10557), .ZN(n7693) );
  ND2D1BWP30P140LVT U11270 ( .A1(n7694), .A2(n7693), .ZN(N5620) );
  AOI22D1BWP30P140LVT U11271 ( .A1(i_data_bus[827]), .A2(n10560), .B1(
        i_data_bus[891]), .B2(n10559), .ZN(n7696) );
  AOI22D1BWP30P140LVT U11272 ( .A1(i_data_bus[795]), .A2(n10558), .B1(
        i_data_bus[859]), .B2(n10557), .ZN(n7695) );
  ND2D1BWP30P140LVT U11273 ( .A1(n7696), .A2(n7695), .ZN(N5642) );
  AOI22D1BWP30P140LVT U11274 ( .A1(i_data_bus[883]), .A2(n10559), .B1(
        i_data_bus[787]), .B2(n10558), .ZN(n7698) );
  AOI22D1BWP30P140LVT U11275 ( .A1(i_data_bus[819]), .A2(n10560), .B1(
        i_data_bus[851]), .B2(n10557), .ZN(n7697) );
  ND2D1BWP30P140LVT U11276 ( .A1(n7698), .A2(n7697), .ZN(N5634) );
  AOI22D1BWP30P140LVT U11277 ( .A1(i_data_bus[878]), .A2(n10559), .B1(
        i_data_bus[782]), .B2(n10558), .ZN(n7700) );
  AOI22D1BWP30P140LVT U11278 ( .A1(i_data_bus[814]), .A2(n10560), .B1(
        i_data_bus[846]), .B2(n10557), .ZN(n7699) );
  ND2D1BWP30P140LVT U11279 ( .A1(n7700), .A2(n7699), .ZN(N5629) );
  AOI22D1BWP30P140LVT U11280 ( .A1(i_data_bus[886]), .A2(n10559), .B1(
        i_data_bus[790]), .B2(n10558), .ZN(n7702) );
  AOI22D1BWP30P140LVT U11281 ( .A1(i_data_bus[822]), .A2(n10560), .B1(
        i_data_bus[854]), .B2(n10557), .ZN(n7701) );
  ND2D1BWP30P140LVT U11282 ( .A1(n7702), .A2(n7701), .ZN(N5637) );
  AOI22D1BWP30P140LVT U11283 ( .A1(i_data_bus[801]), .A2(n10560), .B1(
        i_data_bus[769]), .B2(n10558), .ZN(n7704) );
  AOI22D1BWP30P140LVT U11284 ( .A1(i_data_bus[865]), .A2(n10559), .B1(
        i_data_bus[833]), .B2(n10557), .ZN(n7703) );
  ND2D1BWP30P140LVT U11285 ( .A1(n7704), .A2(n7703), .ZN(N5616) );
  AOI22D1BWP30P140LVT U11286 ( .A1(i_data_bus[885]), .A2(n10559), .B1(
        i_data_bus[821]), .B2(n10560), .ZN(n7706) );
  AOI22D1BWP30P140LVT U11287 ( .A1(i_data_bus[789]), .A2(n10558), .B1(
        i_data_bus[853]), .B2(n10557), .ZN(n7705) );
  ND2D1BWP30P140LVT U11288 ( .A1(n7706), .A2(n7705), .ZN(N5636) );
  AOI22D1BWP30P140LVT U11289 ( .A1(i_data_bus[90]), .A2(n10517), .B1(
        i_data_bus[26]), .B2(n10520), .ZN(n7708) );
  AOI22D1BWP30P140LVT U11290 ( .A1(i_data_bus[122]), .A2(n10519), .B1(
        i_data_bus[58]), .B2(n10518), .ZN(n7707) );
  ND2D1BWP30P140LVT U11291 ( .A1(n7708), .A2(n7707), .ZN(N8093) );
  AOI22D1BWP30P140LVT U11292 ( .A1(i_data_bus[126]), .A2(n10519), .B1(
        i_data_bus[30]), .B2(n10520), .ZN(n7710) );
  AOI22D1BWP30P140LVT U11293 ( .A1(i_data_bus[94]), .A2(n10517), .B1(
        i_data_bus[62]), .B2(n10518), .ZN(n7709) );
  ND2D1BWP30P140LVT U11294 ( .A1(n7710), .A2(n7709), .ZN(N8097) );
  AOI22D1BWP30P140LVT U11295 ( .A1(i_data_bus[98]), .A2(n10519), .B1(
        i_data_bus[2]), .B2(n10520), .ZN(n7712) );
  AOI22D1BWP30P140LVT U11296 ( .A1(i_data_bus[66]), .A2(n10517), .B1(
        i_data_bus[34]), .B2(n10518), .ZN(n7711) );
  ND2D1BWP30P140LVT U11297 ( .A1(n7712), .A2(n7711), .ZN(N8069) );
  AOI22D1BWP30P140LVT U11298 ( .A1(i_data_bus[95]), .A2(n10517), .B1(
        i_data_bus[31]), .B2(n10520), .ZN(n7714) );
  AOI22D1BWP30P140LVT U11299 ( .A1(i_data_bus[127]), .A2(n10519), .B1(
        i_data_bus[63]), .B2(n10518), .ZN(n7713) );
  ND2D1BWP30P140LVT U11300 ( .A1(n7714), .A2(n7713), .ZN(N8098) );
  AOI22D1BWP30P140LVT U11301 ( .A1(i_data_bus[108]), .A2(n10519), .B1(
        i_data_bus[12]), .B2(n10520), .ZN(n7716) );
  AOI22D1BWP30P140LVT U11302 ( .A1(i_data_bus[76]), .A2(n10517), .B1(
        i_data_bus[44]), .B2(n10518), .ZN(n7715) );
  ND2D1BWP30P140LVT U11303 ( .A1(n7716), .A2(n7715), .ZN(N8079) );
  AOI22D1BWP30P140LVT U11304 ( .A1(i_data_bus[8]), .A2(n10520), .B1(
        i_data_bus[104]), .B2(n10519), .ZN(n7718) );
  AOI22D1BWP30P140LVT U11305 ( .A1(i_data_bus[40]), .A2(n10518), .B1(
        i_data_bus[72]), .B2(n10517), .ZN(n7717) );
  ND2D1BWP30P140LVT U11306 ( .A1(n7718), .A2(n7717), .ZN(N8075) );
  AOI22D1BWP30P140LVT U11307 ( .A1(i_data_bus[996]), .A2(n10457), .B1(
        i_data_bus[964]), .B2(n10459), .ZN(n7720) );
  AOI22D1BWP30P140LVT U11308 ( .A1(i_data_bus[932]), .A2(n10460), .B1(
        i_data_bus[900]), .B2(n10458), .ZN(n7719) );
  ND2D1BWP30P140LVT U11309 ( .A1(n7720), .A2(n7719), .ZN(N11457) );
  AOI22D1BWP30P140LVT U11310 ( .A1(i_data_bus[1007]), .A2(n10457), .B1(
        i_data_bus[975]), .B2(n10459), .ZN(n7722) );
  AOI22D1BWP30P140LVT U11311 ( .A1(i_data_bus[943]), .A2(n10460), .B1(
        i_data_bus[911]), .B2(n10458), .ZN(n7721) );
  ND2D1BWP30P140LVT U11312 ( .A1(n7722), .A2(n7721), .ZN(N11468) );
  AOI22D1BWP30P140LVT U11313 ( .A1(i_data_bus[939]), .A2(n10460), .B1(
        i_data_bus[971]), .B2(n10459), .ZN(n7724) );
  AOI22D1BWP30P140LVT U11314 ( .A1(i_data_bus[1003]), .A2(n10457), .B1(
        i_data_bus[907]), .B2(n10458), .ZN(n7723) );
  ND2D1BWP30P140LVT U11315 ( .A1(n7724), .A2(n7723), .ZN(N11464) );
  AOI22D1BWP30P140LVT U11316 ( .A1(i_data_bus[6]), .A2(n10520), .B1(
        i_data_bus[102]), .B2(n10519), .ZN(n7726) );
  AOI22D1BWP30P140LVT U11317 ( .A1(i_data_bus[38]), .A2(n10518), .B1(
        i_data_bus[70]), .B2(n10517), .ZN(n7725) );
  ND2D1BWP30P140LVT U11318 ( .A1(n7726), .A2(n7725), .ZN(N8073) );
  AOI22D1BWP30P140LVT U11319 ( .A1(i_data_bus[100]), .A2(n10519), .B1(
        i_data_bus[36]), .B2(n10518), .ZN(n7728) );
  AOI22D1BWP30P140LVT U11320 ( .A1(i_data_bus[4]), .A2(n10520), .B1(
        i_data_bus[68]), .B2(n10517), .ZN(n7727) );
  ND2D1BWP30P140LVT U11321 ( .A1(n7728), .A2(n7727), .ZN(N8071) );
  AOI22D1BWP30P140LVT U11322 ( .A1(i_data_bus[116]), .A2(n10519), .B1(
        i_data_bus[20]), .B2(n10520), .ZN(n7730) );
  AOI22D1BWP30P140LVT U11323 ( .A1(i_data_bus[52]), .A2(n10518), .B1(
        i_data_bus[84]), .B2(n10517), .ZN(n7729) );
  ND2D1BWP30P140LVT U11324 ( .A1(n7730), .A2(n7729), .ZN(N8087) );
  AOI22D1BWP30P140LVT U11325 ( .A1(i_data_bus[600]), .A2(n10600), .B1(
        i_data_bus[632]), .B2(n10599), .ZN(n7732) );
  AOI22D1BWP30P140LVT U11326 ( .A1(i_data_bus[536]), .A2(n10597), .B1(
        i_data_bus[568]), .B2(n10598), .ZN(n7731) );
  ND2D1BWP30P140LVT U11327 ( .A1(n7732), .A2(n7731), .ZN(N3333) );
  AOI22D1BWP30P140LVT U11328 ( .A1(i_data_bus[531]), .A2(n10597), .B1(
        i_data_bus[627]), .B2(n10599), .ZN(n7734) );
  AOI22D1BWP30P140LVT U11329 ( .A1(i_data_bus[595]), .A2(n10600), .B1(
        i_data_bus[563]), .B2(n10598), .ZN(n7733) );
  ND2D1BWP30P140LVT U11330 ( .A1(n7734), .A2(n7733), .ZN(N3328) );
  AOI22D1BWP30P140LVT U11331 ( .A1(i_data_bus[951]), .A2(n10460), .B1(
        i_data_bus[983]), .B2(n10459), .ZN(n7736) );
  AOI22D1BWP30P140LVT U11332 ( .A1(i_data_bus[919]), .A2(n10458), .B1(
        i_data_bus[1015]), .B2(n10457), .ZN(n7735) );
  ND2D1BWP30P140LVT U11333 ( .A1(n7736), .A2(n7735), .ZN(N11476) );
  AOI22D1BWP30P140LVT U11334 ( .A1(i_data_bus[920]), .A2(n10458), .B1(
        i_data_bus[984]), .B2(n10459), .ZN(n7738) );
  AOI22D1BWP30P140LVT U11335 ( .A1(i_data_bus[952]), .A2(n10460), .B1(
        i_data_bus[1016]), .B2(n10457), .ZN(n7737) );
  ND2D1BWP30P140LVT U11336 ( .A1(n7738), .A2(n7737), .ZN(N11477) );
  AOI22D1BWP30P140LVT U11337 ( .A1(i_data_bus[604]), .A2(n10469), .B1(
        i_data_bus[572]), .B2(n10472), .ZN(n7740) );
  AOI22D1BWP30P140LVT U11338 ( .A1(i_data_bus[636]), .A2(n10470), .B1(
        i_data_bus[540]), .B2(n10471), .ZN(n7739) );
  ND2D1BWP30P140LVT U11339 ( .A1(n7740), .A2(n7739), .ZN(N10833) );
  AOI22D1BWP30P140LVT U11340 ( .A1(i_data_bus[1004]), .A2(n10457), .B1(
        i_data_bus[972]), .B2(n10459), .ZN(n7742) );
  AOI22D1BWP30P140LVT U11341 ( .A1(i_data_bus[908]), .A2(n10458), .B1(
        i_data_bus[940]), .B2(n10460), .ZN(n7741) );
  ND2D1BWP30P140LVT U11342 ( .A1(n7742), .A2(n7741), .ZN(N11465) );
  AOI22D1BWP30P140LVT U11343 ( .A1(i_data_bus[898]), .A2(n10458), .B1(
        i_data_bus[962]), .B2(n10459), .ZN(n7744) );
  AOI22D1BWP30P140LVT U11344 ( .A1(i_data_bus[994]), .A2(n10457), .B1(
        i_data_bus[930]), .B2(n10460), .ZN(n7743) );
  ND2D1BWP30P140LVT U11345 ( .A1(n7744), .A2(n7743), .ZN(N11455) );
  AOI22D1BWP30P140LVT U11346 ( .A1(i_data_bus[616]), .A2(n10470), .B1(
        i_data_bus[584]), .B2(n10469), .ZN(n7746) );
  AOI22D1BWP30P140LVT U11347 ( .A1(i_data_bus[552]), .A2(n10472), .B1(
        i_data_bus[520]), .B2(n10471), .ZN(n7745) );
  ND2D1BWP30P140LVT U11348 ( .A1(n7746), .A2(n7745), .ZN(N10813) );
  AOI22D1BWP30P140LVT U11349 ( .A1(i_data_bus[913]), .A2(n10458), .B1(
        i_data_bus[977]), .B2(n10459), .ZN(n7748) );
  AOI22D1BWP30P140LVT U11350 ( .A1(i_data_bus[1009]), .A2(n10457), .B1(
        i_data_bus[945]), .B2(n10460), .ZN(n7747) );
  ND2D1BWP30P140LVT U11351 ( .A1(n7748), .A2(n7747), .ZN(N11470) );
  AOI22D1BWP30P140LVT U11352 ( .A1(i_data_bus[557]), .A2(n10472), .B1(
        i_data_bus[589]), .B2(n10469), .ZN(n7750) );
  AOI22D1BWP30P140LVT U11353 ( .A1(i_data_bus[621]), .A2(n10470), .B1(
        i_data_bus[525]), .B2(n10471), .ZN(n7749) );
  ND2D1BWP30P140LVT U11354 ( .A1(n7750), .A2(n7749), .ZN(N10818) );
  AOI22D1BWP30P140LVT U11355 ( .A1(i_data_bus[1023]), .A2(n10457), .B1(
        i_data_bus[991]), .B2(n10459), .ZN(n7752) );
  AOI22D1BWP30P140LVT U11356 ( .A1(i_data_bus[927]), .A2(n10458), .B1(
        i_data_bus[959]), .B2(n10460), .ZN(n7751) );
  ND2D1BWP30P140LVT U11357 ( .A1(n7752), .A2(n7751), .ZN(N11484) );
  AOI22D1BWP30P140LVT U11358 ( .A1(i_data_bus[560]), .A2(n10472), .B1(
        i_data_bus[592]), .B2(n10469), .ZN(n7754) );
  AOI22D1BWP30P140LVT U11359 ( .A1(i_data_bus[624]), .A2(n10470), .B1(
        i_data_bus[528]), .B2(n10471), .ZN(n7753) );
  ND2D1BWP30P140LVT U11360 ( .A1(n7754), .A2(n7753), .ZN(N10821) );
  AOI22D1BWP30P140LVT U11361 ( .A1(i_data_bus[568]), .A2(n10472), .B1(
        i_data_bus[632]), .B2(n10470), .ZN(n7756) );
  AOI22D1BWP30P140LVT U11362 ( .A1(i_data_bus[600]), .A2(n10469), .B1(
        i_data_bus[536]), .B2(n10471), .ZN(n7755) );
  ND2D1BWP30P140LVT U11363 ( .A1(n7756), .A2(n7755), .ZN(N10829) );
  AOI22D1BWP30P140LVT U11364 ( .A1(i_data_bus[601]), .A2(n10469), .B1(
        i_data_bus[633]), .B2(n10470), .ZN(n7758) );
  AOI22D1BWP30P140LVT U11365 ( .A1(i_data_bus[569]), .A2(n10472), .B1(
        i_data_bus[537]), .B2(n10471), .ZN(n7757) );
  ND2D1BWP30P140LVT U11366 ( .A1(n7758), .A2(n7757), .ZN(N10830) );
  AOI22D1BWP30P140LVT U11367 ( .A1(i_data_bus[574]), .A2(n10472), .B1(
        i_data_bus[606]), .B2(n10469), .ZN(n7760) );
  AOI22D1BWP30P140LVT U11368 ( .A1(i_data_bus[638]), .A2(n10470), .B1(
        i_data_bus[542]), .B2(n10471), .ZN(n7759) );
  ND2D1BWP30P140LVT U11369 ( .A1(n7760), .A2(n7759), .ZN(N10835) );
  AOI22D1BWP30P140LVT U11370 ( .A1(i_data_bus[586]), .A2(n10600), .B1(
        i_data_bus[618]), .B2(n10599), .ZN(n7762) );
  AOI22D1BWP30P140LVT U11371 ( .A1(i_data_bus[554]), .A2(n10598), .B1(
        i_data_bus[522]), .B2(n10597), .ZN(n7761) );
  ND2D1BWP30P140LVT U11372 ( .A1(n7762), .A2(n7761), .ZN(N3319) );
  AOI22D1BWP30P140LVT U11373 ( .A1(i_data_bus[566]), .A2(n10598), .B1(
        i_data_bus[630]), .B2(n10599), .ZN(n7764) );
  AOI22D1BWP30P140LVT U11374 ( .A1(i_data_bus[598]), .A2(n10600), .B1(
        i_data_bus[534]), .B2(n10597), .ZN(n7763) );
  ND2D1BWP30P140LVT U11375 ( .A1(n7764), .A2(n7763), .ZN(N3331) );
  AOI22D1BWP30P140LVT U11376 ( .A1(i_data_bus[557]), .A2(n10598), .B1(
        i_data_bus[621]), .B2(n10599), .ZN(n7766) );
  AOI22D1BWP30P140LVT U11377 ( .A1(i_data_bus[525]), .A2(n10597), .B1(
        i_data_bus[589]), .B2(n10600), .ZN(n7765) );
  ND2D1BWP30P140LVT U11378 ( .A1(n7766), .A2(n7765), .ZN(N3322) );
  AOI22D1BWP30P140LVT U11379 ( .A1(i_data_bus[602]), .A2(n10600), .B1(
        i_data_bus[634]), .B2(n10599), .ZN(n7768) );
  AOI22D1BWP30P140LVT U11380 ( .A1(i_data_bus[570]), .A2(n10598), .B1(
        i_data_bus[538]), .B2(n10597), .ZN(n7767) );
  ND2D1BWP30P140LVT U11381 ( .A1(n7768), .A2(n7767), .ZN(N3335) );
  AOI22D1BWP30P140LVT U11382 ( .A1(i_data_bus[556]), .A2(n10598), .B1(
        i_data_bus[620]), .B2(n10599), .ZN(n7770) );
  AOI22D1BWP30P140LVT U11383 ( .A1(i_data_bus[524]), .A2(n10597), .B1(
        i_data_bus[588]), .B2(n10600), .ZN(n7769) );
  ND2D1BWP30P140LVT U11384 ( .A1(n7770), .A2(n7769), .ZN(N3321) );
  AOI22D1BWP30P140LVT U11385 ( .A1(i_data_bus[526]), .A2(n10597), .B1(
        i_data_bus[622]), .B2(n10599), .ZN(n7772) );
  AOI22D1BWP30P140LVT U11386 ( .A1(i_data_bus[558]), .A2(n10598), .B1(
        i_data_bus[590]), .B2(n10600), .ZN(n7771) );
  ND2D1BWP30P140LVT U11387 ( .A1(n7772), .A2(n7771), .ZN(N3323) );
  AOI22D1BWP30P140LVT U11388 ( .A1(i_data_bus[593]), .A2(n10600), .B1(
        i_data_bus[625]), .B2(n10599), .ZN(n7774) );
  AOI22D1BWP30P140LVT U11389 ( .A1(i_data_bus[561]), .A2(n10598), .B1(
        i_data_bus[529]), .B2(n10597), .ZN(n7773) );
  ND2D1BWP30P140LVT U11390 ( .A1(n7774), .A2(n7773), .ZN(N3326) );
  AOI22D1BWP30P140LVT U11391 ( .A1(i_data_bus[761]), .A2(n10403), .B1(
        i_data_bus[697]), .B2(n10404), .ZN(n7776) );
  AOI22D1BWP30P140LVT U11392 ( .A1(i_data_bus[665]), .A2(n10401), .B1(
        i_data_bus[729]), .B2(n10402), .ZN(n7775) );
  ND2D1BWP30P140LVT U11393 ( .A1(n7776), .A2(n7775), .ZN(N14794) );
  AOI22D1BWP30P140LVT U11394 ( .A1(i_data_bus[753]), .A2(n10403), .B1(
        i_data_bus[689]), .B2(n10404), .ZN(n7778) );
  AOI22D1BWP30P140LVT U11395 ( .A1(i_data_bus[657]), .A2(n10401), .B1(
        i_data_bus[721]), .B2(n10402), .ZN(n7777) );
  ND2D1BWP30P140LVT U11396 ( .A1(n7778), .A2(n7777), .ZN(N14786) );
  AOI22D1BWP30P140LVT U11397 ( .A1(i_data_bus[695]), .A2(n10404), .B1(
        i_data_bus[759]), .B2(n10403), .ZN(n7780) );
  AOI22D1BWP30P140LVT U11398 ( .A1(i_data_bus[663]), .A2(n10401), .B1(
        i_data_bus[727]), .B2(n10402), .ZN(n7779) );
  ND2D1BWP30P140LVT U11399 ( .A1(n7780), .A2(n7779), .ZN(N14792) );
  AOI22D1BWP30P140LVT U11400 ( .A1(i_data_bus[755]), .A2(n10403), .B1(
        i_data_bus[691]), .B2(n10404), .ZN(n7782) );
  AOI22D1BWP30P140LVT U11401 ( .A1(i_data_bus[659]), .A2(n10401), .B1(
        i_data_bus[723]), .B2(n10402), .ZN(n7781) );
  ND2D1BWP30P140LVT U11402 ( .A1(n7782), .A2(n7781), .ZN(N14788) );
  AOI22D1BWP30P140LVT U11403 ( .A1(i_data_bus[675]), .A2(n10404), .B1(
        i_data_bus[739]), .B2(n10403), .ZN(n7784) );
  AOI22D1BWP30P140LVT U11404 ( .A1(i_data_bus[643]), .A2(n10401), .B1(
        i_data_bus[707]), .B2(n10402), .ZN(n7783) );
  ND2D1BWP30P140LVT U11405 ( .A1(n7784), .A2(n7783), .ZN(N14772) );
  AOI22D1BWP30P140LVT U11406 ( .A1(i_data_bus[767]), .A2(n10403), .B1(
        i_data_bus[671]), .B2(n10401), .ZN(n7786) );
  AOI22D1BWP30P140LVT U11407 ( .A1(i_data_bus[703]), .A2(n10404), .B1(
        i_data_bus[735]), .B2(n10402), .ZN(n7785) );
  ND2D1BWP30P140LVT U11408 ( .A1(n7786), .A2(n7785), .ZN(N14800) );
  AOI22D1BWP30P140LVT U11409 ( .A1(i_data_bus[667]), .A2(n10401), .B1(
        i_data_bus[699]), .B2(n10404), .ZN(n7788) );
  AOI22D1BWP30P140LVT U11410 ( .A1(i_data_bus[763]), .A2(n10403), .B1(
        i_data_bus[731]), .B2(n10402), .ZN(n7787) );
  ND2D1BWP30P140LVT U11411 ( .A1(n7788), .A2(n7787), .ZN(N14796) );
  AOI22D1BWP30P140LVT U11412 ( .A1(i_data_bus[692]), .A2(n10404), .B1(
        i_data_bus[660]), .B2(n10401), .ZN(n7790) );
  AOI22D1BWP30P140LVT U11413 ( .A1(i_data_bus[756]), .A2(n10403), .B1(
        i_data_bus[724]), .B2(n10402), .ZN(n7789) );
  ND2D1BWP30P140LVT U11414 ( .A1(n7790), .A2(n7789), .ZN(N14789) );
  AOI22D1BWP30P140LVT U11415 ( .A1(i_data_bus[236]), .A2(n10418), .B1(
        i_data_bus[140]), .B2(n10417), .ZN(n7792) );
  AOI22D1BWP30P140LVT U11416 ( .A1(i_data_bus[204]), .A2(n10419), .B1(
        i_data_bus[172]), .B2(n10420), .ZN(n7791) );
  ND2D1BWP30P140LVT U11417 ( .A1(n7792), .A2(n7791), .ZN(N13917) );
  AOI22D1BWP30P140LVT U11418 ( .A1(i_data_bus[195]), .A2(n10419), .B1(
        i_data_bus[131]), .B2(n10417), .ZN(n7794) );
  AOI22D1BWP30P140LVT U11419 ( .A1(i_data_bus[227]), .A2(n10418), .B1(
        i_data_bus[163]), .B2(n10420), .ZN(n7793) );
  ND2D1BWP30P140LVT U11420 ( .A1(n7794), .A2(n7793), .ZN(N13908) );
  AOI22D1BWP30P140LVT U11421 ( .A1(i_data_bus[248]), .A2(n10418), .B1(
        i_data_bus[152]), .B2(n10417), .ZN(n7796) );
  AOI22D1BWP30P140LVT U11422 ( .A1(i_data_bus[216]), .A2(n10419), .B1(
        i_data_bus[184]), .B2(n10420), .ZN(n7795) );
  ND2D1BWP30P140LVT U11423 ( .A1(n7796), .A2(n7795), .ZN(N13929) );
  AOI22D1BWP30P140LVT U11424 ( .A1(i_data_bus[143]), .A2(n10417), .B1(
        i_data_bus[239]), .B2(n10418), .ZN(n7798) );
  AOI22D1BWP30P140LVT U11425 ( .A1(i_data_bus[207]), .A2(n10419), .B1(
        i_data_bus[175]), .B2(n10420), .ZN(n7797) );
  ND2D1BWP30P140LVT U11426 ( .A1(n7798), .A2(n7797), .ZN(N13920) );
  AOI22D1BWP30P140LVT U11427 ( .A1(i_data_bus[201]), .A2(n10419), .B1(
        i_data_bus[137]), .B2(n10417), .ZN(n7800) );
  AOI22D1BWP30P140LVT U11428 ( .A1(i_data_bus[233]), .A2(n10418), .B1(
        i_data_bus[169]), .B2(n10420), .ZN(n7799) );
  ND2D1BWP30P140LVT U11429 ( .A1(n7800), .A2(n7799), .ZN(N13914) );
  AOI22D1BWP30P140LVT U11430 ( .A1(i_data_bus[230]), .A2(n10418), .B1(
        i_data_bus[134]), .B2(n10417), .ZN(n7802) );
  AOI22D1BWP30P140LVT U11431 ( .A1(i_data_bus[198]), .A2(n10419), .B1(
        i_data_bus[166]), .B2(n10420), .ZN(n7801) );
  ND2D1BWP30P140LVT U11432 ( .A1(n7802), .A2(n7801), .ZN(N13911) );
  AOI22D1BWP30P140LVT U11433 ( .A1(i_data_bus[150]), .A2(n10417), .B1(
        i_data_bus[246]), .B2(n10418), .ZN(n7804) );
  AOI22D1BWP30P140LVT U11434 ( .A1(i_data_bus[214]), .A2(n10419), .B1(
        i_data_bus[182]), .B2(n10420), .ZN(n7803) );
  ND2D1BWP30P140LVT U11435 ( .A1(n7804), .A2(n7803), .ZN(N13927) );
  AOI22D1BWP30P140LVT U11436 ( .A1(i_data_bus[229]), .A2(n10418), .B1(
        i_data_bus[197]), .B2(n10419), .ZN(n7806) );
  AOI22D1BWP30P140LVT U11437 ( .A1(i_data_bus[133]), .A2(n10417), .B1(
        i_data_bus[165]), .B2(n10420), .ZN(n7805) );
  ND2D1BWP30P140LVT U11438 ( .A1(n7806), .A2(n7805), .ZN(N13910) );
  AOI22D1BWP30P140LVT U11439 ( .A1(i_data_bus[253]), .A2(n10418), .B1(
        i_data_bus[157]), .B2(n10417), .ZN(n7808) );
  AOI22D1BWP30P140LVT U11440 ( .A1(i_data_bus[221]), .A2(n10419), .B1(
        i_data_bus[189]), .B2(n10420), .ZN(n7807) );
  ND2D1BWP30P140LVT U11441 ( .A1(n7808), .A2(n7807), .ZN(N13934) );
  AOI22D1BWP30P140LVT U11442 ( .A1(i_data_bus[217]), .A2(n10419), .B1(
        i_data_bus[153]), .B2(n10417), .ZN(n7810) );
  AOI22D1BWP30P140LVT U11443 ( .A1(i_data_bus[249]), .A2(n10418), .B1(
        i_data_bus[185]), .B2(n10420), .ZN(n7809) );
  ND2D1BWP30P140LVT U11444 ( .A1(n7810), .A2(n7809), .ZN(N13930) );
  AOI22D1BWP30P140LVT U11445 ( .A1(i_data_bus[742]), .A2(n10500), .B1(
        i_data_bus[678]), .B2(n10499), .ZN(n7812) );
  AOI22D1BWP30P140LVT U11446 ( .A1(i_data_bus[646]), .A2(n10498), .B1(
        i_data_bus[710]), .B2(n10497), .ZN(n7811) );
  ND2D1BWP30P140LVT U11447 ( .A1(n7812), .A2(n7811), .ZN(N9153) );
  AOI22D1BWP30P140LVT U11448 ( .A1(i_data_bus[648]), .A2(n10498), .B1(
        i_data_bus[680]), .B2(n10499), .ZN(n7814) );
  AOI22D1BWP30P140LVT U11449 ( .A1(i_data_bus[744]), .A2(n10500), .B1(
        i_data_bus[712]), .B2(n10497), .ZN(n7813) );
  ND2D1BWP30P140LVT U11450 ( .A1(n7814), .A2(n7813), .ZN(N9155) );
  AOI22D1BWP30P140LVT U11451 ( .A1(i_data_bus[663]), .A2(n10498), .B1(
        i_data_bus[759]), .B2(n10500), .ZN(n7816) );
  AOI22D1BWP30P140LVT U11452 ( .A1(i_data_bus[695]), .A2(n10499), .B1(
        i_data_bus[727]), .B2(n10497), .ZN(n7815) );
  ND2D1BWP30P140LVT U11453 ( .A1(n7816), .A2(n7815), .ZN(N9170) );
  AOI22D1BWP30P140LVT U11454 ( .A1(i_data_bus[660]), .A2(n10498), .B1(
        i_data_bus[756]), .B2(n10500), .ZN(n7818) );
  AOI22D1BWP30P140LVT U11455 ( .A1(i_data_bus[692]), .A2(n10499), .B1(
        i_data_bus[724]), .B2(n10497), .ZN(n7817) );
  ND2D1BWP30P140LVT U11456 ( .A1(n7818), .A2(n7817), .ZN(N9167) );
  AOI22D1BWP30P140LVT U11457 ( .A1(i_data_bus[749]), .A2(n10500), .B1(
        i_data_bus[685]), .B2(n10499), .ZN(n7820) );
  AOI22D1BWP30P140LVT U11458 ( .A1(i_data_bus[653]), .A2(n10498), .B1(
        i_data_bus[717]), .B2(n10497), .ZN(n7819) );
  ND2D1BWP30P140LVT U11459 ( .A1(n7820), .A2(n7819), .ZN(N9160) );
  AOI22D1BWP30P140LVT U11460 ( .A1(i_data_bus[657]), .A2(n10498), .B1(
        i_data_bus[753]), .B2(n10500), .ZN(n7822) );
  AOI22D1BWP30P140LVT U11461 ( .A1(i_data_bus[689]), .A2(n10499), .B1(
        i_data_bus[721]), .B2(n10497), .ZN(n7821) );
  ND2D1BWP30P140LVT U11462 ( .A1(n7822), .A2(n7821), .ZN(N9164) );
  AOI22D1BWP30P140LVT U11463 ( .A1(i_data_bus[667]), .A2(n10498), .B1(
        i_data_bus[699]), .B2(n10499), .ZN(n7824) );
  AOI22D1BWP30P140LVT U11464 ( .A1(i_data_bus[763]), .A2(n10500), .B1(
        i_data_bus[731]), .B2(n10497), .ZN(n7823) );
  ND2D1BWP30P140LVT U11465 ( .A1(n7824), .A2(n7823), .ZN(N9174) );
  AOI22D1BWP30P140LVT U11466 ( .A1(i_data_bus[665]), .A2(n10498), .B1(
        i_data_bus[697]), .B2(n10499), .ZN(n7826) );
  AOI22D1BWP30P140LVT U11467 ( .A1(i_data_bus[761]), .A2(n10500), .B1(
        i_data_bus[729]), .B2(n10497), .ZN(n7825) );
  ND2D1BWP30P140LVT U11468 ( .A1(n7826), .A2(n7825), .ZN(N9172) );
  AOI22D1BWP30P140LVT U11469 ( .A1(i_data_bus[698]), .A2(n10499), .B1(
        i_data_bus[762]), .B2(n10500), .ZN(n7828) );
  AOI22D1BWP30P140LVT U11470 ( .A1(i_data_bus[666]), .A2(n10498), .B1(
        i_data_bus[730]), .B2(n10497), .ZN(n7827) );
  ND2D1BWP30P140LVT U11471 ( .A1(n7828), .A2(n7827), .ZN(N9173) );
  AOI22D1BWP30P140LVT U11472 ( .A1(i_data_bus[650]), .A2(n10498), .B1(
        i_data_bus[682]), .B2(n10499), .ZN(n7830) );
  AOI22D1BWP30P140LVT U11473 ( .A1(i_data_bus[746]), .A2(n10500), .B1(
        i_data_bus[714]), .B2(n10497), .ZN(n7829) );
  ND2D1BWP30P140LVT U11474 ( .A1(n7830), .A2(n7829), .ZN(N9157) );
  NR4D1BWP30P140LVT U11475 ( .A1(i_cmd[7]), .A2(n7831), .A3(n10014), .A4(n7832), .ZN(n10422) );
  INR4D1BWP30P140LVT U11476 ( .A1(i_cmd[31]), .B1(i_cmd[15]), .B2(n10019), 
        .B3(n7834), .ZN(n10424) );
  AOI22D1BWP30P140LVT U11477 ( .A1(i_data_bus[73]), .A2(n10422), .B1(
        i_data_bus[105]), .B2(n10424), .ZN(n7836) );
  NR4D1BWP30P140LVT U11478 ( .A1(i_cmd[23]), .A2(n10013), .A3(n7833), .A4(
        n7832), .ZN(n10421) );
  INR4D1BWP30P140LVT U11479 ( .A1(i_cmd[15]), .B1(i_cmd[31]), .B2(n10018), 
        .B3(n7834), .ZN(n10423) );
  AOI22D1BWP30P140LVT U11480 ( .A1(i_data_bus[9]), .A2(n10421), .B1(
        i_data_bus[41]), .B2(n10423), .ZN(n7835) );
  ND2D1BWP30P140LVT U11481 ( .A1(n7836), .A2(n7835), .ZN(N13698) );
  AOI22D1BWP30P140LVT U11482 ( .A1(i_data_bus[23]), .A2(n10421), .B1(
        i_data_bus[119]), .B2(n10424), .ZN(n7838) );
  AOI22D1BWP30P140LVT U11483 ( .A1(i_data_bus[87]), .A2(n10422), .B1(
        i_data_bus[55]), .B2(n10423), .ZN(n7837) );
  ND2D1BWP30P140LVT U11484 ( .A1(n7838), .A2(n7837), .ZN(N13712) );
  AOI22D1BWP30P140LVT U11485 ( .A1(i_data_bus[122]), .A2(n10424), .B1(
        i_data_bus[26]), .B2(n10421), .ZN(n7840) );
  AOI22D1BWP30P140LVT U11486 ( .A1(i_data_bus[90]), .A2(n10422), .B1(
        i_data_bus[58]), .B2(n10423), .ZN(n7839) );
  ND2D1BWP30P140LVT U11487 ( .A1(n7840), .A2(n7839), .ZN(N13715) );
  AOI22D1BWP30P140LVT U11488 ( .A1(i_data_bus[110]), .A2(n10424), .B1(
        i_data_bus[78]), .B2(n10422), .ZN(n7842) );
  AOI22D1BWP30P140LVT U11489 ( .A1(i_data_bus[14]), .A2(n10421), .B1(
        i_data_bus[46]), .B2(n10423), .ZN(n7841) );
  ND2D1BWP30P140LVT U11490 ( .A1(n7842), .A2(n7841), .ZN(N13703) );
  AOI22D1BWP30P140LVT U11491 ( .A1(i_data_bus[121]), .A2(n10424), .B1(
        i_data_bus[25]), .B2(n10421), .ZN(n7844) );
  AOI22D1BWP30P140LVT U11492 ( .A1(i_data_bus[89]), .A2(n10422), .B1(
        i_data_bus[57]), .B2(n10423), .ZN(n7843) );
  ND2D1BWP30P140LVT U11493 ( .A1(n7844), .A2(n7843), .ZN(N13714) );
  AOI22D1BWP30P140LVT U11494 ( .A1(i_data_bus[86]), .A2(n10422), .B1(
        i_data_bus[22]), .B2(n10421), .ZN(n7846) );
  AOI22D1BWP30P140LVT U11495 ( .A1(i_data_bus[118]), .A2(n10424), .B1(
        i_data_bus[54]), .B2(n10423), .ZN(n7845) );
  ND2D1BWP30P140LVT U11496 ( .A1(n7846), .A2(n7845), .ZN(N13711) );
  AOI22D1BWP30P140LVT U11497 ( .A1(i_data_bus[4]), .A2(n10421), .B1(
        i_data_bus[68]), .B2(n10422), .ZN(n7848) );
  AOI22D1BWP30P140LVT U11498 ( .A1(i_data_bus[100]), .A2(n10424), .B1(
        i_data_bus[36]), .B2(n10423), .ZN(n7847) );
  ND2D1BWP30P140LVT U11499 ( .A1(n7848), .A2(n7847), .ZN(N13693) );
  AOI22D1BWP30P140LVT U11500 ( .A1(i_data_bus[120]), .A2(n10424), .B1(
        i_data_bus[24]), .B2(n10421), .ZN(n7850) );
  AOI22D1BWP30P140LVT U11501 ( .A1(i_data_bus[88]), .A2(n10422), .B1(
        i_data_bus[56]), .B2(n10423), .ZN(n7849) );
  ND2D1BWP30P140LVT U11502 ( .A1(n7850), .A2(n7849), .ZN(N13713) );
  AOI22D1BWP30P140LVT U11503 ( .A1(i_data_bus[107]), .A2(n10424), .B1(
        i_data_bus[11]), .B2(n10421), .ZN(n7852) );
  AOI22D1BWP30P140LVT U11504 ( .A1(i_data_bus[75]), .A2(n10422), .B1(
        i_data_bus[43]), .B2(n10423), .ZN(n7851) );
  ND2D1BWP30P140LVT U11505 ( .A1(n7852), .A2(n7851), .ZN(N13700) );
  AOI22D1BWP30P140LVT U11506 ( .A1(i_data_bus[33]), .A2(n10423), .B1(
        i_data_bus[97]), .B2(n10424), .ZN(n7854) );
  AOI22D1BWP30P140LVT U11507 ( .A1(i_data_bus[65]), .A2(n10422), .B1(
        i_data_bus[1]), .B2(n10421), .ZN(n7853) );
  ND2D1BWP30P140LVT U11508 ( .A1(n7854), .A2(n7853), .ZN(N13690) );
  AOI22D1BWP30P140LVT U11509 ( .A1(i_data_bus[127]), .A2(n10424), .B1(
        i_data_bus[63]), .B2(n10423), .ZN(n7856) );
  AOI22D1BWP30P140LVT U11510 ( .A1(i_data_bus[95]), .A2(n10422), .B1(
        i_data_bus[31]), .B2(n10421), .ZN(n7855) );
  ND2D1BWP30P140LVT U11511 ( .A1(n7856), .A2(n7855), .ZN(N13720) );
  AOI22D1BWP30P140LVT U11512 ( .A1(i_data_bus[60]), .A2(n10423), .B1(
        i_data_bus[124]), .B2(n10424), .ZN(n7858) );
  AOI22D1BWP30P140LVT U11513 ( .A1(i_data_bus[92]), .A2(n10422), .B1(
        i_data_bus[28]), .B2(n10421), .ZN(n7857) );
  ND2D1BWP30P140LVT U11514 ( .A1(n7858), .A2(n7857), .ZN(N13717) );
  AOI22D1BWP30P140LVT U11515 ( .A1(i_data_bus[104]), .A2(n10424), .B1(
        i_data_bus[72]), .B2(n10422), .ZN(n7860) );
  AOI22D1BWP30P140LVT U11516 ( .A1(i_data_bus[40]), .A2(n10423), .B1(
        i_data_bus[8]), .B2(n10421), .ZN(n7859) );
  ND2D1BWP30P140LVT U11517 ( .A1(n7860), .A2(n7859), .ZN(N13697) );
  AOI22D1BWP30P140LVT U11518 ( .A1(i_data_bus[94]), .A2(n10422), .B1(
        i_data_bus[62]), .B2(n10423), .ZN(n7862) );
  AOI22D1BWP30P140LVT U11519 ( .A1(i_data_bus[126]), .A2(n10424), .B1(
        i_data_bus[30]), .B2(n10421), .ZN(n7861) );
  ND2D1BWP30P140LVT U11520 ( .A1(n7862), .A2(n7861), .ZN(N13719) );
  AOI22D1BWP30P140LVT U11521 ( .A1(i_data_bus[66]), .A2(n10422), .B1(
        i_data_bus[98]), .B2(n10424), .ZN(n7864) );
  AOI22D1BWP30P140LVT U11522 ( .A1(i_data_bus[34]), .A2(n10423), .B1(
        i_data_bus[2]), .B2(n10421), .ZN(n7863) );
  ND2D1BWP30P140LVT U11523 ( .A1(n7864), .A2(n7863), .ZN(N13691) );
  AOI22D1BWP30P140LVT U11524 ( .A1(i_data_bus[517]), .A2(n10438), .B1(
        i_data_bus[613]), .B2(n10440), .ZN(n7866) );
  AOI22D1BWP30P140LVT U11525 ( .A1(i_data_bus[549]), .A2(n10439), .B1(
        i_data_bus[581]), .B2(n10437), .ZN(n7865) );
  ND2D1BWP30P140LVT U11526 ( .A1(n7866), .A2(n7865), .ZN(N12684) );
  AOI22D1BWP30P140LVT U11527 ( .A1(i_data_bus[81]), .A2(n10422), .B1(
        i_data_bus[113]), .B2(n10424), .ZN(n7868) );
  AOI22D1BWP30P140LVT U11528 ( .A1(i_data_bus[49]), .A2(n10423), .B1(
        i_data_bus[17]), .B2(n10421), .ZN(n7867) );
  ND2D1BWP30P140LVT U11529 ( .A1(n7868), .A2(n7867), .ZN(N13706) );
  AOI22D1BWP30P140LVT U11530 ( .A1(i_data_bus[76]), .A2(n10422), .B1(
        i_data_bus[108]), .B2(n10424), .ZN(n7870) );
  AOI22D1BWP30P140LVT U11531 ( .A1(i_data_bus[44]), .A2(n10423), .B1(
        i_data_bus[12]), .B2(n10421), .ZN(n7869) );
  ND2D1BWP30P140LVT U11532 ( .A1(n7870), .A2(n7869), .ZN(N13701) );
  AOI22D1BWP30P140LVT U11533 ( .A1(i_data_bus[37]), .A2(n10423), .B1(
        i_data_bus[101]), .B2(n10424), .ZN(n7872) );
  AOI22D1BWP30P140LVT U11534 ( .A1(i_data_bus[69]), .A2(n10422), .B1(
        i_data_bus[5]), .B2(n10421), .ZN(n7871) );
  ND2D1BWP30P140LVT U11535 ( .A1(n7872), .A2(n7871), .ZN(N13694) );
  AOI22D1BWP30P140LVT U11536 ( .A1(i_data_bus[524]), .A2(n10438), .B1(
        i_data_bus[620]), .B2(n10440), .ZN(n7874) );
  AOI22D1BWP30P140LVT U11537 ( .A1(i_data_bus[556]), .A2(n10439), .B1(
        i_data_bus[588]), .B2(n10437), .ZN(n7873) );
  ND2D1BWP30P140LVT U11538 ( .A1(n7874), .A2(n7873), .ZN(N12691) );
  AOI22D1BWP30P140LVT U11539 ( .A1(i_data_bus[48]), .A2(n10423), .B1(
        i_data_bus[112]), .B2(n10424), .ZN(n7876) );
  AOI22D1BWP30P140LVT U11540 ( .A1(i_data_bus[80]), .A2(n10422), .B1(
        i_data_bus[16]), .B2(n10421), .ZN(n7875) );
  ND2D1BWP30P140LVT U11541 ( .A1(n7876), .A2(n7875), .ZN(N13705) );
  AOI22D1BWP30P140LVT U11542 ( .A1(i_data_bus[35]), .A2(n10423), .B1(
        i_data_bus[99]), .B2(n10424), .ZN(n7878) );
  AOI22D1BWP30P140LVT U11543 ( .A1(i_data_bus[67]), .A2(n10422), .B1(
        i_data_bus[3]), .B2(n10421), .ZN(n7877) );
  ND2D1BWP30P140LVT U11544 ( .A1(n7878), .A2(n7877), .ZN(N13692) );
  AOI22D1BWP30P140LVT U11545 ( .A1(i_data_bus[116]), .A2(n10424), .B1(
        i_data_bus[84]), .B2(n10422), .ZN(n7880) );
  AOI22D1BWP30P140LVT U11546 ( .A1(i_data_bus[52]), .A2(n10423), .B1(
        i_data_bus[20]), .B2(n10421), .ZN(n7879) );
  ND2D1BWP30P140LVT U11547 ( .A1(n7880), .A2(n7879), .ZN(N13709) );
  AOI22D1BWP30P140LVT U11548 ( .A1(i_data_bus[82]), .A2(n10422), .B1(
        i_data_bus[50]), .B2(n10423), .ZN(n7882) );
  AOI22D1BWP30P140LVT U11549 ( .A1(i_data_bus[114]), .A2(n10424), .B1(
        i_data_bus[18]), .B2(n10421), .ZN(n7881) );
  ND2D1BWP30P140LVT U11550 ( .A1(n7882), .A2(n7881), .ZN(N13707) );
  AOI22D1BWP30P140LVT U11551 ( .A1(i_data_bus[109]), .A2(n10424), .B1(
        i_data_bus[77]), .B2(n10422), .ZN(n7884) );
  AOI22D1BWP30P140LVT U11552 ( .A1(i_data_bus[45]), .A2(n10423), .B1(
        i_data_bus[13]), .B2(n10421), .ZN(n7883) );
  ND2D1BWP30P140LVT U11553 ( .A1(n7884), .A2(n7883), .ZN(N13702) );
  AOI22D1BWP30P140LVT U11554 ( .A1(i_data_bus[519]), .A2(n10438), .B1(
        i_data_bus[615]), .B2(n10440), .ZN(n7886) );
  AOI22D1BWP30P140LVT U11555 ( .A1(i_data_bus[551]), .A2(n10439), .B1(
        i_data_bus[583]), .B2(n10437), .ZN(n7885) );
  ND2D1BWP30P140LVT U11556 ( .A1(n7886), .A2(n7885), .ZN(N12686) );
  AOI22D1BWP30P140LVT U11557 ( .A1(i_data_bus[71]), .A2(n10422), .B1(
        i_data_bus[103]), .B2(n10424), .ZN(n7888) );
  AOI22D1BWP30P140LVT U11558 ( .A1(i_data_bus[39]), .A2(n10423), .B1(
        i_data_bus[7]), .B2(n10421), .ZN(n7887) );
  ND2D1BWP30P140LVT U11559 ( .A1(n7888), .A2(n7887), .ZN(N13696) );
  AOI22D1BWP30P140LVT U11560 ( .A1(i_data_bus[279]), .A2(n10510), .B1(
        i_data_bus[311]), .B2(n10512), .ZN(n7890) );
  AOI22D1BWP30P140LVT U11561 ( .A1(i_data_bus[375]), .A2(n10511), .B1(
        i_data_bus[343]), .B2(n10509), .ZN(n7889) );
  ND2D1BWP30P140LVT U11562 ( .A1(n7890), .A2(n7889), .ZN(N8522) );
  AOI22D1BWP30P140LVT U11563 ( .A1(i_data_bus[353]), .A2(n10511), .B1(
        i_data_bus[289]), .B2(n10512), .ZN(n7892) );
  AOI22D1BWP30P140LVT U11564 ( .A1(i_data_bus[257]), .A2(n10510), .B1(
        i_data_bus[321]), .B2(n10509), .ZN(n7891) );
  ND2D1BWP30P140LVT U11565 ( .A1(n7892), .A2(n7891), .ZN(N8500) );
  AOI22D1BWP30P140LVT U11566 ( .A1(i_data_bus[282]), .A2(n10510), .B1(
        i_data_bus[378]), .B2(n10511), .ZN(n7894) );
  AOI22D1BWP30P140LVT U11567 ( .A1(i_data_bus[314]), .A2(n10512), .B1(
        i_data_bus[346]), .B2(n10509), .ZN(n7893) );
  ND2D1BWP30P140LVT U11568 ( .A1(n7894), .A2(n7893), .ZN(N8525) );
  AOI22D1BWP30P140LVT U11569 ( .A1(i_data_bus[364]), .A2(n10511), .B1(
        i_data_bus[300]), .B2(n10512), .ZN(n7896) );
  AOI22D1BWP30P140LVT U11570 ( .A1(i_data_bus[268]), .A2(n10510), .B1(
        i_data_bus[332]), .B2(n10509), .ZN(n7895) );
  ND2D1BWP30P140LVT U11571 ( .A1(n7896), .A2(n7895), .ZN(N8511) );
  AOI22D1BWP30P140LVT U11572 ( .A1(i_data_bus[281]), .A2(n10510), .B1(
        i_data_bus[377]), .B2(n10511), .ZN(n7898) );
  AOI22D1BWP30P140LVT U11573 ( .A1(i_data_bus[313]), .A2(n10512), .B1(
        i_data_bus[345]), .B2(n10509), .ZN(n7897) );
  ND2D1BWP30P140LVT U11574 ( .A1(n7898), .A2(n7897), .ZN(N8524) );
  AOI22D1BWP30P140LVT U11575 ( .A1(i_data_bus[284]), .A2(n10510), .B1(
        i_data_bus[316]), .B2(n10512), .ZN(n7900) );
  AOI22D1BWP30P140LVT U11576 ( .A1(i_data_bus[380]), .A2(n10511), .B1(
        i_data_bus[348]), .B2(n10509), .ZN(n7899) );
  ND2D1BWP30P140LVT U11577 ( .A1(n7900), .A2(n7899), .ZN(N8527) );
  AOI22D1BWP30P140LVT U11578 ( .A1(i_data_bus[275]), .A2(n10510), .B1(
        i_data_bus[371]), .B2(n10511), .ZN(n7902) );
  AOI22D1BWP30P140LVT U11579 ( .A1(i_data_bus[307]), .A2(n10512), .B1(
        i_data_bus[339]), .B2(n10509), .ZN(n7901) );
  ND2D1BWP30P140LVT U11580 ( .A1(n7902), .A2(n7901), .ZN(N8518) );
  AOI22D1BWP30P140LVT U11581 ( .A1(i_data_bus[267]), .A2(n10510), .B1(
        i_data_bus[299]), .B2(n10512), .ZN(n7904) );
  AOI22D1BWP30P140LVT U11582 ( .A1(i_data_bus[363]), .A2(n10511), .B1(
        i_data_bus[331]), .B2(n10509), .ZN(n7903) );
  ND2D1BWP30P140LVT U11583 ( .A1(n7904), .A2(n7903), .ZN(N8510) );
  AOI22D1BWP30P140LVT U11584 ( .A1(i_data_bus[561]), .A2(n10439), .B1(
        i_data_bus[625]), .B2(n10440), .ZN(n7906) );
  AOI22D1BWP30P140LVT U11585 ( .A1(i_data_bus[593]), .A2(n10437), .B1(
        i_data_bus[529]), .B2(n10438), .ZN(n7905) );
  ND2D1BWP30P140LVT U11586 ( .A1(n7906), .A2(n7905), .ZN(N12696) );
  AOI22D1BWP30P140LVT U11587 ( .A1(i_data_bus[590]), .A2(n10437), .B1(
        i_data_bus[622]), .B2(n10440), .ZN(n7908) );
  AOI22D1BWP30P140LVT U11588 ( .A1(i_data_bus[558]), .A2(n10439), .B1(
        i_data_bus[526]), .B2(n10438), .ZN(n7907) );
  ND2D1BWP30P140LVT U11589 ( .A1(n7908), .A2(n7907), .ZN(N12693) );
  AOI22D1BWP30P140LVT U11590 ( .A1(i_data_bus[569]), .A2(n10439), .B1(
        i_data_bus[633]), .B2(n10440), .ZN(n7910) );
  AOI22D1BWP30P140LVT U11591 ( .A1(i_data_bus[601]), .A2(n10437), .B1(
        i_data_bus[537]), .B2(n10438), .ZN(n7909) );
  ND2D1BWP30P140LVT U11592 ( .A1(n7910), .A2(n7909), .ZN(N12704) );
  AOI22D1BWP30P140LVT U11593 ( .A1(i_data_bus[559]), .A2(n10439), .B1(
        i_data_bus[623]), .B2(n10440), .ZN(n7912) );
  AOI22D1BWP30P140LVT U11594 ( .A1(i_data_bus[591]), .A2(n10437), .B1(
        i_data_bus[527]), .B2(n10438), .ZN(n7911) );
  ND2D1BWP30P140LVT U11595 ( .A1(n7912), .A2(n7911), .ZN(N12694) );
  AOI22D1BWP30P140LVT U11596 ( .A1(i_data_bus[322]), .A2(n10544), .B1(
        i_data_bus[354]), .B2(n10542), .ZN(n7914) );
  AOI22D1BWP30P140LVT U11597 ( .A1(i_data_bus[258]), .A2(n10543), .B1(
        i_data_bus[290]), .B2(n10541), .ZN(n7913) );
  ND2D1BWP30P140LVT U11598 ( .A1(n7914), .A2(n7913), .ZN(N6627) );
  AOI22D1BWP30P140LVT U11599 ( .A1(i_data_bus[270]), .A2(n10543), .B1(
        i_data_bus[366]), .B2(n10542), .ZN(n7916) );
  AOI22D1BWP30P140LVT U11600 ( .A1(i_data_bus[334]), .A2(n10544), .B1(
        i_data_bus[302]), .B2(n10541), .ZN(n7915) );
  ND2D1BWP30P140LVT U11601 ( .A1(n7916), .A2(n7915), .ZN(N6639) );
  AOI22D1BWP30P140LVT U11602 ( .A1(i_data_bus[287]), .A2(n10543), .B1(
        i_data_bus[383]), .B2(n10542), .ZN(n7918) );
  AOI22D1BWP30P140LVT U11603 ( .A1(i_data_bus[351]), .A2(n10544), .B1(
        i_data_bus[319]), .B2(n10541), .ZN(n7917) );
  ND2D1BWP30P140LVT U11604 ( .A1(n7918), .A2(n7917), .ZN(N6656) );
  AOI22D1BWP30P140LVT U11605 ( .A1(i_data_bus[257]), .A2(n10543), .B1(
        i_data_bus[353]), .B2(n10542), .ZN(n7920) );
  AOI22D1BWP30P140LVT U11606 ( .A1(i_data_bus[321]), .A2(n10544), .B1(
        i_data_bus[289]), .B2(n10541), .ZN(n7919) );
  ND2D1BWP30P140LVT U11607 ( .A1(n7920), .A2(n7919), .ZN(N6626) );
  AOI22D1BWP30P140LVT U11608 ( .A1(i_data_bus[324]), .A2(n10544), .B1(
        i_data_bus[356]), .B2(n10542), .ZN(n7922) );
  AOI22D1BWP30P140LVT U11609 ( .A1(i_data_bus[292]), .A2(n10541), .B1(
        i_data_bus[260]), .B2(n10543), .ZN(n7921) );
  ND2D1BWP30P140LVT U11610 ( .A1(n7922), .A2(n7921), .ZN(N6629) );
  AOI22D1BWP30P140LVT U11611 ( .A1(i_data_bus[325]), .A2(n10544), .B1(
        i_data_bus[357]), .B2(n10542), .ZN(n7924) );
  AOI22D1BWP30P140LVT U11612 ( .A1(i_data_bus[293]), .A2(n10541), .B1(
        i_data_bus[261]), .B2(n10543), .ZN(n7923) );
  ND2D1BWP30P140LVT U11613 ( .A1(n7924), .A2(n7923), .ZN(N6630) );
  AOI22D1BWP30P140LVT U11614 ( .A1(i_data_bus[275]), .A2(n10543), .B1(
        i_data_bus[371]), .B2(n10542), .ZN(n7926) );
  AOI22D1BWP30P140LVT U11615 ( .A1(i_data_bus[307]), .A2(n10541), .B1(
        i_data_bus[339]), .B2(n10544), .ZN(n7925) );
  ND2D1BWP30P140LVT U11616 ( .A1(n7926), .A2(n7925), .ZN(N6644) );
  AOI22D1BWP30P140LVT U11617 ( .A1(i_data_bus[298]), .A2(n10541), .B1(
        i_data_bus[362]), .B2(n10542), .ZN(n7928) );
  AOI22D1BWP30P140LVT U11618 ( .A1(i_data_bus[266]), .A2(n10543), .B1(
        i_data_bus[330]), .B2(n10544), .ZN(n7927) );
  ND2D1BWP30P140LVT U11619 ( .A1(n7928), .A2(n7927), .ZN(N6635) );
  AOI22D1BWP30P140LVT U11620 ( .A1(i_data_bus[305]), .A2(n10541), .B1(
        i_data_bus[369]), .B2(n10542), .ZN(n7930) );
  AOI22D1BWP30P140LVT U11621 ( .A1(i_data_bus[273]), .A2(n10543), .B1(
        i_data_bus[337]), .B2(n10544), .ZN(n7929) );
  ND2D1BWP30P140LVT U11622 ( .A1(n7930), .A2(n7929), .ZN(N6642) );
  AOI22D1BWP30P140LVT U11623 ( .A1(i_data_bus[719]), .A2(n10434), .B1(
        i_data_bus[687]), .B2(n10436), .ZN(n7932) );
  AOI22D1BWP30P140LVT U11624 ( .A1(i_data_bus[751]), .A2(n10433), .B1(
        i_data_bus[655]), .B2(n10435), .ZN(n7931) );
  ND2D1BWP30P140LVT U11625 ( .A1(n7932), .A2(n7931), .ZN(N12910) );
  AOI22D1BWP30P140LVT U11626 ( .A1(i_data_bus[766]), .A2(n10433), .B1(
        i_data_bus[702]), .B2(n10436), .ZN(n7934) );
  AOI22D1BWP30P140LVT U11627 ( .A1(i_data_bus[734]), .A2(n10434), .B1(
        i_data_bus[670]), .B2(n10435), .ZN(n7933) );
  ND2D1BWP30P140LVT U11628 ( .A1(n7934), .A2(n7933), .ZN(N12925) );
  AOI22D1BWP30P140LVT U11629 ( .A1(i_data_bus[709]), .A2(n10434), .B1(
        i_data_bus[741]), .B2(n10433), .ZN(n7936) );
  AOI22D1BWP30P140LVT U11630 ( .A1(i_data_bus[677]), .A2(n10436), .B1(
        i_data_bus[645]), .B2(n10435), .ZN(n7935) );
  ND2D1BWP30P140LVT U11631 ( .A1(n7936), .A2(n7935), .ZN(N12900) );
  AOI22D1BWP30P140LVT U11632 ( .A1(i_data_bus[686]), .A2(n10436), .B1(
        i_data_bus[750]), .B2(n10433), .ZN(n7938) );
  AOI22D1BWP30P140LVT U11633 ( .A1(i_data_bus[718]), .A2(n10434), .B1(
        i_data_bus[654]), .B2(n10435), .ZN(n7937) );
  ND2D1BWP30P140LVT U11634 ( .A1(n7938), .A2(n7937), .ZN(N12909) );
  AOI22D1BWP30P140LVT U11635 ( .A1(i_data_bus[679]), .A2(n10436), .B1(
        i_data_bus[743]), .B2(n10433), .ZN(n7940) );
  AOI22D1BWP30P140LVT U11636 ( .A1(i_data_bus[711]), .A2(n10434), .B1(
        i_data_bus[647]), .B2(n10435), .ZN(n7939) );
  ND2D1BWP30P140LVT U11637 ( .A1(n7940), .A2(n7939), .ZN(N12902) );
  AOI22D1BWP30P140LVT U11638 ( .A1(i_data_bus[704]), .A2(n10434), .B1(
        i_data_bus[736]), .B2(n10433), .ZN(n7942) );
  AOI22D1BWP30P140LVT U11639 ( .A1(i_data_bus[672]), .A2(n10436), .B1(
        i_data_bus[640]), .B2(n10435), .ZN(n7941) );
  ND2D1BWP30P140LVT U11640 ( .A1(n7942), .A2(n7941), .ZN(N12895) );
  AOI22D1BWP30P140LVT U11641 ( .A1(i_data_bus[725]), .A2(n10434), .B1(
        i_data_bus[757]), .B2(n10433), .ZN(n7944) );
  AOI22D1BWP30P140LVT U11642 ( .A1(i_data_bus[693]), .A2(n10436), .B1(
        i_data_bus[661]), .B2(n10435), .ZN(n7943) );
  ND2D1BWP30P140LVT U11643 ( .A1(n7944), .A2(n7943), .ZN(N12916) );
  AOI22D1BWP30P140LVT U11644 ( .A1(i_data_bus[728]), .A2(n10434), .B1(
        i_data_bus[760]), .B2(n10433), .ZN(n7946) );
  AOI22D1BWP30P140LVT U11645 ( .A1(i_data_bus[696]), .A2(n10436), .B1(
        i_data_bus[664]), .B2(n10435), .ZN(n7945) );
  ND2D1BWP30P140LVT U11646 ( .A1(n7946), .A2(n7945), .ZN(N12919) );
  AOI22D1BWP30P140LVT U11647 ( .A1(i_data_bus[713]), .A2(n10434), .B1(
        i_data_bus[745]), .B2(n10433), .ZN(n7948) );
  AOI22D1BWP30P140LVT U11648 ( .A1(i_data_bus[681]), .A2(n10436), .B1(
        i_data_bus[649]), .B2(n10435), .ZN(n7947) );
  ND2D1BWP30P140LVT U11649 ( .A1(n7948), .A2(n7947), .ZN(N12904) );
  AOI22D1BWP30P140LVT U11650 ( .A1(i_data_bus[703]), .A2(n10436), .B1(
        i_data_bus[767]), .B2(n10433), .ZN(n7950) );
  AOI22D1BWP30P140LVT U11651 ( .A1(i_data_bus[735]), .A2(n10434), .B1(
        i_data_bus[671]), .B2(n10435), .ZN(n7949) );
  ND2D1BWP30P140LVT U11652 ( .A1(n7950), .A2(n7949), .ZN(N12926) );
  AOI22D1BWP30P140LVT U11653 ( .A1(i_data_bus[389]), .A2(n10441), .B1(
        i_data_bus[453]), .B2(n10442), .ZN(n7952) );
  AOI22D1BWP30P140LVT U11654 ( .A1(i_data_bus[485]), .A2(n10444), .B1(
        i_data_bus[421]), .B2(n10443), .ZN(n7951) );
  ND2D1BWP30P140LVT U11655 ( .A1(n7952), .A2(n7951), .ZN(N12468) );
  AOI22D1BWP30P140LVT U11656 ( .A1(i_data_bus[483]), .A2(n10444), .B1(
        i_data_bus[387]), .B2(n10441), .ZN(n7954) );
  AOI22D1BWP30P140LVT U11657 ( .A1(i_data_bus[451]), .A2(n10442), .B1(
        i_data_bus[419]), .B2(n10443), .ZN(n7953) );
  ND2D1BWP30P140LVT U11658 ( .A1(n7954), .A2(n7953), .ZN(N12466) );
  AOI22D1BWP30P140LVT U11659 ( .A1(i_data_bus[392]), .A2(n10441), .B1(
        i_data_bus[456]), .B2(n10442), .ZN(n7956) );
  AOI22D1BWP30P140LVT U11660 ( .A1(i_data_bus[488]), .A2(n10444), .B1(
        i_data_bus[424]), .B2(n10443), .ZN(n7955) );
  ND2D1BWP30P140LVT U11661 ( .A1(n7956), .A2(n7955), .ZN(N12471) );
  AOI22D1BWP30P140LVT U11662 ( .A1(i_data_bus[487]), .A2(n10444), .B1(
        i_data_bus[391]), .B2(n10441), .ZN(n7958) );
  AOI22D1BWP30P140LVT U11663 ( .A1(i_data_bus[455]), .A2(n10442), .B1(
        i_data_bus[423]), .B2(n10443), .ZN(n7957) );
  ND2D1BWP30P140LVT U11664 ( .A1(n7958), .A2(n7957), .ZN(N12470) );
  AOI22D1BWP30P140LVT U11665 ( .A1(i_data_bus[465]), .A2(n10442), .B1(
        i_data_bus[497]), .B2(n10444), .ZN(n7960) );
  AOI22D1BWP30P140LVT U11666 ( .A1(i_data_bus[401]), .A2(n10441), .B1(
        i_data_bus[433]), .B2(n10443), .ZN(n7959) );
  ND2D1BWP30P140LVT U11667 ( .A1(n7960), .A2(n7959), .ZN(N12480) );
  AOI22D1BWP30P140LVT U11668 ( .A1(i_data_bus[489]), .A2(n10444), .B1(
        i_data_bus[457]), .B2(n10442), .ZN(n7962) );
  AOI22D1BWP30P140LVT U11669 ( .A1(i_data_bus[393]), .A2(n10441), .B1(
        i_data_bus[425]), .B2(n10443), .ZN(n7961) );
  ND2D1BWP30P140LVT U11670 ( .A1(n7962), .A2(n7961), .ZN(N12472) );
  AOI22D1BWP30P140LVT U11671 ( .A1(i_data_bus[578]), .A2(n10565), .B1(
        i_data_bus[546]), .B2(n10567), .ZN(n7964) );
  AOI22D1BWP30P140LVT U11672 ( .A1(i_data_bus[610]), .A2(n10568), .B1(
        i_data_bus[514]), .B2(n10566), .ZN(n7963) );
  ND2D1BWP30P140LVT U11673 ( .A1(n7964), .A2(n7963), .ZN(N5185) );
  AOI22D1BWP30P140LVT U11674 ( .A1(i_data_bus[594]), .A2(n10565), .B1(
        i_data_bus[562]), .B2(n10567), .ZN(n7966) );
  AOI22D1BWP30P140LVT U11675 ( .A1(i_data_bus[626]), .A2(n10568), .B1(
        i_data_bus[530]), .B2(n10566), .ZN(n7965) );
  ND2D1BWP30P140LVT U11676 ( .A1(n7966), .A2(n7965), .ZN(N5201) );
  AOI22D1BWP30P140LVT U11677 ( .A1(i_data_bus[559]), .A2(n10567), .B1(
        i_data_bus[623]), .B2(n10568), .ZN(n7968) );
  AOI22D1BWP30P140LVT U11678 ( .A1(i_data_bus[591]), .A2(n10565), .B1(
        i_data_bus[527]), .B2(n10566), .ZN(n7967) );
  ND2D1BWP30P140LVT U11679 ( .A1(n7968), .A2(n7967), .ZN(N5198) );
  AOI22D1BWP30P140LVT U11680 ( .A1(i_data_bus[560]), .A2(n10567), .B1(
        i_data_bus[624]), .B2(n10568), .ZN(n7970) );
  AOI22D1BWP30P140LVT U11681 ( .A1(i_data_bus[592]), .A2(n10565), .B1(
        i_data_bus[528]), .B2(n10566), .ZN(n7969) );
  ND2D1BWP30P140LVT U11682 ( .A1(n7970), .A2(n7969), .ZN(N5199) );
  AOI22D1BWP30P140LVT U11683 ( .A1(i_data_bus[574]), .A2(n10567), .B1(
        i_data_bus[606]), .B2(n10565), .ZN(n7972) );
  AOI22D1BWP30P140LVT U11684 ( .A1(i_data_bus[638]), .A2(n10568), .B1(
        i_data_bus[542]), .B2(n10566), .ZN(n7971) );
  ND2D1BWP30P140LVT U11685 ( .A1(n7972), .A2(n7971), .ZN(N5213) );
  AOI22D1BWP30P140LVT U11686 ( .A1(i_data_bus[637]), .A2(n10568), .B1(
        i_data_bus[573]), .B2(n10567), .ZN(n7974) );
  AOI22D1BWP30P140LVT U11687 ( .A1(i_data_bus[605]), .A2(n10565), .B1(
        i_data_bus[541]), .B2(n10566), .ZN(n7973) );
  ND2D1BWP30P140LVT U11688 ( .A1(n7974), .A2(n7973), .ZN(N5212) );
  AOI22D1BWP30P140LVT U11689 ( .A1(i_data_bus[557]), .A2(n10567), .B1(
        i_data_bus[589]), .B2(n10565), .ZN(n7976) );
  AOI22D1BWP30P140LVT U11690 ( .A1(i_data_bus[621]), .A2(n10568), .B1(
        i_data_bus[525]), .B2(n10566), .ZN(n7975) );
  ND2D1BWP30P140LVT U11691 ( .A1(n7976), .A2(n7975), .ZN(N5196) );
  AOI22D1BWP30P140LVT U11692 ( .A1(i_data_bus[571]), .A2(n10567), .B1(
        i_data_bus[603]), .B2(n10565), .ZN(n7978) );
  AOI22D1BWP30P140LVT U11693 ( .A1(i_data_bus[635]), .A2(n10568), .B1(
        i_data_bus[539]), .B2(n10566), .ZN(n7977) );
  ND2D1BWP30P140LVT U11694 ( .A1(n7978), .A2(n7977), .ZN(N5210) );
  AOI22D1BWP30P140LVT U11695 ( .A1(i_data_bus[554]), .A2(n10567), .B1(
        i_data_bus[586]), .B2(n10565), .ZN(n7980) );
  AOI22D1BWP30P140LVT U11696 ( .A1(i_data_bus[618]), .A2(n10568), .B1(
        i_data_bus[522]), .B2(n10566), .ZN(n7979) );
  ND2D1BWP30P140LVT U11697 ( .A1(n7980), .A2(n7979), .ZN(N5193) );
  AOI22D1BWP30P140LVT U11698 ( .A1(i_data_bus[969]), .A2(n10555), .B1(
        i_data_bus[937]), .B2(n10553), .ZN(n7982) );
  AOI22D1BWP30P140LVT U11699 ( .A1(i_data_bus[1001]), .A2(n10556), .B1(
        i_data_bus[905]), .B2(n10554), .ZN(n7981) );
  ND2D1BWP30P140LVT U11700 ( .A1(n7982), .A2(n7981), .ZN(N5840) );
  AOI22D1BWP30P140LVT U11701 ( .A1(i_data_bus[998]), .A2(n10556), .B1(
        i_data_bus[966]), .B2(n10555), .ZN(n7984) );
  AOI22D1BWP30P140LVT U11702 ( .A1(i_data_bus[934]), .A2(n10553), .B1(
        i_data_bus[902]), .B2(n10554), .ZN(n7983) );
  ND2D1BWP30P140LVT U11703 ( .A1(n7984), .A2(n7983), .ZN(N5837) );
  AOI22D1BWP30P140LVT U11704 ( .A1(i_data_bus[933]), .A2(n10553), .B1(
        i_data_bus[997]), .B2(n10556), .ZN(n7986) );
  AOI22D1BWP30P140LVT U11705 ( .A1(i_data_bus[965]), .A2(n10555), .B1(
        i_data_bus[901]), .B2(n10554), .ZN(n7985) );
  ND2D1BWP30P140LVT U11706 ( .A1(n7986), .A2(n7985), .ZN(N5836) );
  AOI22D1BWP30P140LVT U11707 ( .A1(i_data_bus[936]), .A2(n10553), .B1(
        i_data_bus[1000]), .B2(n10556), .ZN(n7988) );
  AOI22D1BWP30P140LVT U11708 ( .A1(i_data_bus[968]), .A2(n10555), .B1(
        i_data_bus[904]), .B2(n10554), .ZN(n7987) );
  ND2D1BWP30P140LVT U11709 ( .A1(n7988), .A2(n7987), .ZN(N5839) );
  AOI22D1BWP30P140LVT U11710 ( .A1(i_data_bus[943]), .A2(n10553), .B1(
        i_data_bus[975]), .B2(n10555), .ZN(n7990) );
  AOI22D1BWP30P140LVT U11711 ( .A1(i_data_bus[1007]), .A2(n10556), .B1(
        i_data_bus[911]), .B2(n10554), .ZN(n7989) );
  ND2D1BWP30P140LVT U11712 ( .A1(n7990), .A2(n7989), .ZN(N5846) );
  AOI22D1BWP30P140LVT U11713 ( .A1(i_data_bus[1005]), .A2(n10556), .B1(
        i_data_bus[941]), .B2(n10553), .ZN(n7992) );
  AOI22D1BWP30P140LVT U11714 ( .A1(i_data_bus[973]), .A2(n10555), .B1(
        i_data_bus[909]), .B2(n10554), .ZN(n7991) );
  ND2D1BWP30P140LVT U11715 ( .A1(n7992), .A2(n7991), .ZN(N5844) );
  AOI22D1BWP30P140LVT U11716 ( .A1(i_data_bus[986]), .A2(n10555), .B1(
        i_data_bus[1018]), .B2(n10556), .ZN(n7994) );
  AOI22D1BWP30P140LVT U11717 ( .A1(i_data_bus[954]), .A2(n10553), .B1(
        i_data_bus[922]), .B2(n10554), .ZN(n7993) );
  ND2D1BWP30P140LVT U11718 ( .A1(n7994), .A2(n7993), .ZN(N5857) );
  AOI22D1BWP30P140LVT U11719 ( .A1(i_data_bus[123]), .A2(n10424), .B1(
        i_data_bus[59]), .B2(n10423), .ZN(n7996) );
  AOI22D1BWP30P140LVT U11720 ( .A1(i_data_bus[27]), .A2(n10421), .B1(
        i_data_bus[91]), .B2(n10422), .ZN(n7995) );
  ND2D1BWP30P140LVT U11721 ( .A1(n7996), .A2(n7995), .ZN(N13716) );
  AOI22D1BWP30P140LVT U11722 ( .A1(i_data_bus[117]), .A2(n10424), .B1(
        i_data_bus[21]), .B2(n10421), .ZN(n7998) );
  AOI22D1BWP30P140LVT U11723 ( .A1(i_data_bus[53]), .A2(n10423), .B1(
        i_data_bus[85]), .B2(n10422), .ZN(n7997) );
  ND2D1BWP30P140LVT U11724 ( .A1(n7998), .A2(n7997), .ZN(N13710) );
  AOI22D1BWP30P140LVT U11725 ( .A1(i_data_bus[15]), .A2(n10421), .B1(
        i_data_bus[47]), .B2(n10423), .ZN(n8000) );
  AOI22D1BWP30P140LVT U11726 ( .A1(i_data_bus[111]), .A2(n10424), .B1(
        i_data_bus[79]), .B2(n10422), .ZN(n7999) );
  ND2D1BWP30P140LVT U11727 ( .A1(n8000), .A2(n7999), .ZN(N13704) );
  AOI22D1BWP30P140LVT U11728 ( .A1(i_data_bus[443]), .A2(n10443), .B1(
        i_data_bus[475]), .B2(n10442), .ZN(n8002) );
  AOI22D1BWP30P140LVT U11729 ( .A1(i_data_bus[507]), .A2(n10444), .B1(
        i_data_bus[411]), .B2(n10441), .ZN(n8001) );
  ND2D1BWP30P140LVT U11730 ( .A1(n8002), .A2(n8001), .ZN(N12490) );
  AOI22D1BWP30P140LVT U11731 ( .A1(i_data_bus[470]), .A2(n10442), .B1(
        i_data_bus[438]), .B2(n10443), .ZN(n8004) );
  AOI22D1BWP30P140LVT U11732 ( .A1(i_data_bus[502]), .A2(n10444), .B1(
        i_data_bus[406]), .B2(n10441), .ZN(n8003) );
  ND2D1BWP30P140LVT U11733 ( .A1(n8004), .A2(n8003), .ZN(N12485) );
  AOI22D1BWP30P140LVT U11734 ( .A1(i_data_bus[439]), .A2(n10443), .B1(
        i_data_bus[503]), .B2(n10444), .ZN(n8006) );
  AOI22D1BWP30P140LVT U11735 ( .A1(i_data_bus[471]), .A2(n10442), .B1(
        i_data_bus[407]), .B2(n10441), .ZN(n8005) );
  ND2D1BWP30P140LVT U11736 ( .A1(n8006), .A2(n8005), .ZN(N12486) );
  AOI22D1BWP30P140LVT U11737 ( .A1(i_data_bus[482]), .A2(n10444), .B1(
        i_data_bus[450]), .B2(n10442), .ZN(n8008) );
  AOI22D1BWP30P140LVT U11738 ( .A1(i_data_bus[418]), .A2(n10443), .B1(
        i_data_bus[386]), .B2(n10441), .ZN(n8007) );
  ND2D1BWP30P140LVT U11739 ( .A1(n8008), .A2(n8007), .ZN(N12465) );
  AOI22D1BWP30P140LVT U11740 ( .A1(i_data_bus[432]), .A2(n10443), .B1(
        i_data_bus[464]), .B2(n10442), .ZN(n8010) );
  AOI22D1BWP30P140LVT U11741 ( .A1(i_data_bus[496]), .A2(n10444), .B1(
        i_data_bus[400]), .B2(n10441), .ZN(n8009) );
  ND2D1BWP30P140LVT U11742 ( .A1(n8010), .A2(n8009), .ZN(N12479) );
  AOI22D1BWP30P140LVT U11743 ( .A1(i_data_bus[422]), .A2(n10443), .B1(
        i_data_bus[454]), .B2(n10442), .ZN(n8012) );
  AOI22D1BWP30P140LVT U11744 ( .A1(i_data_bus[486]), .A2(n10444), .B1(
        i_data_bus[390]), .B2(n10441), .ZN(n8011) );
  ND2D1BWP30P140LVT U11745 ( .A1(n8012), .A2(n8011), .ZN(N12469) );
  AOI22D1BWP30P140LVT U11746 ( .A1(i_data_bus[447]), .A2(n10443), .B1(
        i_data_bus[511]), .B2(n10444), .ZN(n8014) );
  AOI22D1BWP30P140LVT U11747 ( .A1(i_data_bus[479]), .A2(n10442), .B1(
        i_data_bus[415]), .B2(n10441), .ZN(n8013) );
  ND2D1BWP30P140LVT U11748 ( .A1(n8014), .A2(n8013), .ZN(N12494) );
  AOI22D1BWP30P140LVT U11749 ( .A1(i_data_bus[492]), .A2(n10444), .B1(
        i_data_bus[428]), .B2(n10443), .ZN(n8016) );
  AOI22D1BWP30P140LVT U11750 ( .A1(i_data_bus[460]), .A2(n10442), .B1(
        i_data_bus[396]), .B2(n10441), .ZN(n8015) );
  ND2D1BWP30P140LVT U11751 ( .A1(n8016), .A2(n8015), .ZN(N12475) );
  AOI22D1BWP30P140LVT U11752 ( .A1(i_data_bus[467]), .A2(n10442), .B1(
        i_data_bus[435]), .B2(n10443), .ZN(n8018) );
  AOI22D1BWP30P140LVT U11753 ( .A1(i_data_bus[499]), .A2(n10444), .B1(
        i_data_bus[403]), .B2(n10441), .ZN(n8017) );
  ND2D1BWP30P140LVT U11754 ( .A1(n8018), .A2(n8017), .ZN(N12482) );
  AOI22D1BWP30P140LVT U11755 ( .A1(i_data_bus[151]), .A2(n10417), .B1(
        i_data_bus[215]), .B2(n10419), .ZN(n8020) );
  AOI22D1BWP30P140LVT U11756 ( .A1(i_data_bus[183]), .A2(n10420), .B1(
        i_data_bus[247]), .B2(n10418), .ZN(n8019) );
  ND2D1BWP30P140LVT U11757 ( .A1(n8020), .A2(n8019), .ZN(N13928) );
  AOI22D1BWP30P140LVT U11758 ( .A1(i_data_bus[366]), .A2(n10445), .B1(
        i_data_bus[302]), .B2(n10448), .ZN(n8022) );
  AOI22D1BWP30P140LVT U11759 ( .A1(i_data_bus[270]), .A2(n10447), .B1(
        i_data_bus[334]), .B2(n10446), .ZN(n8021) );
  ND2D1BWP30P140LVT U11760 ( .A1(n8022), .A2(n8021), .ZN(N12261) );
  AOI22D1BWP30P140LVT U11761 ( .A1(i_data_bus[178]), .A2(n10420), .B1(
        i_data_bus[210]), .B2(n10419), .ZN(n8024) );
  AOI22D1BWP30P140LVT U11762 ( .A1(i_data_bus[146]), .A2(n10417), .B1(
        i_data_bus[242]), .B2(n10418), .ZN(n8023) );
  ND2D1BWP30P140LVT U11763 ( .A1(n8024), .A2(n8023), .ZN(N13923) );
  AOI22D1BWP30P140LVT U11764 ( .A1(i_data_bus[380]), .A2(n10445), .B1(
        i_data_bus[316]), .B2(n10448), .ZN(n8026) );
  AOI22D1BWP30P140LVT U11765 ( .A1(i_data_bus[284]), .A2(n10447), .B1(
        i_data_bus[348]), .B2(n10446), .ZN(n8025) );
  ND2D1BWP30P140LVT U11766 ( .A1(n8026), .A2(n8025), .ZN(N12275) );
  AOI22D1BWP30P140LVT U11767 ( .A1(i_data_bus[278]), .A2(n10447), .B1(
        i_data_bus[374]), .B2(n10445), .ZN(n8028) );
  AOI22D1BWP30P140LVT U11768 ( .A1(i_data_bus[310]), .A2(n10448), .B1(
        i_data_bus[342]), .B2(n10446), .ZN(n8027) );
  ND2D1BWP30P140LVT U11769 ( .A1(n8028), .A2(n8027), .ZN(N12269) );
  AOI22D1BWP30P140LVT U11770 ( .A1(i_data_bus[205]), .A2(n10419), .B1(
        i_data_bus[141]), .B2(n10417), .ZN(n8030) );
  AOI22D1BWP30P140LVT U11771 ( .A1(i_data_bus[173]), .A2(n10420), .B1(
        i_data_bus[237]), .B2(n10418), .ZN(n8029) );
  ND2D1BWP30P140LVT U11772 ( .A1(n8030), .A2(n8029), .ZN(N13918) );
  AOI22D1BWP30P140LVT U11773 ( .A1(i_data_bus[275]), .A2(n10447), .B1(
        i_data_bus[307]), .B2(n10448), .ZN(n8032) );
  AOI22D1BWP30P140LVT U11774 ( .A1(i_data_bus[371]), .A2(n10445), .B1(
        i_data_bus[339]), .B2(n10446), .ZN(n8031) );
  ND2D1BWP30P140LVT U11775 ( .A1(n8032), .A2(n8031), .ZN(N12266) );
  AOI22D1BWP30P140LVT U11776 ( .A1(i_data_bus[358]), .A2(n10445), .B1(
        i_data_bus[294]), .B2(n10448), .ZN(n8034) );
  AOI22D1BWP30P140LVT U11777 ( .A1(i_data_bus[262]), .A2(n10447), .B1(
        i_data_bus[326]), .B2(n10446), .ZN(n8033) );
  ND2D1BWP30P140LVT U11778 ( .A1(n8034), .A2(n8033), .ZN(N12253) );
  AOI22D1BWP30P140LVT U11779 ( .A1(i_data_bus[269]), .A2(n10447), .B1(
        i_data_bus[301]), .B2(n10448), .ZN(n8036) );
  AOI22D1BWP30P140LVT U11780 ( .A1(i_data_bus[365]), .A2(n10445), .B1(
        i_data_bus[333]), .B2(n10446), .ZN(n8035) );
  ND2D1BWP30P140LVT U11781 ( .A1(n8036), .A2(n8035), .ZN(N12260) );
  AOI22D1BWP30P140LVT U11782 ( .A1(i_data_bus[355]), .A2(n10445), .B1(
        i_data_bus[259]), .B2(n10447), .ZN(n8038) );
  AOI22D1BWP30P140LVT U11783 ( .A1(i_data_bus[291]), .A2(n10448), .B1(
        i_data_bus[323]), .B2(n10446), .ZN(n8037) );
  ND2D1BWP30P140LVT U11784 ( .A1(n8038), .A2(n8037), .ZN(N12250) );
  AOI22D1BWP30P140LVT U11785 ( .A1(i_data_bus[271]), .A2(n10447), .B1(
        i_data_bus[303]), .B2(n10448), .ZN(n8040) );
  AOI22D1BWP30P140LVT U11786 ( .A1(i_data_bus[367]), .A2(n10445), .B1(
        i_data_bus[335]), .B2(n10446), .ZN(n8039) );
  ND2D1BWP30P140LVT U11787 ( .A1(n8040), .A2(n8039), .ZN(N12262) );
  AOI22D1BWP30P140LVT U11788 ( .A1(i_data_bus[311]), .A2(n10448), .B1(
        i_data_bus[375]), .B2(n10445), .ZN(n8042) );
  AOI22D1BWP30P140LVT U11789 ( .A1(i_data_bus[279]), .A2(n10447), .B1(
        i_data_bus[343]), .B2(n10446), .ZN(n8041) );
  ND2D1BWP30P140LVT U11790 ( .A1(n8042), .A2(n8041), .ZN(N12270) );
  AOI22D1BWP30P140LVT U11791 ( .A1(i_data_bus[144]), .A2(n10417), .B1(
        i_data_bus[176]), .B2(n10420), .ZN(n8044) );
  AOI22D1BWP30P140LVT U11792 ( .A1(i_data_bus[208]), .A2(n10419), .B1(
        i_data_bus[240]), .B2(n10418), .ZN(n8043) );
  ND2D1BWP30P140LVT U11793 ( .A1(n8044), .A2(n8043), .ZN(N13921) );
  AOI22D1BWP30P140LVT U11794 ( .A1(i_data_bus[281]), .A2(n10447), .B1(
        i_data_bus[377]), .B2(n10445), .ZN(n8046) );
  AOI22D1BWP30P140LVT U11795 ( .A1(i_data_bus[313]), .A2(n10448), .B1(
        i_data_bus[345]), .B2(n10446), .ZN(n8045) );
  ND2D1BWP30P140LVT U11796 ( .A1(n8046), .A2(n8045), .ZN(N12272) );
  AOI22D1BWP30P140LVT U11797 ( .A1(i_data_bus[148]), .A2(n10417), .B1(
        i_data_bus[212]), .B2(n10419), .ZN(n8048) );
  AOI22D1BWP30P140LVT U11798 ( .A1(i_data_bus[180]), .A2(n10420), .B1(
        i_data_bus[244]), .B2(n10418), .ZN(n8047) );
  ND2D1BWP30P140LVT U11799 ( .A1(n8048), .A2(n8047), .ZN(N13925) );
  AOI22D1BWP30P140LVT U11800 ( .A1(i_data_bus[282]), .A2(n10447), .B1(
        i_data_bus[378]), .B2(n10445), .ZN(n8050) );
  AOI22D1BWP30P140LVT U11801 ( .A1(i_data_bus[314]), .A2(n10448), .B1(
        i_data_bus[346]), .B2(n10446), .ZN(n8049) );
  ND2D1BWP30P140LVT U11802 ( .A1(n8050), .A2(n8049), .ZN(N12273) );
  AOI22D1BWP30P140LVT U11803 ( .A1(i_data_bus[372]), .A2(n10479), .B1(
        i_data_bus[276]), .B2(n10480), .ZN(n8052) );
  AOI22D1BWP30P140LVT U11804 ( .A1(i_data_bus[308]), .A2(n10477), .B1(
        i_data_bus[340]), .B2(n10478), .ZN(n8051) );
  ND2D1BWP30P140LVT U11805 ( .A1(n8052), .A2(n8051), .ZN(N10393) );
  AOI22D1BWP30P140LVT U11806 ( .A1(i_data_bus[181]), .A2(n10420), .B1(
        i_data_bus[213]), .B2(n10419), .ZN(n8054) );
  AOI22D1BWP30P140LVT U11807 ( .A1(i_data_bus[149]), .A2(n10417), .B1(
        i_data_bus[245]), .B2(n10418), .ZN(n8053) );
  ND2D1BWP30P140LVT U11808 ( .A1(n8054), .A2(n8053), .ZN(N13926) );
  AOI22D1BWP30P140LVT U11809 ( .A1(i_data_bus[262]), .A2(n10480), .B1(
        i_data_bus[294]), .B2(n10477), .ZN(n8056) );
  AOI22D1BWP30P140LVT U11810 ( .A1(i_data_bus[358]), .A2(n10479), .B1(
        i_data_bus[326]), .B2(n10478), .ZN(n8055) );
  ND2D1BWP30P140LVT U11811 ( .A1(n8056), .A2(n8055), .ZN(N10379) );
  AOI22D1BWP30P140LVT U11812 ( .A1(i_data_bus[359]), .A2(n10479), .B1(
        i_data_bus[263]), .B2(n10480), .ZN(n8058) );
  AOI22D1BWP30P140LVT U11813 ( .A1(i_data_bus[295]), .A2(n10477), .B1(
        i_data_bus[327]), .B2(n10478), .ZN(n8057) );
  ND2D1BWP30P140LVT U11814 ( .A1(n8058), .A2(n8057), .ZN(N10380) );
  AOI22D1BWP30P140LVT U11815 ( .A1(i_data_bus[269]), .A2(n10480), .B1(
        i_data_bus[301]), .B2(n10477), .ZN(n8060) );
  AOI22D1BWP30P140LVT U11816 ( .A1(i_data_bus[365]), .A2(n10479), .B1(
        i_data_bus[333]), .B2(n10478), .ZN(n8059) );
  ND2D1BWP30P140LVT U11817 ( .A1(n8060), .A2(n8059), .ZN(N10386) );
  AOI22D1BWP30P140LVT U11818 ( .A1(i_data_bus[363]), .A2(n10479), .B1(
        i_data_bus[299]), .B2(n10477), .ZN(n8062) );
  AOI22D1BWP30P140LVT U11819 ( .A1(i_data_bus[267]), .A2(n10480), .B1(
        i_data_bus[331]), .B2(n10478), .ZN(n8061) );
  ND2D1BWP30P140LVT U11820 ( .A1(n8062), .A2(n8061), .ZN(N10384) );
  AOI22D1BWP30P140LVT U11821 ( .A1(i_data_bus[286]), .A2(n10480), .B1(
        i_data_bus[318]), .B2(n10477), .ZN(n8064) );
  AOI22D1BWP30P140LVT U11822 ( .A1(i_data_bus[382]), .A2(n10479), .B1(
        i_data_bus[350]), .B2(n10478), .ZN(n8063) );
  ND2D1BWP30P140LVT U11823 ( .A1(n8064), .A2(n8063), .ZN(N10403) );
  AOI22D1BWP30P140LVT U11824 ( .A1(i_data_bus[355]), .A2(n10479), .B1(
        i_data_bus[259]), .B2(n10480), .ZN(n8066) );
  AOI22D1BWP30P140LVT U11825 ( .A1(i_data_bus[291]), .A2(n10477), .B1(
        i_data_bus[323]), .B2(n10478), .ZN(n8065) );
  ND2D1BWP30P140LVT U11826 ( .A1(n8066), .A2(n8065), .ZN(N10376) );
  AOI22D1BWP30P140LVT U11827 ( .A1(i_data_bus[284]), .A2(n10480), .B1(
        i_data_bus[316]), .B2(n10477), .ZN(n8068) );
  AOI22D1BWP30P140LVT U11828 ( .A1(i_data_bus[380]), .A2(n10479), .B1(
        i_data_bus[348]), .B2(n10478), .ZN(n8067) );
  ND2D1BWP30P140LVT U11829 ( .A1(n8068), .A2(n8067), .ZN(N10401) );
  AOI22D1BWP30P140LVT U11830 ( .A1(i_data_bus[10]), .A2(n10615), .B1(
        i_data_bus[42]), .B2(n10614), .ZN(n8070) );
  AOI22D1BWP30P140LVT U11831 ( .A1(i_data_bus[74]), .A2(n10613), .B1(
        i_data_bus[106]), .B2(n10616), .ZN(n8069) );
  ND2D1BWP30P140LVT U11832 ( .A1(n8070), .A2(n8069), .ZN(N2455) );
  AOI22D1BWP30P140LVT U11833 ( .A1(i_data_bus[80]), .A2(n10613), .B1(
        i_data_bus[16]), .B2(n10615), .ZN(n8072) );
  AOI22D1BWP30P140LVT U11834 ( .A1(i_data_bus[48]), .A2(n10614), .B1(
        i_data_bus[112]), .B2(n10616), .ZN(n8071) );
  ND2D1BWP30P140LVT U11835 ( .A1(n8072), .A2(n8071), .ZN(N2461) );
  AOI22D1BWP30P140LVT U11836 ( .A1(i_data_bus[49]), .A2(n10614), .B1(
        i_data_bus[81]), .B2(n10613), .ZN(n8074) );
  AOI22D1BWP30P140LVT U11837 ( .A1(i_data_bus[17]), .A2(n10615), .B1(
        i_data_bus[113]), .B2(n10616), .ZN(n8073) );
  ND2D1BWP30P140LVT U11838 ( .A1(n8074), .A2(n8073), .ZN(N2462) );
  AOI22D1BWP30P140LVT U11839 ( .A1(i_data_bus[93]), .A2(n10613), .B1(
        i_data_bus[29]), .B2(n10615), .ZN(n8076) );
  AOI22D1BWP30P140LVT U11840 ( .A1(i_data_bus[61]), .A2(n10614), .B1(
        i_data_bus[125]), .B2(n10616), .ZN(n8075) );
  ND2D1BWP30P140LVT U11841 ( .A1(n8076), .A2(n8075), .ZN(N2474) );
  AOI22D1BWP30P140LVT U11842 ( .A1(i_data_bus[37]), .A2(n10614), .B1(
        i_data_bus[69]), .B2(n10613), .ZN(n8078) );
  AOI22D1BWP30P140LVT U11843 ( .A1(i_data_bus[5]), .A2(n10615), .B1(
        i_data_bus[101]), .B2(n10616), .ZN(n8077) );
  ND2D1BWP30P140LVT U11844 ( .A1(n8078), .A2(n8077), .ZN(N2450) );
  AOI22D1BWP30P140LVT U11845 ( .A1(i_data_bus[47]), .A2(n10614), .B1(
        i_data_bus[79]), .B2(n10613), .ZN(n8080) );
  AOI22D1BWP30P140LVT U11846 ( .A1(i_data_bus[15]), .A2(n10615), .B1(
        i_data_bus[111]), .B2(n10616), .ZN(n8079) );
  ND2D1BWP30P140LVT U11847 ( .A1(n8080), .A2(n8079), .ZN(N2460) );
  AOI22D1BWP30P140LVT U11848 ( .A1(i_data_bus[65]), .A2(n10613), .B1(
        i_data_bus[1]), .B2(n10615), .ZN(n8082) );
  AOI22D1BWP30P140LVT U11849 ( .A1(i_data_bus[33]), .A2(n10614), .B1(
        i_data_bus[97]), .B2(n10616), .ZN(n8081) );
  ND2D1BWP30P140LVT U11850 ( .A1(n8082), .A2(n8081), .ZN(N2446) );
  AOI22D1BWP30P140LVT U11851 ( .A1(i_data_bus[626]), .A2(n10501), .B1(
        i_data_bus[562]), .B2(n10504), .ZN(n8084) );
  AOI22D1BWP30P140LVT U11852 ( .A1(i_data_bus[594]), .A2(n10502), .B1(
        i_data_bus[530]), .B2(n10503), .ZN(n8083) );
  ND2D1BWP30P140LVT U11853 ( .A1(n8084), .A2(n8083), .ZN(N8949) );
  AOI22D1BWP30P140LVT U11854 ( .A1(i_data_bus[572]), .A2(n10504), .B1(
        i_data_bus[636]), .B2(n10501), .ZN(n8086) );
  AOI22D1BWP30P140LVT U11855 ( .A1(i_data_bus[604]), .A2(n10502), .B1(
        i_data_bus[540]), .B2(n10503), .ZN(n8085) );
  ND2D1BWP30P140LVT U11856 ( .A1(n8086), .A2(n8085), .ZN(N8959) );
  AOI22D1BWP30P140LVT U11857 ( .A1(i_data_bus[552]), .A2(n10504), .B1(
        i_data_bus[584]), .B2(n10502), .ZN(n8088) );
  AOI22D1BWP30P140LVT U11858 ( .A1(i_data_bus[616]), .A2(n10501), .B1(
        i_data_bus[520]), .B2(n10503), .ZN(n8087) );
  ND2D1BWP30P140LVT U11859 ( .A1(n8088), .A2(n8087), .ZN(N8939) );
  AOI22D1BWP30P140LVT U11860 ( .A1(i_data_bus[586]), .A2(n10502), .B1(
        i_data_bus[618]), .B2(n10501), .ZN(n8090) );
  AOI22D1BWP30P140LVT U11861 ( .A1(i_data_bus[554]), .A2(n10504), .B1(
        i_data_bus[522]), .B2(n10503), .ZN(n8089) );
  ND2D1BWP30P140LVT U11862 ( .A1(n8090), .A2(n8089), .ZN(N8941) );
  AOI22D1BWP30P140LVT U11863 ( .A1(i_data_bus[550]), .A2(n10504), .B1(
        i_data_bus[582]), .B2(n10502), .ZN(n8092) );
  AOI22D1BWP30P140LVT U11864 ( .A1(i_data_bus[614]), .A2(n10501), .B1(
        i_data_bus[518]), .B2(n10503), .ZN(n8091) );
  ND2D1BWP30P140LVT U11865 ( .A1(n8092), .A2(n8091), .ZN(N8937) );
  AOI22D1BWP30P140LVT U11866 ( .A1(i_data_bus[569]), .A2(n10504), .B1(
        i_data_bus[633]), .B2(n10501), .ZN(n8094) );
  AOI22D1BWP30P140LVT U11867 ( .A1(i_data_bus[601]), .A2(n10502), .B1(
        i_data_bus[537]), .B2(n10503), .ZN(n8093) );
  ND2D1BWP30P140LVT U11868 ( .A1(n8094), .A2(n8093), .ZN(N8956) );
  AOI22D1BWP30P140LVT U11869 ( .A1(i_data_bus[568]), .A2(n10504), .B1(
        i_data_bus[632]), .B2(n10501), .ZN(n8096) );
  AOI22D1BWP30P140LVT U11870 ( .A1(i_data_bus[600]), .A2(n10502), .B1(
        i_data_bus[536]), .B2(n10503), .ZN(n8095) );
  ND2D1BWP30P140LVT U11871 ( .A1(n8096), .A2(n8095), .ZN(N8955) );
  AOI22D1BWP30P140LVT U11872 ( .A1(i_data_bus[564]), .A2(n10504), .B1(
        i_data_bus[628]), .B2(n10501), .ZN(n8098) );
  AOI22D1BWP30P140LVT U11873 ( .A1(i_data_bus[596]), .A2(n10502), .B1(
        i_data_bus[532]), .B2(n10503), .ZN(n8097) );
  ND2D1BWP30P140LVT U11874 ( .A1(n8098), .A2(n8097), .ZN(N8951) );
  AOI22D1BWP30P140LVT U11875 ( .A1(i_data_bus[630]), .A2(n10501), .B1(
        i_data_bus[598]), .B2(n10502), .ZN(n8100) );
  AOI22D1BWP30P140LVT U11876 ( .A1(i_data_bus[566]), .A2(n10504), .B1(
        i_data_bus[534]), .B2(n10503), .ZN(n8099) );
  ND2D1BWP30P140LVT U11877 ( .A1(n8100), .A2(n8099), .ZN(N8953) );
  AOI22D1BWP30P140LVT U11878 ( .A1(i_data_bus[610]), .A2(n10501), .B1(
        i_data_bus[546]), .B2(n10504), .ZN(n8102) );
  AOI22D1BWP30P140LVT U11879 ( .A1(i_data_bus[578]), .A2(n10502), .B1(
        i_data_bus[514]), .B2(n10503), .ZN(n8101) );
  ND2D1BWP30P140LVT U11880 ( .A1(n8102), .A2(n8101), .ZN(N8933) );
  AOI22D1BWP30P140LVT U11881 ( .A1(i_data_bus[570]), .A2(n10504), .B1(
        i_data_bus[634]), .B2(n10501), .ZN(n8104) );
  AOI22D1BWP30P140LVT U11882 ( .A1(i_data_bus[602]), .A2(n10502), .B1(
        i_data_bus[538]), .B2(n10503), .ZN(n8103) );
  ND2D1BWP30P140LVT U11883 ( .A1(n8104), .A2(n8103), .ZN(N8957) );
  AOI22D1BWP30P140LVT U11884 ( .A1(i_data_bus[588]), .A2(n10502), .B1(
        i_data_bus[620]), .B2(n10501), .ZN(n8106) );
  AOI22D1BWP30P140LVT U11885 ( .A1(i_data_bus[556]), .A2(n10504), .B1(
        i_data_bus[524]), .B2(n10503), .ZN(n8105) );
  ND2D1BWP30P140LVT U11886 ( .A1(n8106), .A2(n8105), .ZN(N8943) );
  AOI22D1BWP30P140LVT U11887 ( .A1(i_data_bus[100]), .A2(n10584), .B1(
        i_data_bus[4]), .B2(n10581), .ZN(n8108) );
  AOI22D1BWP30P140LVT U11888 ( .A1(i_data_bus[68]), .A2(n10582), .B1(
        i_data_bus[36]), .B2(n10583), .ZN(n8107) );
  ND2D1BWP30P140LVT U11889 ( .A1(n8108), .A2(n8107), .ZN(N4323) );
  AOI22D1BWP30P140LVT U11890 ( .A1(i_data_bus[82]), .A2(n10582), .B1(
        i_data_bus[18]), .B2(n10581), .ZN(n8110) );
  AOI22D1BWP30P140LVT U11891 ( .A1(i_data_bus[114]), .A2(n10584), .B1(
        i_data_bus[50]), .B2(n10583), .ZN(n8109) );
  ND2D1BWP30P140LVT U11892 ( .A1(n8110), .A2(n8109), .ZN(N4337) );
  AOI22D1BWP30P140LVT U11893 ( .A1(i_data_bus[121]), .A2(n10584), .B1(
        i_data_bus[25]), .B2(n10581), .ZN(n8112) );
  AOI22D1BWP30P140LVT U11894 ( .A1(i_data_bus[89]), .A2(n10582), .B1(
        i_data_bus[57]), .B2(n10583), .ZN(n8111) );
  ND2D1BWP30P140LVT U11895 ( .A1(n8112), .A2(n8111), .ZN(N4344) );
  AOI22D1BWP30P140LVT U11896 ( .A1(i_data_bus[94]), .A2(n10582), .B1(
        i_data_bus[30]), .B2(n10581), .ZN(n8114) );
  AOI22D1BWP30P140LVT U11897 ( .A1(i_data_bus[126]), .A2(n10584), .B1(
        i_data_bus[62]), .B2(n10583), .ZN(n8113) );
  ND2D1BWP30P140LVT U11898 ( .A1(n8114), .A2(n8113), .ZN(N4349) );
  AOI22D1BWP30P140LVT U11899 ( .A1(i_data_bus[77]), .A2(n10582), .B1(
        i_data_bus[13]), .B2(n10581), .ZN(n8116) );
  AOI22D1BWP30P140LVT U11900 ( .A1(i_data_bus[109]), .A2(n10584), .B1(
        i_data_bus[45]), .B2(n10583), .ZN(n8115) );
  ND2D1BWP30P140LVT U11901 ( .A1(n8116), .A2(n8115), .ZN(N4332) );
  AOI22D1BWP30P140LVT U11902 ( .A1(i_data_bus[27]), .A2(n10581), .B1(
        i_data_bus[91]), .B2(n10582), .ZN(n8118) );
  AOI22D1BWP30P140LVT U11903 ( .A1(i_data_bus[123]), .A2(n10584), .B1(
        i_data_bus[59]), .B2(n10583), .ZN(n8117) );
  ND2D1BWP30P140LVT U11904 ( .A1(n8118), .A2(n8117), .ZN(N4346) );
  AOI22D1BWP30P140LVT U11905 ( .A1(i_data_bus[695]), .A2(n10564), .B1(
        i_data_bus[759]), .B2(n10562), .ZN(n8120) );
  AOI22D1BWP30P140LVT U11906 ( .A1(i_data_bus[663]), .A2(n10563), .B1(
        i_data_bus[727]), .B2(n10561), .ZN(n8119) );
  ND2D1BWP30P140LVT U11907 ( .A1(n8120), .A2(n8119), .ZN(N5422) );
  AOI22D1BWP30P140LVT U11908 ( .A1(i_data_bus[156]), .A2(n10452), .B1(
        i_data_bus[220]), .B2(n10451), .ZN(n8122) );
  AOI22D1BWP30P140LVT U11909 ( .A1(i_data_bus[252]), .A2(n10449), .B1(
        i_data_bus[188]), .B2(n10450), .ZN(n8121) );
  ND2D1BWP30P140LVT U11910 ( .A1(n8122), .A2(n8121), .ZN(N12059) );
  AOI22D1BWP30P140LVT U11911 ( .A1(i_data_bus[653]), .A2(n10563), .B1(
        i_data_bus[685]), .B2(n10564), .ZN(n8124) );
  AOI22D1BWP30P140LVT U11912 ( .A1(i_data_bus[749]), .A2(n10562), .B1(
        i_data_bus[717]), .B2(n10561), .ZN(n8123) );
  ND2D1BWP30P140LVT U11913 ( .A1(n8124), .A2(n8123), .ZN(N5412) );
  AOI22D1BWP30P140LVT U11914 ( .A1(i_data_bus[223]), .A2(n10451), .B1(
        i_data_bus[255]), .B2(n10449), .ZN(n8126) );
  AOI22D1BWP30P140LVT U11915 ( .A1(i_data_bus[159]), .A2(n10452), .B1(
        i_data_bus[191]), .B2(n10450), .ZN(n8125) );
  ND2D1BWP30P140LVT U11916 ( .A1(n8126), .A2(n8125), .ZN(N12062) );
  AOI22D1BWP30P140LVT U11917 ( .A1(i_data_bus[253]), .A2(n10449), .B1(
        i_data_bus[157]), .B2(n10452), .ZN(n8128) );
  AOI22D1BWP30P140LVT U11918 ( .A1(i_data_bus[221]), .A2(n10451), .B1(
        i_data_bus[189]), .B2(n10450), .ZN(n8127) );
  ND2D1BWP30P140LVT U11919 ( .A1(n8128), .A2(n8127), .ZN(N12060) );
  AOI22D1BWP30P140LVT U11920 ( .A1(i_data_bus[141]), .A2(n10452), .B1(
        i_data_bus[237]), .B2(n10449), .ZN(n8130) );
  AOI22D1BWP30P140LVT U11921 ( .A1(i_data_bus[205]), .A2(n10451), .B1(
        i_data_bus[173]), .B2(n10450), .ZN(n8129) );
  ND2D1BWP30P140LVT U11922 ( .A1(n8130), .A2(n8129), .ZN(N12044) );
  AOI22D1BWP30P140LVT U11923 ( .A1(i_data_bus[229]), .A2(n10449), .B1(
        i_data_bus[197]), .B2(n10451), .ZN(n8132) );
  AOI22D1BWP30P140LVT U11924 ( .A1(i_data_bus[133]), .A2(n10452), .B1(
        i_data_bus[165]), .B2(n10450), .ZN(n8131) );
  ND2D1BWP30P140LVT U11925 ( .A1(n8132), .A2(n8131), .ZN(N12036) );
  AOI22D1BWP30P140LVT U11926 ( .A1(i_data_bus[248]), .A2(n10449), .B1(
        i_data_bus[152]), .B2(n10452), .ZN(n8134) );
  AOI22D1BWP30P140LVT U11927 ( .A1(i_data_bus[216]), .A2(n10451), .B1(
        i_data_bus[184]), .B2(n10450), .ZN(n8133) );
  ND2D1BWP30P140LVT U11928 ( .A1(n8134), .A2(n8133), .ZN(N12055) );
  AOI22D1BWP30P140LVT U11929 ( .A1(i_data_bus[698]), .A2(n10564), .B1(
        i_data_bus[762]), .B2(n10562), .ZN(n8136) );
  AOI22D1BWP30P140LVT U11930 ( .A1(i_data_bus[666]), .A2(n10563), .B1(
        i_data_bus[730]), .B2(n10561), .ZN(n8135) );
  ND2D1BWP30P140LVT U11931 ( .A1(n8136), .A2(n8135), .ZN(N5425) );
  AOI22D1BWP30P140LVT U11932 ( .A1(i_data_bus[673]), .A2(n10564), .B1(
        i_data_bus[641]), .B2(n10563), .ZN(n8138) );
  AOI22D1BWP30P140LVT U11933 ( .A1(i_data_bus[737]), .A2(n10562), .B1(
        i_data_bus[705]), .B2(n10561), .ZN(n8137) );
  ND2D1BWP30P140LVT U11934 ( .A1(n8138), .A2(n8137), .ZN(N5400) );
  AOI22D1BWP30P140LVT U11935 ( .A1(i_data_bus[746]), .A2(n10562), .B1(
        i_data_bus[682]), .B2(n10564), .ZN(n8140) );
  AOI22D1BWP30P140LVT U11936 ( .A1(i_data_bus[650]), .A2(n10563), .B1(
        i_data_bus[714]), .B2(n10561), .ZN(n8139) );
  ND2D1BWP30P140LVT U11937 ( .A1(n8140), .A2(n8139), .ZN(N5409) );
  AOI22D1BWP30P140LVT U11938 ( .A1(i_data_bus[665]), .A2(n10563), .B1(
        i_data_bus[761]), .B2(n10562), .ZN(n8142) );
  AOI22D1BWP30P140LVT U11939 ( .A1(i_data_bus[697]), .A2(n10564), .B1(
        i_data_bus[729]), .B2(n10561), .ZN(n8141) );
  ND2D1BWP30P140LVT U11940 ( .A1(n8142), .A2(n8141), .ZN(N5424) );
  AOI22D1BWP30P140LVT U11941 ( .A1(i_data_bus[208]), .A2(n10451), .B1(
        i_data_bus[240]), .B2(n10449), .ZN(n8144) );
  AOI22D1BWP30P140LVT U11942 ( .A1(i_data_bus[144]), .A2(n10452), .B1(
        i_data_bus[176]), .B2(n10450), .ZN(n8143) );
  ND2D1BWP30P140LVT U11943 ( .A1(n8144), .A2(n8143), .ZN(N12047) );
  AOI22D1BWP30P140LVT U11944 ( .A1(i_data_bus[733]), .A2(n10531), .B1(
        i_data_bus[765]), .B2(n10530), .ZN(n8146) );
  AOI22D1BWP30P140LVT U11945 ( .A1(i_data_bus[669]), .A2(n10529), .B1(
        i_data_bus[701]), .B2(n10532), .ZN(n8145) );
  ND2D1BWP30P140LVT U11946 ( .A1(n8146), .A2(n8145), .ZN(N7302) );
  AOI22D1BWP30P140LVT U11947 ( .A1(i_data_bus[658]), .A2(n10529), .B1(
        i_data_bus[754]), .B2(n10530), .ZN(n8148) );
  AOI22D1BWP30P140LVT U11948 ( .A1(i_data_bus[722]), .A2(n10531), .B1(
        i_data_bus[690]), .B2(n10532), .ZN(n8147) );
  ND2D1BWP30P140LVT U11949 ( .A1(n8148), .A2(n8147), .ZN(N7291) );
  AOI22D1BWP30P140LVT U11950 ( .A1(i_data_bus[650]), .A2(n10435), .B1(
        i_data_bus[714]), .B2(n10434), .ZN(n8150) );
  AOI22D1BWP30P140LVT U11951 ( .A1(i_data_bus[746]), .A2(n10433), .B1(
        i_data_bus[682]), .B2(n10436), .ZN(n8149) );
  ND2D1BWP30P140LVT U11952 ( .A1(n8150), .A2(n8149), .ZN(N12905) );
  AOI22D1BWP30P140LVT U11953 ( .A1(i_data_bus[707]), .A2(n10434), .B1(
        i_data_bus[739]), .B2(n10433), .ZN(n8152) );
  AOI22D1BWP30P140LVT U11954 ( .A1(i_data_bus[643]), .A2(n10435), .B1(
        i_data_bus[675]), .B2(n10436), .ZN(n8151) );
  ND2D1BWP30P140LVT U11955 ( .A1(n8152), .A2(n8151), .ZN(N12898) );
  AOI22D1BWP30P140LVT U11956 ( .A1(i_data_bus[665]), .A2(n10435), .B1(
        i_data_bus[729]), .B2(n10434), .ZN(n8154) );
  AOI22D1BWP30P140LVT U11957 ( .A1(i_data_bus[761]), .A2(n10433), .B1(
        i_data_bus[697]), .B2(n10436), .ZN(n8153) );
  ND2D1BWP30P140LVT U11958 ( .A1(n8154), .A2(n8153), .ZN(N12920) );
  AOI22D1BWP30P140LVT U11959 ( .A1(i_data_bus[652]), .A2(n10529), .B1(
        i_data_bus[748]), .B2(n10530), .ZN(n8156) );
  AOI22D1BWP30P140LVT U11960 ( .A1(i_data_bus[716]), .A2(n10531), .B1(
        i_data_bus[684]), .B2(n10532), .ZN(n8155) );
  ND2D1BWP30P140LVT U11961 ( .A1(n8156), .A2(n8155), .ZN(N7285) );
  AOI22D1BWP30P140LVT U11962 ( .A1(i_data_bus[733]), .A2(n10434), .B1(
        i_data_bus[765]), .B2(n10433), .ZN(n8158) );
  AOI22D1BWP30P140LVT U11963 ( .A1(i_data_bus[669]), .A2(n10435), .B1(
        i_data_bus[701]), .B2(n10436), .ZN(n8157) );
  ND2D1BWP30P140LVT U11964 ( .A1(n8158), .A2(n8157), .ZN(N12924) );
  AOI22D1BWP30P140LVT U11965 ( .A1(i_data_bus[766]), .A2(n10530), .B1(
        i_data_bus[670]), .B2(n10529), .ZN(n8160) );
  AOI22D1BWP30P140LVT U11966 ( .A1(i_data_bus[734]), .A2(n10531), .B1(
        i_data_bus[702]), .B2(n10532), .ZN(n8159) );
  ND2D1BWP30P140LVT U11967 ( .A1(n8160), .A2(n8159), .ZN(N7303) );
  AOI22D1BWP30P140LVT U11968 ( .A1(i_data_bus[715]), .A2(n10531), .B1(
        i_data_bus[651]), .B2(n10529), .ZN(n8162) );
  AOI22D1BWP30P140LVT U11969 ( .A1(i_data_bus[747]), .A2(n10530), .B1(
        i_data_bus[683]), .B2(n10532), .ZN(n8161) );
  ND2D1BWP30P140LVT U11970 ( .A1(n8162), .A2(n8161), .ZN(N7284) );
  AOI22D1BWP30P140LVT U11971 ( .A1(i_data_bus[722]), .A2(n10434), .B1(
        i_data_bus[754]), .B2(n10433), .ZN(n8164) );
  AOI22D1BWP30P140LVT U11972 ( .A1(i_data_bus[658]), .A2(n10435), .B1(
        i_data_bus[690]), .B2(n10436), .ZN(n8163) );
  ND2D1BWP30P140LVT U11973 ( .A1(n8164), .A2(n8163), .ZN(N12913) );
  AOI22D1BWP30P140LVT U11974 ( .A1(i_data_bus[665]), .A2(n10529), .B1(
        i_data_bus[729]), .B2(n10531), .ZN(n8166) );
  AOI22D1BWP30P140LVT U11975 ( .A1(i_data_bus[761]), .A2(n10530), .B1(
        i_data_bus[697]), .B2(n10532), .ZN(n8165) );
  ND2D1BWP30P140LVT U11976 ( .A1(n8166), .A2(n8165), .ZN(N7298) );
  AOI22D1BWP30P140LVT U11977 ( .A1(i_data_bus[757]), .A2(n10530), .B1(
        i_data_bus[661]), .B2(n10529), .ZN(n8168) );
  AOI22D1BWP30P140LVT U11978 ( .A1(i_data_bus[725]), .A2(n10531), .B1(
        i_data_bus[693]), .B2(n10532), .ZN(n8167) );
  ND2D1BWP30P140LVT U11979 ( .A1(n8168), .A2(n8167), .ZN(N7294) );
  AOI22D1BWP30P140LVT U11980 ( .A1(i_data_bus[746]), .A2(n10530), .B1(
        i_data_bus[650]), .B2(n10529), .ZN(n8170) );
  AOI22D1BWP30P140LVT U11981 ( .A1(i_data_bus[714]), .A2(n10531), .B1(
        i_data_bus[682]), .B2(n10532), .ZN(n8169) );
  ND2D1BWP30P140LVT U11982 ( .A1(n8170), .A2(n8169), .ZN(N7283) );
  AOI22D1BWP30P140LVT U11983 ( .A1(i_data_bus[659]), .A2(n10529), .B1(
        i_data_bus[723]), .B2(n10531), .ZN(n8172) );
  AOI22D1BWP30P140LVT U11984 ( .A1(i_data_bus[755]), .A2(n10530), .B1(
        i_data_bus[691]), .B2(n10532), .ZN(n8171) );
  ND2D1BWP30P140LVT U11985 ( .A1(n8172), .A2(n8171), .ZN(N7292) );
  AOI22D1BWP30P140LVT U11986 ( .A1(i_data_bus[706]), .A2(n10531), .B1(
        i_data_bus[738]), .B2(n10530), .ZN(n8174) );
  AOI22D1BWP30P140LVT U11987 ( .A1(i_data_bus[642]), .A2(n10529), .B1(
        i_data_bus[674]), .B2(n10532), .ZN(n8173) );
  ND2D1BWP30P140LVT U11988 ( .A1(n8174), .A2(n8173), .ZN(N7275) );
  AOI22D1BWP30P140LVT U11989 ( .A1(i_data_bus[752]), .A2(n10433), .B1(
        i_data_bus[656]), .B2(n10435), .ZN(n8176) );
  AOI22D1BWP30P140LVT U11990 ( .A1(i_data_bus[720]), .A2(n10434), .B1(
        i_data_bus[688]), .B2(n10436), .ZN(n8175) );
  ND2D1BWP30P140LVT U11991 ( .A1(n8176), .A2(n8175), .ZN(N12911) );
  AOI22D1BWP30P140LVT U11992 ( .A1(i_data_bus[642]), .A2(n10435), .B1(
        i_data_bus[738]), .B2(n10433), .ZN(n8178) );
  AOI22D1BWP30P140LVT U11993 ( .A1(i_data_bus[706]), .A2(n10434), .B1(
        i_data_bus[674]), .B2(n10436), .ZN(n8177) );
  ND2D1BWP30P140LVT U11994 ( .A1(n8178), .A2(n8177), .ZN(N12897) );
  AOI22D1BWP30P140LVT U11995 ( .A1(i_data_bus[652]), .A2(n10435), .B1(
        i_data_bus[748]), .B2(n10433), .ZN(n8180) );
  AOI22D1BWP30P140LVT U11996 ( .A1(i_data_bus[716]), .A2(n10434), .B1(
        i_data_bus[684]), .B2(n10436), .ZN(n8179) );
  ND2D1BWP30P140LVT U11997 ( .A1(n8180), .A2(n8179), .ZN(N12907) );
  AOI22D1BWP30P140LVT U11998 ( .A1(i_data_bus[446]), .A2(n10474), .B1(
        i_data_bus[510]), .B2(n10475), .ZN(n8182) );
  AOI22D1BWP30P140LVT U11999 ( .A1(i_data_bus[414]), .A2(n10473), .B1(
        i_data_bus[478]), .B2(n10476), .ZN(n8181) );
  ND2D1BWP30P140LVT U12000 ( .A1(n8182), .A2(n8181), .ZN(N10619) );
  AOI22D1BWP30P140LVT U12001 ( .A1(i_data_bus[418]), .A2(n10474), .B1(
        i_data_bus[386]), .B2(n10473), .ZN(n8184) );
  AOI22D1BWP30P140LVT U12002 ( .A1(i_data_bus[482]), .A2(n10475), .B1(
        i_data_bus[450]), .B2(n10476), .ZN(n8183) );
  ND2D1BWP30P140LVT U12003 ( .A1(n8184), .A2(n8183), .ZN(N10591) );
  AOI22D1BWP30P140LVT U12004 ( .A1(i_data_bus[443]), .A2(n10474), .B1(
        i_data_bus[507]), .B2(n10475), .ZN(n8186) );
  AOI22D1BWP30P140LVT U12005 ( .A1(i_data_bus[411]), .A2(n10473), .B1(
        i_data_bus[475]), .B2(n10476), .ZN(n8185) );
  ND2D1BWP30P140LVT U12006 ( .A1(n8186), .A2(n8185), .ZN(N10616) );
  AOI22D1BWP30P140LVT U12007 ( .A1(i_data_bus[417]), .A2(n10474), .B1(
        i_data_bus[481]), .B2(n10475), .ZN(n8188) );
  AOI22D1BWP30P140LVT U12008 ( .A1(i_data_bus[385]), .A2(n10473), .B1(
        i_data_bus[449]), .B2(n10476), .ZN(n8187) );
  ND2D1BWP30P140LVT U12009 ( .A1(n8188), .A2(n8187), .ZN(N10590) );
  AOI22D1BWP30P140LVT U12010 ( .A1(i_data_bus[498]), .A2(n10475), .B1(
        i_data_bus[434]), .B2(n10474), .ZN(n8190) );
  AOI22D1BWP30P140LVT U12011 ( .A1(i_data_bus[402]), .A2(n10473), .B1(
        i_data_bus[466]), .B2(n10476), .ZN(n8189) );
  ND2D1BWP30P140LVT U12012 ( .A1(n8190), .A2(n8189), .ZN(N10607) );
  AOI22D1BWP30P140LVT U12013 ( .A1(i_data_bus[430]), .A2(n10474), .B1(
        i_data_bus[494]), .B2(n10475), .ZN(n8192) );
  AOI22D1BWP30P140LVT U12014 ( .A1(i_data_bus[398]), .A2(n10473), .B1(
        i_data_bus[462]), .B2(n10476), .ZN(n8191) );
  ND2D1BWP30P140LVT U12015 ( .A1(n8192), .A2(n8191), .ZN(N10603) );
  AOI22D1BWP30P140LVT U12016 ( .A1(i_data_bus[392]), .A2(n10473), .B1(
        i_data_bus[424]), .B2(n10474), .ZN(n8194) );
  AOI22D1BWP30P140LVT U12017 ( .A1(i_data_bus[488]), .A2(n10475), .B1(
        i_data_bus[456]), .B2(n10476), .ZN(n8193) );
  ND2D1BWP30P140LVT U12018 ( .A1(n8194), .A2(n8193), .ZN(N10597) );
  AOI22D1BWP30P140LVT U12019 ( .A1(i_data_bus[406]), .A2(n10473), .B1(
        i_data_bus[438]), .B2(n10474), .ZN(n8196) );
  AOI22D1BWP30P140LVT U12020 ( .A1(i_data_bus[502]), .A2(n10475), .B1(
        i_data_bus[470]), .B2(n10476), .ZN(n8195) );
  ND2D1BWP30P140LVT U12021 ( .A1(n8196), .A2(n8195), .ZN(N10611) );
  AOI22D1BWP30P140LVT U12022 ( .A1(i_data_bus[49]), .A2(n10518), .B1(
        i_data_bus[17]), .B2(n10520), .ZN(n8198) );
  AOI22D1BWP30P140LVT U12023 ( .A1(i_data_bus[81]), .A2(n10517), .B1(
        i_data_bus[113]), .B2(n10519), .ZN(n8197) );
  ND2D1BWP30P140LVT U12024 ( .A1(n8198), .A2(n8197), .ZN(N8084) );
  AOI22D1BWP30P140LVT U12025 ( .A1(i_data_bus[43]), .A2(n10518), .B1(
        i_data_bus[11]), .B2(n10520), .ZN(n8200) );
  AOI22D1BWP30P140LVT U12026 ( .A1(i_data_bus[75]), .A2(n10517), .B1(
        i_data_bus[107]), .B2(n10519), .ZN(n8199) );
  ND2D1BWP30P140LVT U12027 ( .A1(n8200), .A2(n8199), .ZN(N8078) );
  AOI22D1BWP30P140LVT U12028 ( .A1(i_data_bus[92]), .A2(n10517), .B1(
        i_data_bus[28]), .B2(n10520), .ZN(n8202) );
  AOI22D1BWP30P140LVT U12029 ( .A1(i_data_bus[60]), .A2(n10518), .B1(
        i_data_bus[124]), .B2(n10519), .ZN(n8201) );
  ND2D1BWP30P140LVT U12030 ( .A1(n8202), .A2(n8201), .ZN(N8095) );
  AOI22D1BWP30P140LVT U12031 ( .A1(i_data_bus[80]), .A2(n10517), .B1(
        i_data_bus[16]), .B2(n10520), .ZN(n8204) );
  AOI22D1BWP30P140LVT U12032 ( .A1(i_data_bus[48]), .A2(n10518), .B1(
        i_data_bus[112]), .B2(n10519), .ZN(n8203) );
  ND2D1BWP30P140LVT U12033 ( .A1(n8204), .A2(n8203), .ZN(N8083) );
  AOI22D1BWP30P140LVT U12034 ( .A1(i_data_bus[87]), .A2(n10517), .B1(
        i_data_bus[55]), .B2(n10518), .ZN(n8206) );
  AOI22D1BWP30P140LVT U12035 ( .A1(i_data_bus[23]), .A2(n10520), .B1(
        i_data_bus[119]), .B2(n10519), .ZN(n8205) );
  ND2D1BWP30P140LVT U12036 ( .A1(n8206), .A2(n8205), .ZN(N8090) );
  AOI22D1BWP30P140LVT U12037 ( .A1(i_data_bus[46]), .A2(n10518), .B1(
        i_data_bus[78]), .B2(n10517), .ZN(n8208) );
  AOI22D1BWP30P140LVT U12038 ( .A1(i_data_bus[14]), .A2(n10520), .B1(
        i_data_bus[110]), .B2(n10519), .ZN(n8207) );
  ND2D1BWP30P140LVT U12039 ( .A1(n8208), .A2(n8207), .ZN(N8081) );
  AOI22D1BWP30P140LVT U12040 ( .A1(i_data_bus[611]), .A2(n10501), .B1(
        i_data_bus[579]), .B2(n10502), .ZN(n8210) );
  AOI22D1BWP30P140LVT U12041 ( .A1(i_data_bus[515]), .A2(n10503), .B1(
        i_data_bus[547]), .B2(n10504), .ZN(n8209) );
  ND2D1BWP30P140LVT U12042 ( .A1(n8210), .A2(n8209), .ZN(N8934) );
  AOI22D1BWP30P140LVT U12043 ( .A1(i_data_bus[631]), .A2(n10501), .B1(
        i_data_bus[535]), .B2(n10503), .ZN(n8212) );
  AOI22D1BWP30P140LVT U12044 ( .A1(i_data_bus[599]), .A2(n10502), .B1(
        i_data_bus[567]), .B2(n10504), .ZN(n8211) );
  ND2D1BWP30P140LVT U12045 ( .A1(n8212), .A2(n8211), .ZN(N8954) );
  AOI22D1BWP30P140LVT U12046 ( .A1(i_data_bus[605]), .A2(n10502), .B1(
        i_data_bus[541]), .B2(n10503), .ZN(n8214) );
  AOI22D1BWP30P140LVT U12047 ( .A1(i_data_bus[637]), .A2(n10501), .B1(
        i_data_bus[573]), .B2(n10504), .ZN(n8213) );
  ND2D1BWP30P140LVT U12048 ( .A1(n8214), .A2(n8213), .ZN(N8960) );
  AOI22D1BWP30P140LVT U12049 ( .A1(i_data_bus[533]), .A2(n10503), .B1(
        i_data_bus[629]), .B2(n10501), .ZN(n8216) );
  AOI22D1BWP30P140LVT U12050 ( .A1(i_data_bus[597]), .A2(n10502), .B1(
        i_data_bus[565]), .B2(n10504), .ZN(n8215) );
  ND2D1BWP30P140LVT U12051 ( .A1(n8216), .A2(n8215), .ZN(N8952) );
  AOI22D1BWP30P140LVT U12052 ( .A1(i_data_bus[608]), .A2(n10501), .B1(
        i_data_bus[576]), .B2(n10502), .ZN(n8218) );
  AOI22D1BWP30P140LVT U12053 ( .A1(i_data_bus[512]), .A2(n10503), .B1(
        i_data_bus[544]), .B2(n10504), .ZN(n8217) );
  ND2D1BWP30P140LVT U12054 ( .A1(n8218), .A2(n8217), .ZN(N8931) );
  AOI22D1BWP30P140LVT U12055 ( .A1(i_data_bus[9]), .A2(n10581), .B1(
        i_data_bus[41]), .B2(n10583), .ZN(n8220) );
  AOI22D1BWP30P140LVT U12056 ( .A1(i_data_bus[73]), .A2(n10582), .B1(
        i_data_bus[105]), .B2(n10584), .ZN(n8219) );
  ND2D1BWP30P140LVT U12057 ( .A1(n8220), .A2(n8219), .ZN(N4328) );
  AOI22D1BWP30P140LVT U12058 ( .A1(i_data_bus[17]), .A2(n10581), .B1(
        i_data_bus[81]), .B2(n10582), .ZN(n8222) );
  AOI22D1BWP30P140LVT U12059 ( .A1(i_data_bus[49]), .A2(n10583), .B1(
        i_data_bus[113]), .B2(n10584), .ZN(n8221) );
  ND2D1BWP30P140LVT U12060 ( .A1(n8222), .A2(n8221), .ZN(N4336) );
  AOI22D1BWP30P140LVT U12061 ( .A1(i_data_bus[51]), .A2(n10423), .B1(
        i_data_bus[19]), .B2(n10421), .ZN(n8224) );
  AOI22D1BWP30P140LVT U12062 ( .A1(i_data_bus[83]), .A2(n10422), .B1(
        i_data_bus[115]), .B2(n10424), .ZN(n8223) );
  ND2D1BWP30P140LVT U12063 ( .A1(n8224), .A2(n8223), .ZN(N13708) );
  AOI22D1BWP30P140LVT U12064 ( .A1(i_data_bus[455]), .A2(n10604), .B1(
        i_data_bus[391]), .B2(n10603), .ZN(n8226) );
  AOI22D1BWP30P140LVT U12065 ( .A1(i_data_bus[487]), .A2(n10602), .B1(
        i_data_bus[423]), .B2(n10601), .ZN(n8225) );
  ND2D1BWP30P140LVT U12066 ( .A1(n8226), .A2(n8225), .ZN(N3100) );
  AOI22D1BWP30P140LVT U12067 ( .A1(i_data_bus[69]), .A2(n10582), .B1(
        i_data_bus[5]), .B2(n10581), .ZN(n8228) );
  AOI22D1BWP30P140LVT U12068 ( .A1(i_data_bus[37]), .A2(n10583), .B1(
        i_data_bus[101]), .B2(n10584), .ZN(n8227) );
  ND2D1BWP30P140LVT U12069 ( .A1(n8228), .A2(n8227), .ZN(N4324) );
  AOI22D1BWP30P140LVT U12070 ( .A1(i_data_bus[87]), .A2(n10582), .B1(
        i_data_bus[55]), .B2(n10583), .ZN(n8230) );
  AOI22D1BWP30P140LVT U12071 ( .A1(i_data_bus[23]), .A2(n10581), .B1(
        i_data_bus[119]), .B2(n10584), .ZN(n8229) );
  ND2D1BWP30P140LVT U12072 ( .A1(n8230), .A2(n8229), .ZN(N4342) );
  AOI22D1BWP30P140LVT U12073 ( .A1(i_data_bus[499]), .A2(n10602), .B1(
        i_data_bus[403]), .B2(n10603), .ZN(n8232) );
  AOI22D1BWP30P140LVT U12074 ( .A1(i_data_bus[467]), .A2(n10604), .B1(
        i_data_bus[435]), .B2(n10601), .ZN(n8231) );
  ND2D1BWP30P140LVT U12075 ( .A1(n8232), .A2(n8231), .ZN(N3112) );
  AOI22D1BWP30P140LVT U12076 ( .A1(i_data_bus[67]), .A2(n10582), .B1(
        i_data_bus[3]), .B2(n10581), .ZN(n8234) );
  AOI22D1BWP30P140LVT U12077 ( .A1(i_data_bus[35]), .A2(n10583), .B1(
        i_data_bus[99]), .B2(n10584), .ZN(n8233) );
  ND2D1BWP30P140LVT U12078 ( .A1(n8234), .A2(n8233), .ZN(N4322) );
  AOI22D1BWP30P140LVT U12079 ( .A1(i_data_bus[462]), .A2(n10604), .B1(
        i_data_bus[494]), .B2(n10602), .ZN(n8236) );
  AOI22D1BWP30P140LVT U12080 ( .A1(i_data_bus[398]), .A2(n10603), .B1(
        i_data_bus[430]), .B2(n10601), .ZN(n8235) );
  ND2D1BWP30P140LVT U12081 ( .A1(n8236), .A2(n8235), .ZN(N3107) );
  AOI22D1BWP30P140LVT U12082 ( .A1(i_data_bus[10]), .A2(n10421), .B1(
        i_data_bus[42]), .B2(n10423), .ZN(n8238) );
  AOI22D1BWP30P140LVT U12083 ( .A1(i_data_bus[74]), .A2(n10422), .B1(
        i_data_bus[106]), .B2(n10424), .ZN(n8237) );
  ND2D1BWP30P140LVT U12084 ( .A1(n8238), .A2(n8237), .ZN(N13699) );
  AOI22D1BWP30P140LVT U12085 ( .A1(i_data_bus[38]), .A2(n10583), .B1(
        i_data_bus[6]), .B2(n10581), .ZN(n8240) );
  AOI22D1BWP30P140LVT U12086 ( .A1(i_data_bus[70]), .A2(n10582), .B1(
        i_data_bus[102]), .B2(n10584), .ZN(n8239) );
  ND2D1BWP30P140LVT U12087 ( .A1(n8240), .A2(n8239), .ZN(N4325) );
  AOI22D1BWP30P140LVT U12088 ( .A1(i_data_bus[93]), .A2(n10422), .B1(
        i_data_bus[29]), .B2(n10421), .ZN(n8242) );
  AOI22D1BWP30P140LVT U12089 ( .A1(i_data_bus[61]), .A2(n10423), .B1(
        i_data_bus[125]), .B2(n10424), .ZN(n8241) );
  ND2D1BWP30P140LVT U12090 ( .A1(n8242), .A2(n8241), .ZN(N13718) );
  AOI22D1BWP30P140LVT U12091 ( .A1(i_data_bus[409]), .A2(n10603), .B1(
        i_data_bus[505]), .B2(n10602), .ZN(n8244) );
  AOI22D1BWP30P140LVT U12092 ( .A1(i_data_bus[473]), .A2(n10604), .B1(
        i_data_bus[441]), .B2(n10601), .ZN(n8243) );
  ND2D1BWP30P140LVT U12093 ( .A1(n8244), .A2(n8243), .ZN(N3118) );
  AOI22D1BWP30P140LVT U12094 ( .A1(i_data_bus[39]), .A2(n10583), .B1(
        i_data_bus[7]), .B2(n10581), .ZN(n8246) );
  AOI22D1BWP30P140LVT U12095 ( .A1(i_data_bus[71]), .A2(n10582), .B1(
        i_data_bus[103]), .B2(n10584), .ZN(n8245) );
  ND2D1BWP30P140LVT U12096 ( .A1(n8246), .A2(n8245), .ZN(N4326) );
  AOI22D1BWP30P140LVT U12097 ( .A1(i_data_bus[0]), .A2(n10581), .B1(
        i_data_bus[64]), .B2(n10582), .ZN(n8248) );
  AOI22D1BWP30P140LVT U12098 ( .A1(i_data_bus[32]), .A2(n10583), .B1(
        i_data_bus[96]), .B2(n10584), .ZN(n8247) );
  ND2D1BWP30P140LVT U12099 ( .A1(n8248), .A2(n8247), .ZN(N4319) );
  AOI22D1BWP30P140LVT U12100 ( .A1(i_data_bus[38]), .A2(n10423), .B1(
        i_data_bus[6]), .B2(n10421), .ZN(n8250) );
  AOI22D1BWP30P140LVT U12101 ( .A1(i_data_bus[70]), .A2(n10422), .B1(
        i_data_bus[102]), .B2(n10424), .ZN(n8249) );
  ND2D1BWP30P140LVT U12102 ( .A1(n8250), .A2(n8249), .ZN(N13695) );
  AOI22D1BWP30P140LVT U12103 ( .A1(i_data_bus[392]), .A2(n10603), .B1(
        i_data_bus[456]), .B2(n10604), .ZN(n8252) );
  AOI22D1BWP30P140LVT U12104 ( .A1(i_data_bus[488]), .A2(n10602), .B1(
        i_data_bus[424]), .B2(n10601), .ZN(n8251) );
  ND2D1BWP30P140LVT U12105 ( .A1(n8252), .A2(n8251), .ZN(N3101) );
  AOI22D1BWP30P140LVT U12106 ( .A1(i_data_bus[74]), .A2(n10582), .B1(
        i_data_bus[42]), .B2(n10583), .ZN(n8254) );
  AOI22D1BWP30P140LVT U12107 ( .A1(i_data_bus[10]), .A2(n10581), .B1(
        i_data_bus[106]), .B2(n10584), .ZN(n8253) );
  ND2D1BWP30P140LVT U12108 ( .A1(n8254), .A2(n8253), .ZN(N4329) );
  AOI22D1BWP30P140LVT U12109 ( .A1(i_data_bus[65]), .A2(n10582), .B1(
        i_data_bus[1]), .B2(n10581), .ZN(n8256) );
  AOI22D1BWP30P140LVT U12110 ( .A1(i_data_bus[33]), .A2(n10583), .B1(
        i_data_bus[97]), .B2(n10584), .ZN(n8255) );
  ND2D1BWP30P140LVT U12111 ( .A1(n8256), .A2(n8255), .ZN(N4320) );
  AOI22D1BWP30P140LVT U12112 ( .A1(i_data_bus[0]), .A2(n10421), .B1(
        i_data_bus[64]), .B2(n10422), .ZN(n8258) );
  AOI22D1BWP30P140LVT U12113 ( .A1(i_data_bus[32]), .A2(n10423), .B1(
        i_data_bus[96]), .B2(n10424), .ZN(n8257) );
  ND2D1BWP30P140LVT U12114 ( .A1(n8258), .A2(n8257), .ZN(N13689) );
  AOI22D1BWP30P140LVT U12115 ( .A1(i_data_bus[827]), .A2(n10592), .B1(
        i_data_bus[891]), .B2(n10591), .ZN(n8260) );
  AOI22D1BWP30P140LVT U12116 ( .A1(i_data_bus[795]), .A2(n10589), .B1(
        i_data_bus[859]), .B2(n10590), .ZN(n8259) );
  ND2D1BWP30P140LVT U12117 ( .A1(n8260), .A2(n8259), .ZN(N3768) );
  AOI22D1BWP30P140LVT U12118 ( .A1(i_data_bus[829]), .A2(n10592), .B1(
        i_data_bus[797]), .B2(n10589), .ZN(n8262) );
  AOI22D1BWP30P140LVT U12119 ( .A1(i_data_bus[893]), .A2(n10591), .B1(
        i_data_bus[861]), .B2(n10590), .ZN(n8261) );
  ND2D1BWP30P140LVT U12120 ( .A1(n8262), .A2(n8261), .ZN(N3770) );
  AOI22D1BWP30P140LVT U12121 ( .A1(i_data_bus[870]), .A2(n10591), .B1(
        i_data_bus[774]), .B2(n10589), .ZN(n8264) );
  AOI22D1BWP30P140LVT U12122 ( .A1(i_data_bus[806]), .A2(n10592), .B1(
        i_data_bus[838]), .B2(n10590), .ZN(n8263) );
  ND2D1BWP30P140LVT U12123 ( .A1(n8264), .A2(n8263), .ZN(N3747) );
  AOI22D1BWP30P140LVT U12124 ( .A1(i_data_bus[818]), .A2(n10592), .B1(
        i_data_bus[786]), .B2(n10589), .ZN(n8266) );
  AOI22D1BWP30P140LVT U12125 ( .A1(i_data_bus[882]), .A2(n10591), .B1(
        i_data_bus[850]), .B2(n10590), .ZN(n8265) );
  ND2D1BWP30P140LVT U12126 ( .A1(n8266), .A2(n8265), .ZN(N3759) );
  AOI22D1BWP30P140LVT U12127 ( .A1(i_data_bus[787]), .A2(n10589), .B1(
        i_data_bus[819]), .B2(n10592), .ZN(n8268) );
  AOI22D1BWP30P140LVT U12128 ( .A1(i_data_bus[883]), .A2(n10591), .B1(
        i_data_bus[851]), .B2(n10590), .ZN(n8267) );
  ND2D1BWP30P140LVT U12129 ( .A1(n8268), .A2(n8267), .ZN(N3760) );
  AOI22D1BWP30P140LVT U12130 ( .A1(i_data_bus[810]), .A2(n10592), .B1(
        i_data_bus[874]), .B2(n10591), .ZN(n8270) );
  AOI22D1BWP30P140LVT U12131 ( .A1(i_data_bus[778]), .A2(n10589), .B1(
        i_data_bus[842]), .B2(n10590), .ZN(n8269) );
  ND2D1BWP30P140LVT U12132 ( .A1(n8270), .A2(n8269), .ZN(N3751) );
  AOI22D1BWP30P140LVT U12133 ( .A1(i_data_bus[850]), .A2(n10463), .B1(
        i_data_bus[818]), .B2(n10464), .ZN(n8272) );
  AOI22D1BWP30P140LVT U12134 ( .A1(i_data_bus[882]), .A2(n10461), .B1(
        i_data_bus[786]), .B2(n10462), .ZN(n8271) );
  ND2D1BWP30P140LVT U12135 ( .A1(n8272), .A2(n8271), .ZN(N11255) );
  AOI22D1BWP30P140LVT U12136 ( .A1(i_data_bus[878]), .A2(n10461), .B1(
        i_data_bus[846]), .B2(n10463), .ZN(n8274) );
  AOI22D1BWP30P140LVT U12137 ( .A1(i_data_bus[814]), .A2(n10464), .B1(
        i_data_bus[782]), .B2(n10462), .ZN(n8273) );
  ND2D1BWP30P140LVT U12138 ( .A1(n8274), .A2(n8273), .ZN(N11251) );
  AOI22D1BWP30P140LVT U12139 ( .A1(i_data_bus[862]), .A2(n10463), .B1(
        i_data_bus[830]), .B2(n10464), .ZN(n8276) );
  AOI22D1BWP30P140LVT U12140 ( .A1(i_data_bus[894]), .A2(n10461), .B1(
        i_data_bus[798]), .B2(n10462), .ZN(n8275) );
  ND2D1BWP30P140LVT U12141 ( .A1(n8276), .A2(n8275), .ZN(N11267) );
  AOI22D1BWP30P140LVT U12142 ( .A1(i_data_bus[856]), .A2(n10463), .B1(
        i_data_bus[824]), .B2(n10464), .ZN(n8278) );
  AOI22D1BWP30P140LVT U12143 ( .A1(i_data_bus[888]), .A2(n10461), .B1(
        i_data_bus[792]), .B2(n10462), .ZN(n8277) );
  ND2D1BWP30P140LVT U12144 ( .A1(n8278), .A2(n8277), .ZN(N11261) );
  AOI22D1BWP30P140LVT U12145 ( .A1(i_data_bus[819]), .A2(n10464), .B1(
        i_data_bus[851]), .B2(n10463), .ZN(n8280) );
  AOI22D1BWP30P140LVT U12146 ( .A1(i_data_bus[883]), .A2(n10461), .B1(
        i_data_bus[787]), .B2(n10462), .ZN(n8279) );
  ND2D1BWP30P140LVT U12147 ( .A1(n8280), .A2(n8279), .ZN(N11256) );
  AOI22D1BWP30P140LVT U12148 ( .A1(i_data_bus[863]), .A2(n10463), .B1(
        i_data_bus[831]), .B2(n10464), .ZN(n8282) );
  AOI22D1BWP30P140LVT U12149 ( .A1(i_data_bus[895]), .A2(n10461), .B1(
        i_data_bus[799]), .B2(n10462), .ZN(n8281) );
  ND2D1BWP30P140LVT U12150 ( .A1(n8282), .A2(n8281), .ZN(N11268) );
  AOI22D1BWP30P140LVT U12151 ( .A1(i_data_bus[849]), .A2(n10463), .B1(
        i_data_bus[817]), .B2(n10464), .ZN(n8284) );
  AOI22D1BWP30P140LVT U12152 ( .A1(i_data_bus[881]), .A2(n10461), .B1(
        i_data_bus[785]), .B2(n10462), .ZN(n8283) );
  ND2D1BWP30P140LVT U12153 ( .A1(n8284), .A2(n8283), .ZN(N11254) );
  AOI22D1BWP30P140LVT U12154 ( .A1(i_data_bus[893]), .A2(n10461), .B1(
        i_data_bus[861]), .B2(n10463), .ZN(n8286) );
  AOI22D1BWP30P140LVT U12155 ( .A1(i_data_bus[829]), .A2(n10464), .B1(
        i_data_bus[797]), .B2(n10462), .ZN(n8285) );
  ND2D1BWP30P140LVT U12156 ( .A1(n8286), .A2(n8285), .ZN(N11266) );
  AOI22D1BWP30P140LVT U12157 ( .A1(i_data_bus[305]), .A2(n10606), .B1(
        i_data_bus[273]), .B2(n10605), .ZN(n8288) );
  AOI22D1BWP30P140LVT U12158 ( .A1(i_data_bus[369]), .A2(n10608), .B1(
        i_data_bus[337]), .B2(n10607), .ZN(n8287) );
  ND2D1BWP30P140LVT U12159 ( .A1(n8288), .A2(n8287), .ZN(N2894) );
  AOI22D1BWP30P140LVT U12160 ( .A1(i_data_bus[281]), .A2(n10605), .B1(
        i_data_bus[377]), .B2(n10608), .ZN(n8290) );
  AOI22D1BWP30P140LVT U12161 ( .A1(i_data_bus[313]), .A2(n10606), .B1(
        i_data_bus[345]), .B2(n10607), .ZN(n8289) );
  ND2D1BWP30P140LVT U12162 ( .A1(n8290), .A2(n8289), .ZN(N2902) );
  AOI22D1BWP30P140LVT U12163 ( .A1(i_data_bus[268]), .A2(n10605), .B1(
        i_data_bus[300]), .B2(n10606), .ZN(n8292) );
  AOI22D1BWP30P140LVT U12164 ( .A1(i_data_bus[364]), .A2(n10608), .B1(
        i_data_bus[332]), .B2(n10607), .ZN(n8291) );
  ND2D1BWP30P140LVT U12165 ( .A1(n8292), .A2(n8291), .ZN(N2889) );
  AOI22D1BWP30P140LVT U12166 ( .A1(i_data_bus[376]), .A2(n10608), .B1(
        i_data_bus[312]), .B2(n10606), .ZN(n8294) );
  AOI22D1BWP30P140LVT U12167 ( .A1(i_data_bus[280]), .A2(n10605), .B1(
        i_data_bus[344]), .B2(n10607), .ZN(n8293) );
  ND2D1BWP30P140LVT U12168 ( .A1(n8294), .A2(n8293), .ZN(N2901) );
  AOI22D1BWP30P140LVT U12169 ( .A1(i_data_bus[270]), .A2(n10605), .B1(
        i_data_bus[302]), .B2(n10606), .ZN(n8296) );
  AOI22D1BWP30P140LVT U12170 ( .A1(i_data_bus[366]), .A2(n10608), .B1(
        i_data_bus[334]), .B2(n10607), .ZN(n8295) );
  ND2D1BWP30P140LVT U12171 ( .A1(n8296), .A2(n8295), .ZN(N2891) );
  AOI22D1BWP30P140LVT U12172 ( .A1(i_data_bus[267]), .A2(n10605), .B1(
        i_data_bus[363]), .B2(n10608), .ZN(n8298) );
  AOI22D1BWP30P140LVT U12173 ( .A1(i_data_bus[299]), .A2(n10606), .B1(
        i_data_bus[331]), .B2(n10607), .ZN(n8297) );
  ND2D1BWP30P140LVT U12174 ( .A1(n8298), .A2(n8297), .ZN(N2888) );
  AOI22D1BWP30P140LVT U12175 ( .A1(i_data_bus[288]), .A2(n10606), .B1(
        i_data_bus[256]), .B2(n10605), .ZN(n8300) );
  AOI22D1BWP30P140LVT U12176 ( .A1(i_data_bus[352]), .A2(n10608), .B1(
        i_data_bus[320]), .B2(n10607), .ZN(n8299) );
  ND2D1BWP30P140LVT U12177 ( .A1(n8300), .A2(n8299), .ZN(N2877) );
  AOI22D1BWP30P140LVT U12178 ( .A1(i_data_bus[816]), .A2(n10525), .B1(
        i_data_bus[880]), .B2(n10526), .ZN(n8302) );
  AOI22D1BWP30P140LVT U12179 ( .A1(i_data_bus[784]), .A2(n10528), .B1(
        i_data_bus[848]), .B2(n10527), .ZN(n8301) );
  ND2D1BWP30P140LVT U12180 ( .A1(n8302), .A2(n8301), .ZN(N7505) );
  AOI22D1BWP30P140LVT U12181 ( .A1(i_data_bus[781]), .A2(n10528), .B1(
        i_data_bus[877]), .B2(n10526), .ZN(n8304) );
  AOI22D1BWP30P140LVT U12182 ( .A1(i_data_bus[813]), .A2(n10525), .B1(
        i_data_bus[845]), .B2(n10527), .ZN(n8303) );
  ND2D1BWP30P140LVT U12183 ( .A1(n8304), .A2(n8303), .ZN(N7502) );
  AOI22D1BWP30P140LVT U12184 ( .A1(i_data_bus[822]), .A2(n10525), .B1(
        i_data_bus[790]), .B2(n10528), .ZN(n8306) );
  AOI22D1BWP30P140LVT U12185 ( .A1(i_data_bus[886]), .A2(n10526), .B1(
        i_data_bus[854]), .B2(n10527), .ZN(n8305) );
  ND2D1BWP30P140LVT U12186 ( .A1(n8306), .A2(n8305), .ZN(N7511) );
  AOI22D1BWP30P140LVT U12187 ( .A1(i_data_bus[785]), .A2(n10528), .B1(
        i_data_bus[817]), .B2(n10525), .ZN(n8308) );
  AOI22D1BWP30P140LVT U12188 ( .A1(i_data_bus[881]), .A2(n10526), .B1(
        i_data_bus[849]), .B2(n10527), .ZN(n8307) );
  ND2D1BWP30P140LVT U12189 ( .A1(n8308), .A2(n8307), .ZN(N7506) );
  AOI22D1BWP30P140LVT U12190 ( .A1(i_data_bus[820]), .A2(n10525), .B1(
        i_data_bus[884]), .B2(n10526), .ZN(n8310) );
  AOI22D1BWP30P140LVT U12191 ( .A1(i_data_bus[788]), .A2(n10528), .B1(
        i_data_bus[852]), .B2(n10527), .ZN(n8309) );
  ND2D1BWP30P140LVT U12192 ( .A1(n8310), .A2(n8309), .ZN(N7509) );
  AOI22D1BWP30P140LVT U12193 ( .A1(i_data_bus[805]), .A2(n10525), .B1(
        i_data_bus[869]), .B2(n10526), .ZN(n8312) );
  AOI22D1BWP30P140LVT U12194 ( .A1(i_data_bus[773]), .A2(n10528), .B1(
        i_data_bus[837]), .B2(n10527), .ZN(n8311) );
  ND2D1BWP30P140LVT U12195 ( .A1(n8312), .A2(n8311), .ZN(N7494) );
  AOI22D1BWP30P140LVT U12196 ( .A1(i_data_bus[827]), .A2(n10525), .B1(
        i_data_bus[795]), .B2(n10528), .ZN(n8314) );
  AOI22D1BWP30P140LVT U12197 ( .A1(i_data_bus[891]), .A2(n10526), .B1(
        i_data_bus[859]), .B2(n10527), .ZN(n8313) );
  ND2D1BWP30P140LVT U12198 ( .A1(n8314), .A2(n8313), .ZN(N7516) );
  AOI22D1BWP30P140LVT U12199 ( .A1(i_data_bus[879]), .A2(n10526), .B1(
        i_data_bus[815]), .B2(n10525), .ZN(n8316) );
  AOI22D1BWP30P140LVT U12200 ( .A1(i_data_bus[783]), .A2(n10528), .B1(
        i_data_bus[847]), .B2(n10527), .ZN(n8315) );
  ND2D1BWP30P140LVT U12201 ( .A1(n8316), .A2(n8315), .ZN(N7504) );
  AOI22D1BWP30P140LVT U12202 ( .A1(i_data_bus[807]), .A2(n10592), .B1(
        i_data_bus[839]), .B2(n10590), .ZN(n8318) );
  AOI22D1BWP30P140LVT U12203 ( .A1(i_data_bus[871]), .A2(n10591), .B1(
        i_data_bus[775]), .B2(n10589), .ZN(n8317) );
  ND2D1BWP30P140LVT U12204 ( .A1(n8318), .A2(n8317), .ZN(N3748) );
  AOI22D1BWP30P140LVT U12205 ( .A1(i_data_bus[866]), .A2(n10591), .B1(
        i_data_bus[802]), .B2(n10592), .ZN(n8320) );
  AOI22D1BWP30P140LVT U12206 ( .A1(i_data_bus[834]), .A2(n10590), .B1(
        i_data_bus[770]), .B2(n10589), .ZN(n8319) );
  ND2D1BWP30P140LVT U12207 ( .A1(n8320), .A2(n8319), .ZN(N3743) );
  AOI22D1BWP30P140LVT U12208 ( .A1(i_data_bus[886]), .A2(n10591), .B1(
        i_data_bus[854]), .B2(n10590), .ZN(n8322) );
  AOI22D1BWP30P140LVT U12209 ( .A1(i_data_bus[822]), .A2(n10592), .B1(
        i_data_bus[790]), .B2(n10589), .ZN(n8321) );
  ND2D1BWP30P140LVT U12210 ( .A1(n8322), .A2(n8321), .ZN(N3763) );
  AOI22D1BWP30P140LVT U12211 ( .A1(i_data_bus[836]), .A2(n10590), .B1(
        i_data_bus[804]), .B2(n10592), .ZN(n8324) );
  AOI22D1BWP30P140LVT U12212 ( .A1(i_data_bus[868]), .A2(n10591), .B1(
        i_data_bus[772]), .B2(n10589), .ZN(n8323) );
  ND2D1BWP30P140LVT U12213 ( .A1(n8324), .A2(n8323), .ZN(N3745) );
  AOI22D1BWP30P140LVT U12214 ( .A1(i_data_bus[881]), .A2(n10591), .B1(
        i_data_bus[817]), .B2(n10592), .ZN(n8326) );
  AOI22D1BWP30P140LVT U12215 ( .A1(i_data_bus[849]), .A2(n10590), .B1(
        i_data_bus[785]), .B2(n10589), .ZN(n8325) );
  ND2D1BWP30P140LVT U12216 ( .A1(n8326), .A2(n8325), .ZN(N3758) );
  AOI22D1BWP30P140LVT U12217 ( .A1(i_data_bus[856]), .A2(n10590), .B1(
        i_data_bus[824]), .B2(n10592), .ZN(n8328) );
  AOI22D1BWP30P140LVT U12218 ( .A1(i_data_bus[888]), .A2(n10591), .B1(
        i_data_bus[792]), .B2(n10589), .ZN(n8327) );
  ND2D1BWP30P140LVT U12219 ( .A1(n8328), .A2(n8327), .ZN(N3765) );
  AOI22D1BWP30P140LVT U12220 ( .A1(i_data_bus[869]), .A2(n10591), .B1(
        i_data_bus[837]), .B2(n10590), .ZN(n8330) );
  AOI22D1BWP30P140LVT U12221 ( .A1(i_data_bus[805]), .A2(n10592), .B1(
        i_data_bus[773]), .B2(n10589), .ZN(n8329) );
  ND2D1BWP30P140LVT U12222 ( .A1(n8330), .A2(n8329), .ZN(N3746) );
  AOI22D1BWP30P140LVT U12223 ( .A1(i_data_bus[814]), .A2(n10592), .B1(
        i_data_bus[846]), .B2(n10590), .ZN(n8332) );
  AOI22D1BWP30P140LVT U12224 ( .A1(i_data_bus[878]), .A2(n10591), .B1(
        i_data_bus[782]), .B2(n10589), .ZN(n8331) );
  ND2D1BWP30P140LVT U12225 ( .A1(n8332), .A2(n8331), .ZN(N3755) );
  AOI22D1BWP30P140LVT U12226 ( .A1(i_data_bus[855]), .A2(n10590), .B1(
        i_data_bus[887]), .B2(n10591), .ZN(n8334) );
  AOI22D1BWP30P140LVT U12227 ( .A1(i_data_bus[823]), .A2(n10592), .B1(
        i_data_bus[791]), .B2(n10589), .ZN(n8333) );
  ND2D1BWP30P140LVT U12228 ( .A1(n8334), .A2(n8333), .ZN(N3764) );
  AOI22D1BWP30P140LVT U12229 ( .A1(i_data_bus[189]), .A2(n10545), .B1(
        i_data_bus[157]), .B2(n10546), .ZN(n8336) );
  AOI22D1BWP30P140LVT U12230 ( .A1(i_data_bus[253]), .A2(n10547), .B1(
        i_data_bus[221]), .B2(n10548), .ZN(n8335) );
  ND2D1BWP30P140LVT U12231 ( .A1(n8336), .A2(n8335), .ZN(N6438) );
  AOI22D1BWP30P140LVT U12232 ( .A1(i_data_bus[161]), .A2(n10545), .B1(
        i_data_bus[225]), .B2(n10547), .ZN(n8338) );
  AOI22D1BWP30P140LVT U12233 ( .A1(i_data_bus[129]), .A2(n10546), .B1(
        i_data_bus[193]), .B2(n10548), .ZN(n8337) );
  ND2D1BWP30P140LVT U12234 ( .A1(n8338), .A2(n8337), .ZN(N6410) );
  AOI22D1BWP30P140LVT U12235 ( .A1(i_data_bus[163]), .A2(n10545), .B1(
        i_data_bus[131]), .B2(n10546), .ZN(n8340) );
  AOI22D1BWP30P140LVT U12236 ( .A1(i_data_bus[227]), .A2(n10547), .B1(
        i_data_bus[195]), .B2(n10548), .ZN(n8339) );
  ND2D1BWP30P140LVT U12237 ( .A1(n8340), .A2(n8339), .ZN(N6412) );
  AOI22D1BWP30P140LVT U12238 ( .A1(i_data_bus[128]), .A2(n10546), .B1(
        i_data_bus[160]), .B2(n10545), .ZN(n8342) );
  AOI22D1BWP30P140LVT U12239 ( .A1(i_data_bus[224]), .A2(n10547), .B1(
        i_data_bus[192]), .B2(n10548), .ZN(n8341) );
  ND2D1BWP30P140LVT U12240 ( .A1(n8342), .A2(n8341), .ZN(N6409) );
  AOI22D1BWP30P140LVT U12241 ( .A1(i_data_bus[179]), .A2(n10545), .B1(
        i_data_bus[243]), .B2(n10547), .ZN(n8344) );
  AOI22D1BWP30P140LVT U12242 ( .A1(i_data_bus[147]), .A2(n10546), .B1(
        i_data_bus[211]), .B2(n10548), .ZN(n8343) );
  ND2D1BWP30P140LVT U12243 ( .A1(n8344), .A2(n8343), .ZN(N6428) );
  AOI22D1BWP30P140LVT U12244 ( .A1(i_data_bus[148]), .A2(n10546), .B1(
        i_data_bus[244]), .B2(n10547), .ZN(n8346) );
  AOI22D1BWP30P140LVT U12245 ( .A1(i_data_bus[180]), .A2(n10545), .B1(
        i_data_bus[212]), .B2(n10548), .ZN(n8345) );
  ND2D1BWP30P140LVT U12246 ( .A1(n8346), .A2(n8345), .ZN(N6429) );
  AOI22D1BWP30P140LVT U12247 ( .A1(i_data_bus[184]), .A2(n10545), .B1(
        i_data_bus[152]), .B2(n10546), .ZN(n8348) );
  AOI22D1BWP30P140LVT U12248 ( .A1(i_data_bus[248]), .A2(n10547), .B1(
        i_data_bus[216]), .B2(n10548), .ZN(n8347) );
  ND2D1BWP30P140LVT U12249 ( .A1(n8348), .A2(n8347), .ZN(N6433) );
  AOI22D1BWP30P140LVT U12250 ( .A1(i_data_bus[155]), .A2(n10546), .B1(
        i_data_bus[251]), .B2(n10547), .ZN(n8350) );
  AOI22D1BWP30P140LVT U12251 ( .A1(i_data_bus[187]), .A2(n10545), .B1(
        i_data_bus[219]), .B2(n10548), .ZN(n8349) );
  ND2D1BWP30P140LVT U12252 ( .A1(n8350), .A2(n8349), .ZN(N6436) );
  AOI22D1BWP30P140LVT U12253 ( .A1(i_data_bus[270]), .A2(n10480), .B1(
        i_data_bus[366]), .B2(n10479), .ZN(n8352) );
  AOI22D1BWP30P140LVT U12254 ( .A1(i_data_bus[334]), .A2(n10478), .B1(
        i_data_bus[302]), .B2(n10477), .ZN(n8351) );
  ND2D1BWP30P140LVT U12255 ( .A1(n8352), .A2(n8351), .ZN(N10387) );
  AOI22D1BWP30P140LVT U12256 ( .A1(i_data_bus[266]), .A2(n10480), .B1(
        i_data_bus[362]), .B2(n10479), .ZN(n8354) );
  AOI22D1BWP30P140LVT U12257 ( .A1(i_data_bus[330]), .A2(n10478), .B1(
        i_data_bus[298]), .B2(n10477), .ZN(n8353) );
  ND2D1BWP30P140LVT U12258 ( .A1(n8354), .A2(n8353), .ZN(N10383) );
  AOI22D1BWP30P140LVT U12259 ( .A1(i_data_bus[945]), .A2(n10588), .B1(
        i_data_bus[977]), .B2(n10586), .ZN(n8356) );
  AOI22D1BWP30P140LVT U12260 ( .A1(i_data_bus[1009]), .A2(n10585), .B1(
        i_data_bus[913]), .B2(n10587), .ZN(n8355) );
  ND2D1BWP30P140LVT U12261 ( .A1(n8356), .A2(n8355), .ZN(N3974) );
  AOI22D1BWP30P140LVT U12262 ( .A1(i_data_bus[931]), .A2(n10588), .B1(
        i_data_bus[963]), .B2(n10586), .ZN(n8358) );
  AOI22D1BWP30P140LVT U12263 ( .A1(i_data_bus[995]), .A2(n10585), .B1(
        i_data_bus[899]), .B2(n10587), .ZN(n8357) );
  ND2D1BWP30P140LVT U12264 ( .A1(n8358), .A2(n8357), .ZN(N3960) );
  AOI22D1BWP30P140LVT U12265 ( .A1(i_data_bus[292]), .A2(n10477), .B1(
        i_data_bus[356]), .B2(n10479), .ZN(n8360) );
  AOI22D1BWP30P140LVT U12266 ( .A1(i_data_bus[324]), .A2(n10478), .B1(
        i_data_bus[260]), .B2(n10480), .ZN(n8359) );
  ND2D1BWP30P140LVT U12267 ( .A1(n8360), .A2(n8359), .ZN(N10377) );
  AOI22D1BWP30P140LVT U12268 ( .A1(i_data_bus[954]), .A2(n10588), .B1(
        i_data_bus[986]), .B2(n10586), .ZN(n8362) );
  AOI22D1BWP30P140LVT U12269 ( .A1(i_data_bus[1018]), .A2(n10585), .B1(
        i_data_bus[922]), .B2(n10587), .ZN(n8361) );
  ND2D1BWP30P140LVT U12270 ( .A1(n8362), .A2(n8361), .ZN(N3983) );
  AOI22D1BWP30P140LVT U12271 ( .A1(i_data_bus[309]), .A2(n10477), .B1(
        i_data_bus[373]), .B2(n10479), .ZN(n8364) );
  AOI22D1BWP30P140LVT U12272 ( .A1(i_data_bus[341]), .A2(n10478), .B1(
        i_data_bus[277]), .B2(n10480), .ZN(n8363) );
  ND2D1BWP30P140LVT U12273 ( .A1(n8364), .A2(n8363), .ZN(N10394) );
  AOI22D1BWP30P140LVT U12274 ( .A1(i_data_bus[947]), .A2(n10588), .B1(
        i_data_bus[1011]), .B2(n10585), .ZN(n8366) );
  AOI22D1BWP30P140LVT U12275 ( .A1(i_data_bus[979]), .A2(n10586), .B1(
        i_data_bus[915]), .B2(n10587), .ZN(n8365) );
  ND2D1BWP30P140LVT U12276 ( .A1(n8366), .A2(n8365), .ZN(N3976) );
  AOI22D1BWP30P140LVT U12277 ( .A1(i_data_bus[1005]), .A2(n10585), .B1(
        i_data_bus[941]), .B2(n10588), .ZN(n8368) );
  AOI22D1BWP30P140LVT U12278 ( .A1(i_data_bus[973]), .A2(n10586), .B1(
        i_data_bus[909]), .B2(n10587), .ZN(n8367) );
  ND2D1BWP30P140LVT U12279 ( .A1(n8368), .A2(n8367), .ZN(N3970) );
  AOI22D1BWP30P140LVT U12280 ( .A1(i_data_bus[968]), .A2(n10586), .B1(
        i_data_bus[1000]), .B2(n10585), .ZN(n8370) );
  AOI22D1BWP30P140LVT U12281 ( .A1(i_data_bus[936]), .A2(n10588), .B1(
        i_data_bus[904]), .B2(n10587), .ZN(n8369) );
  ND2D1BWP30P140LVT U12282 ( .A1(n8370), .A2(n8369), .ZN(N3965) );
  AOI22D1BWP30P140LVT U12283 ( .A1(i_data_bus[315]), .A2(n10477), .B1(
        i_data_bus[379]), .B2(n10479), .ZN(n8372) );
  AOI22D1BWP30P140LVT U12284 ( .A1(i_data_bus[347]), .A2(n10478), .B1(
        i_data_bus[283]), .B2(n10480), .ZN(n8371) );
  ND2D1BWP30P140LVT U12285 ( .A1(n8372), .A2(n8371), .ZN(N10400) );
  AOI22D1BWP30P140LVT U12286 ( .A1(i_data_bus[1013]), .A2(n10585), .B1(
        i_data_bus[949]), .B2(n10588), .ZN(n8374) );
  AOI22D1BWP30P140LVT U12287 ( .A1(i_data_bus[981]), .A2(n10586), .B1(
        i_data_bus[917]), .B2(n10587), .ZN(n8373) );
  ND2D1BWP30P140LVT U12288 ( .A1(n8374), .A2(n8373), .ZN(N3978) );
  AOI22D1BWP30P140LVT U12289 ( .A1(i_data_bus[965]), .A2(n10586), .B1(
        i_data_bus[997]), .B2(n10585), .ZN(n8376) );
  AOI22D1BWP30P140LVT U12290 ( .A1(i_data_bus[933]), .A2(n10588), .B1(
        i_data_bus[901]), .B2(n10587), .ZN(n8375) );
  ND2D1BWP30P140LVT U12291 ( .A1(n8376), .A2(n8375), .ZN(N3962) );
  AOI22D1BWP30P140LVT U12292 ( .A1(i_data_bus[275]), .A2(n10480), .B1(
        i_data_bus[371]), .B2(n10479), .ZN(n8378) );
  AOI22D1BWP30P140LVT U12293 ( .A1(i_data_bus[307]), .A2(n10477), .B1(
        i_data_bus[339]), .B2(n10478), .ZN(n8377) );
  ND2D1BWP30P140LVT U12294 ( .A1(n8378), .A2(n8377), .ZN(N10392) );
  AOI22D1BWP30P140LVT U12295 ( .A1(i_data_bus[314]), .A2(n10477), .B1(
        i_data_bus[378]), .B2(n10479), .ZN(n8380) );
  AOI22D1BWP30P140LVT U12296 ( .A1(i_data_bus[282]), .A2(n10480), .B1(
        i_data_bus[346]), .B2(n10478), .ZN(n8379) );
  ND2D1BWP30P140LVT U12297 ( .A1(n8380), .A2(n8379), .ZN(N10399) );
  AOI22D1BWP30P140LVT U12298 ( .A1(i_data_bus[273]), .A2(n10480), .B1(
        i_data_bus[369]), .B2(n10479), .ZN(n8382) );
  AOI22D1BWP30P140LVT U12299 ( .A1(i_data_bus[305]), .A2(n10477), .B1(
        i_data_bus[337]), .B2(n10478), .ZN(n8381) );
  ND2D1BWP30P140LVT U12300 ( .A1(n8382), .A2(n8381), .ZN(N10390) );
  AOI22D1BWP30P140LVT U12301 ( .A1(i_data_bus[460]), .A2(n10538), .B1(
        i_data_bus[492]), .B2(n10539), .ZN(n8384) );
  AOI22D1BWP30P140LVT U12302 ( .A1(i_data_bus[428]), .A2(n10540), .B1(
        i_data_bus[396]), .B2(n10537), .ZN(n8383) );
  ND2D1BWP30P140LVT U12303 ( .A1(n8384), .A2(n8383), .ZN(N6853) );
  AOI22D1BWP30P140LVT U12304 ( .A1(i_data_bus[483]), .A2(n10539), .B1(
        i_data_bus[419]), .B2(n10540), .ZN(n8386) );
  AOI22D1BWP30P140LVT U12305 ( .A1(i_data_bus[451]), .A2(n10538), .B1(
        i_data_bus[387]), .B2(n10537), .ZN(n8385) );
  ND2D1BWP30P140LVT U12306 ( .A1(n8386), .A2(n8385), .ZN(N6844) );
  AOI22D1BWP30P140LVT U12307 ( .A1(i_data_bus[496]), .A2(n10539), .B1(
        i_data_bus[432]), .B2(n10540), .ZN(n8388) );
  AOI22D1BWP30P140LVT U12308 ( .A1(i_data_bus[464]), .A2(n10538), .B1(
        i_data_bus[400]), .B2(n10537), .ZN(n8387) );
  ND2D1BWP30P140LVT U12309 ( .A1(n8388), .A2(n8387), .ZN(N6857) );
  AOI22D1BWP30P140LVT U12310 ( .A1(i_data_bus[310]), .A2(n10477), .B1(
        i_data_bus[374]), .B2(n10479), .ZN(n8390) );
  AOI22D1BWP30P140LVT U12311 ( .A1(i_data_bus[278]), .A2(n10480), .B1(
        i_data_bus[342]), .B2(n10478), .ZN(n8389) );
  ND2D1BWP30P140LVT U12312 ( .A1(n8390), .A2(n8389), .ZN(N10395) );
  AOI22D1BWP30P140LVT U12313 ( .A1(i_data_bus[280]), .A2(n10480), .B1(
        i_data_bus[376]), .B2(n10479), .ZN(n8392) );
  AOI22D1BWP30P140LVT U12314 ( .A1(i_data_bus[312]), .A2(n10477), .B1(
        i_data_bus[344]), .B2(n10478), .ZN(n8391) );
  ND2D1BWP30P140LVT U12315 ( .A1(n8392), .A2(n8391), .ZN(N10397) );
  AOI22D1BWP30P140LVT U12316 ( .A1(i_data_bus[505]), .A2(n10539), .B1(
        i_data_bus[441]), .B2(n10540), .ZN(n8394) );
  AOI22D1BWP30P140LVT U12317 ( .A1(i_data_bus[473]), .A2(n10538), .B1(
        i_data_bus[409]), .B2(n10537), .ZN(n8393) );
  ND2D1BWP30P140LVT U12318 ( .A1(n8394), .A2(n8393), .ZN(N6866) );
  AOI22D1BWP30P140LVT U12319 ( .A1(i_data_bus[471]), .A2(n10538), .B1(
        i_data_bus[503]), .B2(n10539), .ZN(n8396) );
  AOI22D1BWP30P140LVT U12320 ( .A1(i_data_bus[439]), .A2(n10540), .B1(
        i_data_bus[407]), .B2(n10537), .ZN(n8395) );
  ND2D1BWP30P140LVT U12321 ( .A1(n8396), .A2(n8395), .ZN(N6864) );
  AOI22D1BWP30P140LVT U12322 ( .A1(i_data_bus[467]), .A2(n10538), .B1(
        i_data_bus[435]), .B2(n10540), .ZN(n8398) );
  AOI22D1BWP30P140LVT U12323 ( .A1(i_data_bus[499]), .A2(n10539), .B1(
        i_data_bus[403]), .B2(n10537), .ZN(n8397) );
  ND2D1BWP30P140LVT U12324 ( .A1(n8398), .A2(n8397), .ZN(N6860) );
  AOI22D1BWP30P140LVT U12325 ( .A1(i_data_bus[447]), .A2(n10540), .B1(
        i_data_bus[511]), .B2(n10539), .ZN(n8400) );
  AOI22D1BWP30P140LVT U12326 ( .A1(i_data_bus[479]), .A2(n10538), .B1(
        i_data_bus[415]), .B2(n10537), .ZN(n8399) );
  ND2D1BWP30P140LVT U12327 ( .A1(n8400), .A2(n8399), .ZN(N6872) );
  AOI22D1BWP30P140LVT U12328 ( .A1(i_data_bus[281]), .A2(n10480), .B1(
        i_data_bus[377]), .B2(n10479), .ZN(n8402) );
  AOI22D1BWP30P140LVT U12329 ( .A1(i_data_bus[313]), .A2(n10477), .B1(
        i_data_bus[345]), .B2(n10478), .ZN(n8401) );
  ND2D1BWP30P140LVT U12330 ( .A1(n8402), .A2(n8401), .ZN(N10398) );
  AOI22D1BWP30P140LVT U12331 ( .A1(i_data_bus[684]), .A2(n10564), .B1(
        i_data_bus[652]), .B2(n10563), .ZN(n8404) );
  AOI22D1BWP30P140LVT U12332 ( .A1(i_data_bus[716]), .A2(n10561), .B1(
        i_data_bus[748]), .B2(n10562), .ZN(n8403) );
  ND2D1BWP30P140LVT U12333 ( .A1(n8404), .A2(n8403), .ZN(N5411) );
  AOI22D1BWP30P140LVT U12334 ( .A1(i_data_bus[728]), .A2(n10561), .B1(
        i_data_bus[696]), .B2(n10564), .ZN(n8406) );
  AOI22D1BWP30P140LVT U12335 ( .A1(i_data_bus[664]), .A2(n10563), .B1(
        i_data_bus[760]), .B2(n10562), .ZN(n8405) );
  ND2D1BWP30P140LVT U12336 ( .A1(n8406), .A2(n8405), .ZN(N5423) );
  AOI22D1BWP30P140LVT U12337 ( .A1(i_data_bus[719]), .A2(n10561), .B1(
        i_data_bus[655]), .B2(n10563), .ZN(n8408) );
  AOI22D1BWP30P140LVT U12338 ( .A1(i_data_bus[687]), .A2(n10564), .B1(
        i_data_bus[751]), .B2(n10562), .ZN(n8407) );
  ND2D1BWP30P140LVT U12339 ( .A1(n8408), .A2(n8407), .ZN(N5414) );
  AOI22D1BWP30P140LVT U12340 ( .A1(i_data_bus[713]), .A2(n10561), .B1(
        i_data_bus[649]), .B2(n10563), .ZN(n8410) );
  AOI22D1BWP30P140LVT U12341 ( .A1(i_data_bus[681]), .A2(n10564), .B1(
        i_data_bus[745]), .B2(n10562), .ZN(n8409) );
  ND2D1BWP30P140LVT U12342 ( .A1(n8410), .A2(n8409), .ZN(N5408) );
  AOI22D1BWP30P140LVT U12343 ( .A1(i_data_bus[699]), .A2(n10564), .B1(
        i_data_bus[731]), .B2(n10561), .ZN(n8412) );
  AOI22D1BWP30P140LVT U12344 ( .A1(i_data_bus[667]), .A2(n10563), .B1(
        i_data_bus[763]), .B2(n10562), .ZN(n8411) );
  ND2D1BWP30P140LVT U12345 ( .A1(n8412), .A2(n8411), .ZN(N5426) );
  AOI22D1BWP30P140LVT U12346 ( .A1(i_data_bus[707]), .A2(n10561), .B1(
        i_data_bus[675]), .B2(n10564), .ZN(n8414) );
  AOI22D1BWP30P140LVT U12347 ( .A1(i_data_bus[643]), .A2(n10563), .B1(
        i_data_bus[739]), .B2(n10562), .ZN(n8413) );
  ND2D1BWP30P140LVT U12348 ( .A1(n8414), .A2(n8413), .ZN(N5402) );
  AOI22D1BWP30P140LVT U12349 ( .A1(i_data_bus[691]), .A2(n10564), .B1(
        i_data_bus[723]), .B2(n10561), .ZN(n8416) );
  AOI22D1BWP30P140LVT U12350 ( .A1(i_data_bus[659]), .A2(n10563), .B1(
        i_data_bus[755]), .B2(n10562), .ZN(n8415) );
  ND2D1BWP30P140LVT U12351 ( .A1(n8416), .A2(n8415), .ZN(N5418) );
  AOI22D1BWP30P140LVT U12352 ( .A1(i_data_bus[692]), .A2(n10564), .B1(
        i_data_bus[724]), .B2(n10561), .ZN(n8418) );
  AOI22D1BWP30P140LVT U12353 ( .A1(i_data_bus[660]), .A2(n10563), .B1(
        i_data_bus[756]), .B2(n10562), .ZN(n8417) );
  ND2D1BWP30P140LVT U12354 ( .A1(n8418), .A2(n8417), .ZN(N5419) );
  AOI22D1BWP30P140LVT U12355 ( .A1(i_data_bus[706]), .A2(n10561), .B1(
        i_data_bus[642]), .B2(n10563), .ZN(n8420) );
  AOI22D1BWP30P140LVT U12356 ( .A1(i_data_bus[674]), .A2(n10564), .B1(
        i_data_bus[738]), .B2(n10562), .ZN(n8419) );
  ND2D1BWP30P140LVT U12357 ( .A1(n8420), .A2(n8419), .ZN(N5401) );
  AOI22D1BWP30P140LVT U12358 ( .A1(i_data_bus[119]), .A2(n10616), .B1(
        i_data_bus[55]), .B2(n10614), .ZN(n8422) );
  AOI22D1BWP30P140LVT U12359 ( .A1(i_data_bus[23]), .A2(n10615), .B1(
        i_data_bus[87]), .B2(n10613), .ZN(n8421) );
  ND2D1BWP30P140LVT U12360 ( .A1(n8422), .A2(n8421), .ZN(N2468) );
  AOI22D1BWP30P140LVT U12361 ( .A1(i_data_bus[4]), .A2(n10615), .B1(
        i_data_bus[36]), .B2(n10614), .ZN(n8424) );
  AOI22D1BWP30P140LVT U12362 ( .A1(i_data_bus[100]), .A2(n10616), .B1(
        i_data_bus[68]), .B2(n10613), .ZN(n8423) );
  ND2D1BWP30P140LVT U12363 ( .A1(n8424), .A2(n8423), .ZN(N2449) );
  AOI22D1BWP30P140LVT U12364 ( .A1(i_data_bus[38]), .A2(n10614), .B1(
        i_data_bus[102]), .B2(n10616), .ZN(n8426) );
  AOI22D1BWP30P140LVT U12365 ( .A1(i_data_bus[6]), .A2(n10615), .B1(
        i_data_bus[70]), .B2(n10613), .ZN(n8425) );
  ND2D1BWP30P140LVT U12366 ( .A1(n8426), .A2(n8425), .ZN(N2451) );
  AOI22D1BWP30P140LVT U12367 ( .A1(i_data_bus[60]), .A2(n10614), .B1(
        i_data_bus[28]), .B2(n10615), .ZN(n8428) );
  AOI22D1BWP30P140LVT U12368 ( .A1(i_data_bus[124]), .A2(n10616), .B1(
        i_data_bus[92]), .B2(n10613), .ZN(n8427) );
  ND2D1BWP30P140LVT U12369 ( .A1(n8428), .A2(n8427), .ZN(N2473) );
  AOI22D1BWP30P140LVT U12370 ( .A1(i_data_bus[120]), .A2(n10616), .B1(
        i_data_bus[56]), .B2(n10614), .ZN(n8430) );
  AOI22D1BWP30P140LVT U12371 ( .A1(i_data_bus[24]), .A2(n10615), .B1(
        i_data_bus[88]), .B2(n10613), .ZN(n8429) );
  ND2D1BWP30P140LVT U12372 ( .A1(n8430), .A2(n8429), .ZN(N2469) );
  AOI22D1BWP30P140LVT U12373 ( .A1(i_data_bus[771]), .A2(n10397), .B1(
        i_data_bus[803]), .B2(n10400), .ZN(n8432) );
  AOI22D1BWP30P140LVT U12374 ( .A1(i_data_bus[867]), .A2(n10398), .B1(
        i_data_bus[835]), .B2(n10399), .ZN(n8431) );
  ND2D1BWP30P140LVT U12375 ( .A1(n8432), .A2(n8431), .ZN(N14988) );
  AOI22D1BWP30P140LVT U12376 ( .A1(i_data_bus[805]), .A2(n10400), .B1(
        i_data_bus[869]), .B2(n10398), .ZN(n8434) );
  AOI22D1BWP30P140LVT U12377 ( .A1(i_data_bus[773]), .A2(n10397), .B1(
        i_data_bus[837]), .B2(n10399), .ZN(n8433) );
  ND2D1BWP30P140LVT U12378 ( .A1(n8434), .A2(n8433), .ZN(N14990) );
  AOI22D1BWP30P140LVT U12379 ( .A1(i_data_bus[893]), .A2(n10398), .B1(
        i_data_bus[797]), .B2(n10397), .ZN(n8436) );
  AOI22D1BWP30P140LVT U12380 ( .A1(i_data_bus[829]), .A2(n10400), .B1(
        i_data_bus[861]), .B2(n10399), .ZN(n8435) );
  ND2D1BWP30P140LVT U12381 ( .A1(n8436), .A2(n8435), .ZN(N15014) );
  AOI22D1BWP30P140LVT U12382 ( .A1(i_data_bus[885]), .A2(n10398), .B1(
        i_data_bus[821]), .B2(n10400), .ZN(n8438) );
  AOI22D1BWP30P140LVT U12383 ( .A1(i_data_bus[789]), .A2(n10397), .B1(
        i_data_bus[853]), .B2(n10399), .ZN(n8437) );
  ND2D1BWP30P140LVT U12384 ( .A1(n8438), .A2(n8437), .ZN(N15006) );
  AOI22D1BWP30P140LVT U12385 ( .A1(i_data_bus[780]), .A2(n10397), .B1(
        i_data_bus[876]), .B2(n10398), .ZN(n8440) );
  AOI22D1BWP30P140LVT U12386 ( .A1(i_data_bus[812]), .A2(n10400), .B1(
        i_data_bus[844]), .B2(n10399), .ZN(n8439) );
  ND2D1BWP30P140LVT U12387 ( .A1(n8440), .A2(n8439), .ZN(N14997) );
  AOI22D1BWP30P140LVT U12388 ( .A1(i_data_bus[883]), .A2(n10398), .B1(
        i_data_bus[787]), .B2(n10397), .ZN(n8442) );
  AOI22D1BWP30P140LVT U12389 ( .A1(i_data_bus[819]), .A2(n10400), .B1(
        i_data_bus[851]), .B2(n10399), .ZN(n8441) );
  ND2D1BWP30P140LVT U12390 ( .A1(n8442), .A2(n8441), .ZN(N15004) );
  AOI22D1BWP30P140LVT U12391 ( .A1(i_data_bus[322]), .A2(n10413), .B1(
        i_data_bus[354]), .B2(n10416), .ZN(n8444) );
  AOI22D1BWP30P140LVT U12392 ( .A1(i_data_bus[258]), .A2(n10415), .B1(
        i_data_bus[290]), .B2(n10414), .ZN(n8443) );
  ND2D1BWP30P140LVT U12393 ( .A1(n8444), .A2(n8443), .ZN(N14123) );
  AOI22D1BWP30P140LVT U12394 ( .A1(i_data_bus[270]), .A2(n10415), .B1(
        i_data_bus[366]), .B2(n10416), .ZN(n8446) );
  AOI22D1BWP30P140LVT U12395 ( .A1(i_data_bus[334]), .A2(n10413), .B1(
        i_data_bus[302]), .B2(n10414), .ZN(n8445) );
  ND2D1BWP30P140LVT U12396 ( .A1(n8446), .A2(n8445), .ZN(N14135) );
  AOI22D1BWP30P140LVT U12397 ( .A1(i_data_bus[271]), .A2(n10415), .B1(
        i_data_bus[367]), .B2(n10416), .ZN(n8448) );
  AOI22D1BWP30P140LVT U12398 ( .A1(i_data_bus[303]), .A2(n10414), .B1(
        i_data_bus[335]), .B2(n10413), .ZN(n8447) );
  ND2D1BWP30P140LVT U12399 ( .A1(n8448), .A2(n8447), .ZN(N14136) );
  AOI22D1BWP30P140LVT U12400 ( .A1(i_data_bus[314]), .A2(n10414), .B1(
        i_data_bus[378]), .B2(n10416), .ZN(n8450) );
  AOI22D1BWP30P140LVT U12401 ( .A1(i_data_bus[282]), .A2(n10415), .B1(
        i_data_bus[346]), .B2(n10413), .ZN(n8449) );
  ND2D1BWP30P140LVT U12402 ( .A1(n8450), .A2(n8449), .ZN(N14147) );
  AOI22D1BWP30P140LVT U12403 ( .A1(i_data_bus[328]), .A2(n10413), .B1(
        i_data_bus[360]), .B2(n10416), .ZN(n8452) );
  AOI22D1BWP30P140LVT U12404 ( .A1(i_data_bus[296]), .A2(n10414), .B1(
        i_data_bus[264]), .B2(n10415), .ZN(n8451) );
  ND2D1BWP30P140LVT U12405 ( .A1(n8452), .A2(n8451), .ZN(N14129) );
  AOI22D1BWP30P140LVT U12406 ( .A1(i_data_bus[267]), .A2(n10415), .B1(
        i_data_bus[363]), .B2(n10416), .ZN(n8454) );
  AOI22D1BWP30P140LVT U12407 ( .A1(i_data_bus[299]), .A2(n10414), .B1(
        i_data_bus[331]), .B2(n10413), .ZN(n8453) );
  ND2D1BWP30P140LVT U12408 ( .A1(n8454), .A2(n8453), .ZN(N14132) );
  AOI22D1BWP30P140LVT U12409 ( .A1(i_data_bus[349]), .A2(n10413), .B1(
        i_data_bus[381]), .B2(n10416), .ZN(n8456) );
  AOI22D1BWP30P140LVT U12410 ( .A1(i_data_bus[317]), .A2(n10414), .B1(
        i_data_bus[285]), .B2(n10415), .ZN(n8455) );
  ND2D1BWP30P140LVT U12411 ( .A1(n8456), .A2(n8455), .ZN(N14150) );
  AOI22D1BWP30P140LVT U12412 ( .A1(i_data_bus[260]), .A2(n10415), .B1(
        i_data_bus[356]), .B2(n10416), .ZN(n8458) );
  AOI22D1BWP30P140LVT U12413 ( .A1(i_data_bus[292]), .A2(n10414), .B1(
        i_data_bus[324]), .B2(n10413), .ZN(n8457) );
  ND2D1BWP30P140LVT U12414 ( .A1(n8458), .A2(n8457), .ZN(N14125) );
  AOI22D1BWP30P140LVT U12415 ( .A1(i_data_bus[862]), .A2(n10495), .B1(
        i_data_bus[830]), .B2(n10496), .ZN(n8460) );
  AOI22D1BWP30P140LVT U12416 ( .A1(i_data_bus[894]), .A2(n10494), .B1(
        i_data_bus[798]), .B2(n10493), .ZN(n8459) );
  ND2D1BWP30P140LVT U12417 ( .A1(n8460), .A2(n8459), .ZN(N9393) );
  AOI22D1BWP30P140LVT U12418 ( .A1(i_data_bus[882]), .A2(n10494), .B1(
        i_data_bus[850]), .B2(n10495), .ZN(n8462) );
  AOI22D1BWP30P140LVT U12419 ( .A1(i_data_bus[818]), .A2(n10496), .B1(
        i_data_bus[786]), .B2(n10493), .ZN(n8461) );
  ND2D1BWP30P140LVT U12420 ( .A1(n8462), .A2(n8461), .ZN(N9381) );
  AOI22D1BWP30P140LVT U12421 ( .A1(i_data_bus[870]), .A2(n10494), .B1(
        i_data_bus[838]), .B2(n10495), .ZN(n8464) );
  AOI22D1BWP30P140LVT U12422 ( .A1(i_data_bus[806]), .A2(n10496), .B1(
        i_data_bus[774]), .B2(n10493), .ZN(n8463) );
  ND2D1BWP30P140LVT U12423 ( .A1(n8464), .A2(n8463), .ZN(N9369) );
  AOI22D1BWP30P140LVT U12424 ( .A1(i_data_bus[887]), .A2(n10494), .B1(
        i_data_bus[823]), .B2(n10496), .ZN(n8466) );
  AOI22D1BWP30P140LVT U12425 ( .A1(i_data_bus[855]), .A2(n10495), .B1(
        i_data_bus[791]), .B2(n10493), .ZN(n8465) );
  ND2D1BWP30P140LVT U12426 ( .A1(n8466), .A2(n8465), .ZN(N9386) );
  AOI22D1BWP30P140LVT U12427 ( .A1(i_data_bus[857]), .A2(n10495), .B1(
        i_data_bus[825]), .B2(n10496), .ZN(n8468) );
  AOI22D1BWP30P140LVT U12428 ( .A1(i_data_bus[889]), .A2(n10494), .B1(
        i_data_bus[793]), .B2(n10493), .ZN(n8467) );
  ND2D1BWP30P140LVT U12429 ( .A1(n8468), .A2(n8467), .ZN(N9388) );
  AOI22D1BWP30P140LVT U12430 ( .A1(i_data_bus[849]), .A2(n10495), .B1(
        i_data_bus[817]), .B2(n10496), .ZN(n8470) );
  AOI22D1BWP30P140LVT U12431 ( .A1(i_data_bus[881]), .A2(n10494), .B1(
        i_data_bus[785]), .B2(n10493), .ZN(n8469) );
  ND2D1BWP30P140LVT U12432 ( .A1(n8470), .A2(n8469), .ZN(N9380) );
  AOI22D1BWP30P140LVT U12433 ( .A1(i_data_bus[895]), .A2(n10494), .B1(
        i_data_bus[831]), .B2(n10496), .ZN(n8472) );
  AOI22D1BWP30P140LVT U12434 ( .A1(i_data_bus[863]), .A2(n10495), .B1(
        i_data_bus[799]), .B2(n10493), .ZN(n8471) );
  ND2D1BWP30P140LVT U12435 ( .A1(n8472), .A2(n8471), .ZN(N9394) );
  AOI22D1BWP30P140LVT U12436 ( .A1(i_data_bus[840]), .A2(n10495), .B1(
        i_data_bus[808]), .B2(n10496), .ZN(n8474) );
  AOI22D1BWP30P140LVT U12437 ( .A1(i_data_bus[872]), .A2(n10494), .B1(
        i_data_bus[776]), .B2(n10493), .ZN(n8473) );
  ND2D1BWP30P140LVT U12438 ( .A1(n8474), .A2(n8473), .ZN(N9371) );
  AOI22D1BWP30P140LVT U12439 ( .A1(i_data_bus[836]), .A2(n10495), .B1(
        i_data_bus[804]), .B2(n10496), .ZN(n8476) );
  AOI22D1BWP30P140LVT U12440 ( .A1(i_data_bus[868]), .A2(n10494), .B1(
        i_data_bus[772]), .B2(n10493), .ZN(n8475) );
  ND2D1BWP30P140LVT U12441 ( .A1(n8476), .A2(n8475), .ZN(N9367) );
  AOI22D1BWP30P140LVT U12442 ( .A1(i_data_bus[996]), .A2(n10489), .B1(
        i_data_bus[964]), .B2(n10490), .ZN(n8478) );
  AOI22D1BWP30P140LVT U12443 ( .A1(i_data_bus[932]), .A2(n10491), .B1(
        i_data_bus[900]), .B2(n10492), .ZN(n8477) );
  ND2D1BWP30P140LVT U12444 ( .A1(n8478), .A2(n8477), .ZN(N9583) );
  AOI22D1BWP30P140LVT U12445 ( .A1(i_data_bus[993]), .A2(n10489), .B1(
        i_data_bus[961]), .B2(n10490), .ZN(n8480) );
  AOI22D1BWP30P140LVT U12446 ( .A1(i_data_bus[929]), .A2(n10491), .B1(
        i_data_bus[897]), .B2(n10492), .ZN(n8479) );
  ND2D1BWP30P140LVT U12447 ( .A1(n8480), .A2(n8479), .ZN(N9580) );
  AOI22D1BWP30P140LVT U12448 ( .A1(i_data_bus[946]), .A2(n10491), .B1(
        i_data_bus[1010]), .B2(n10489), .ZN(n8482) );
  AOI22D1BWP30P140LVT U12449 ( .A1(i_data_bus[978]), .A2(n10490), .B1(
        i_data_bus[914]), .B2(n10492), .ZN(n8481) );
  ND2D1BWP30P140LVT U12450 ( .A1(n8482), .A2(n8481), .ZN(N9597) );
  AOI22D1BWP30P140LVT U12451 ( .A1(i_data_bus[938]), .A2(n10491), .B1(
        i_data_bus[1002]), .B2(n10489), .ZN(n8484) );
  AOI22D1BWP30P140LVT U12452 ( .A1(i_data_bus[970]), .A2(n10490), .B1(
        i_data_bus[906]), .B2(n10492), .ZN(n8483) );
  ND2D1BWP30P140LVT U12453 ( .A1(n8484), .A2(n8483), .ZN(N9589) );
  AOI22D1BWP30P140LVT U12454 ( .A1(i_data_bus[1011]), .A2(n10489), .B1(
        i_data_bus[979]), .B2(n10490), .ZN(n8486) );
  AOI22D1BWP30P140LVT U12455 ( .A1(i_data_bus[947]), .A2(n10491), .B1(
        i_data_bus[915]), .B2(n10492), .ZN(n8485) );
  ND2D1BWP30P140LVT U12456 ( .A1(n8486), .A2(n8485), .ZN(N9598) );
  AOI22D1BWP30P140LVT U12457 ( .A1(i_data_bus[965]), .A2(n10490), .B1(
        i_data_bus[997]), .B2(n10489), .ZN(n8488) );
  AOI22D1BWP30P140LVT U12458 ( .A1(i_data_bus[933]), .A2(n10491), .B1(
        i_data_bus[901]), .B2(n10492), .ZN(n8487) );
  ND2D1BWP30P140LVT U12459 ( .A1(n8488), .A2(n8487), .ZN(N9584) );
  AOI22D1BWP30P140LVT U12460 ( .A1(i_data_bus[939]), .A2(n10491), .B1(
        i_data_bus[971]), .B2(n10490), .ZN(n8490) );
  AOI22D1BWP30P140LVT U12461 ( .A1(i_data_bus[1003]), .A2(n10489), .B1(
        i_data_bus[907]), .B2(n10492), .ZN(n8489) );
  ND2D1BWP30P140LVT U12462 ( .A1(n8490), .A2(n8489), .ZN(N9590) );
  AOI22D1BWP30P140LVT U12463 ( .A1(i_data_bus[706]), .A2(n10594), .B1(
        i_data_bus[642]), .B2(n10596), .ZN(n8492) );
  AOI22D1BWP30P140LVT U12464 ( .A1(i_data_bus[674]), .A2(n10593), .B1(
        i_data_bus[738]), .B2(n10595), .ZN(n8491) );
  ND2D1BWP30P140LVT U12465 ( .A1(n8492), .A2(n8491), .ZN(N3527) );
  AOI22D1BWP30P140LVT U12466 ( .A1(i_data_bus[710]), .A2(n10594), .B1(
        i_data_bus[678]), .B2(n10593), .ZN(n8494) );
  AOI22D1BWP30P140LVT U12467 ( .A1(i_data_bus[646]), .A2(n10596), .B1(
        i_data_bus[742]), .B2(n10595), .ZN(n8493) );
  ND2D1BWP30P140LVT U12468 ( .A1(n8494), .A2(n8493), .ZN(N3531) );
  AOI22D1BWP30P140LVT U12469 ( .A1(i_data_bus[686]), .A2(n10593), .B1(
        i_data_bus[654]), .B2(n10596), .ZN(n8496) );
  AOI22D1BWP30P140LVT U12470 ( .A1(i_data_bus[718]), .A2(n10594), .B1(
        i_data_bus[750]), .B2(n10595), .ZN(n8495) );
  ND2D1BWP30P140LVT U12471 ( .A1(n8496), .A2(n8495), .ZN(N3539) );
  AOI22D1BWP30P140LVT U12472 ( .A1(i_data_bus[695]), .A2(n10593), .B1(
        i_data_bus[727]), .B2(n10594), .ZN(n8498) );
  AOI22D1BWP30P140LVT U12473 ( .A1(i_data_bus[663]), .A2(n10596), .B1(
        i_data_bus[759]), .B2(n10595), .ZN(n8497) );
  ND2D1BWP30P140LVT U12474 ( .A1(n8498), .A2(n8497), .ZN(N3548) );
  AOI22D1BWP30P140LVT U12475 ( .A1(i_data_bus[709]), .A2(n10594), .B1(
        i_data_bus[677]), .B2(n10593), .ZN(n8500) );
  AOI22D1BWP30P140LVT U12476 ( .A1(i_data_bus[645]), .A2(n10596), .B1(
        i_data_bus[741]), .B2(n10595), .ZN(n8499) );
  ND2D1BWP30P140LVT U12477 ( .A1(n8500), .A2(n8499), .ZN(N3530) );
  AOI22D1BWP30P140LVT U12478 ( .A1(i_data_bus[673]), .A2(n10593), .B1(
        i_data_bus[705]), .B2(n10594), .ZN(n8502) );
  AOI22D1BWP30P140LVT U12479 ( .A1(i_data_bus[641]), .A2(n10596), .B1(
        i_data_bus[737]), .B2(n10595), .ZN(n8501) );
  ND2D1BWP30P140LVT U12480 ( .A1(n8502), .A2(n8501), .ZN(N3526) );
  AOI22D1BWP30P140LVT U12481 ( .A1(i_data_bus[672]), .A2(n10593), .B1(
        i_data_bus[704]), .B2(n10594), .ZN(n8504) );
  AOI22D1BWP30P140LVT U12482 ( .A1(i_data_bus[640]), .A2(n10596), .B1(
        i_data_bus[736]), .B2(n10595), .ZN(n8503) );
  ND2D1BWP30P140LVT U12483 ( .A1(n8504), .A2(n8503), .ZN(N3525) );
  AOI22D1BWP30P140LVT U12484 ( .A1(i_data_bus[728]), .A2(n10594), .B1(
        i_data_bus[696]), .B2(n10593), .ZN(n8506) );
  AOI22D1BWP30P140LVT U12485 ( .A1(i_data_bus[664]), .A2(n10596), .B1(
        i_data_bus[760]), .B2(n10595), .ZN(n8505) );
  ND2D1BWP30P140LVT U12486 ( .A1(n8506), .A2(n8505), .ZN(N3549) );
  AOI22D1BWP30P140LVT U12487 ( .A1(i_data_bus[702]), .A2(n10593), .B1(
        i_data_bus[670]), .B2(n10596), .ZN(n8508) );
  AOI22D1BWP30P140LVT U12488 ( .A1(i_data_bus[734]), .A2(n10594), .B1(
        i_data_bus[766]), .B2(n10595), .ZN(n8507) );
  ND2D1BWP30P140LVT U12489 ( .A1(n8508), .A2(n8507), .ZN(N3555) );
  AOI22D1BWP30P140LVT U12490 ( .A1(i_data_bus[711]), .A2(n10594), .B1(
        i_data_bus[647]), .B2(n10596), .ZN(n8510) );
  AOI22D1BWP30P140LVT U12491 ( .A1(i_data_bus[679]), .A2(n10593), .B1(
        i_data_bus[743]), .B2(n10595), .ZN(n8509) );
  ND2D1BWP30P140LVT U12492 ( .A1(n8510), .A2(n8509), .ZN(N3532) );
  AOI22D1BWP30P140LVT U12493 ( .A1(i_data_bus[693]), .A2(n10593), .B1(
        i_data_bus[661]), .B2(n10596), .ZN(n8512) );
  AOI22D1BWP30P140LVT U12494 ( .A1(i_data_bus[725]), .A2(n10594), .B1(
        i_data_bus[757]), .B2(n10595), .ZN(n8511) );
  ND2D1BWP30P140LVT U12495 ( .A1(n8512), .A2(n8511), .ZN(N3546) );
  AOI22D1BWP30P140LVT U12496 ( .A1(i_data_bus[692]), .A2(n10593), .B1(
        i_data_bus[724]), .B2(n10594), .ZN(n8514) );
  AOI22D1BWP30P140LVT U12497 ( .A1(i_data_bus[660]), .A2(n10596), .B1(
        i_data_bus[756]), .B2(n10595), .ZN(n8513) );
  ND2D1BWP30P140LVT U12498 ( .A1(n8514), .A2(n8513), .ZN(N3545) );
  AOI22D1BWP30P140LVT U12499 ( .A1(i_data_bus[485]), .A2(n10412), .B1(
        i_data_bus[453]), .B2(n10410), .ZN(n8516) );
  AOI22D1BWP30P140LVT U12500 ( .A1(i_data_bus[389]), .A2(n10409), .B1(
        i_data_bus[421]), .B2(n10411), .ZN(n8515) );
  ND2D1BWP30P140LVT U12501 ( .A1(n8516), .A2(n8515), .ZN(N14342) );
  AOI22D1BWP30P140LVT U12502 ( .A1(i_data_bus[469]), .A2(n10410), .B1(
        i_data_bus[501]), .B2(n10412), .ZN(n8518) );
  AOI22D1BWP30P140LVT U12503 ( .A1(i_data_bus[405]), .A2(n10409), .B1(
        i_data_bus[437]), .B2(n10411), .ZN(n8517) );
  ND2D1BWP30P140LVT U12504 ( .A1(n8518), .A2(n8517), .ZN(N14358) );
  AOI22D1BWP30P140LVT U12505 ( .A1(i_data_bus[457]), .A2(n10410), .B1(
        i_data_bus[393]), .B2(n10409), .ZN(n8520) );
  AOI22D1BWP30P140LVT U12506 ( .A1(i_data_bus[489]), .A2(n10412), .B1(
        i_data_bus[425]), .B2(n10411), .ZN(n8519) );
  ND2D1BWP30P140LVT U12507 ( .A1(n8520), .A2(n8519), .ZN(N14346) );
  AOI22D1BWP30P140LVT U12508 ( .A1(i_data_bus[451]), .A2(n10410), .B1(
        i_data_bus[483]), .B2(n10412), .ZN(n8522) );
  AOI22D1BWP30P140LVT U12509 ( .A1(i_data_bus[387]), .A2(n10409), .B1(
        i_data_bus[419]), .B2(n10411), .ZN(n8521) );
  ND2D1BWP30P140LVT U12510 ( .A1(n8522), .A2(n8521), .ZN(N14340) );
  AOI22D1BWP30P140LVT U12511 ( .A1(i_data_bus[473]), .A2(n10410), .B1(
        i_data_bus[505]), .B2(n10412), .ZN(n8524) );
  AOI22D1BWP30P140LVT U12512 ( .A1(i_data_bus[409]), .A2(n10409), .B1(
        i_data_bus[441]), .B2(n10411), .ZN(n8523) );
  ND2D1BWP30P140LVT U12513 ( .A1(n8524), .A2(n8523), .ZN(N14362) );
  AOI22D1BWP30P140LVT U12514 ( .A1(i_data_bus[437]), .A2(n10601), .B1(
        i_data_bus[501]), .B2(n10602), .ZN(n8526) );
  AOI22D1BWP30P140LVT U12515 ( .A1(i_data_bus[405]), .A2(n10603), .B1(
        i_data_bus[469]), .B2(n10604), .ZN(n8525) );
  ND2D1BWP30P140LVT U12516 ( .A1(n8526), .A2(n8525), .ZN(N3114) );
  AOI22D1BWP30P140LVT U12517 ( .A1(i_data_bus[502]), .A2(n10602), .B1(
        i_data_bus[438]), .B2(n10601), .ZN(n8528) );
  AOI22D1BWP30P140LVT U12518 ( .A1(i_data_bus[406]), .A2(n10603), .B1(
        i_data_bus[470]), .B2(n10604), .ZN(n8527) );
  ND2D1BWP30P140LVT U12519 ( .A1(n8528), .A2(n8527), .ZN(N3115) );
  AOI22D1BWP30P140LVT U12520 ( .A1(i_data_bus[416]), .A2(n10601), .B1(
        i_data_bus[480]), .B2(n10602), .ZN(n8530) );
  AOI22D1BWP30P140LVT U12521 ( .A1(i_data_bus[384]), .A2(n10603), .B1(
        i_data_bus[448]), .B2(n10604), .ZN(n8529) );
  ND2D1BWP30P140LVT U12522 ( .A1(n8530), .A2(n8529), .ZN(N3093) );
  AOI22D1BWP30P140LVT U12523 ( .A1(i_data_bus[429]), .A2(n10601), .B1(
        i_data_bus[493]), .B2(n10602), .ZN(n8532) );
  AOI22D1BWP30P140LVT U12524 ( .A1(i_data_bus[397]), .A2(n10603), .B1(
        i_data_bus[461]), .B2(n10604), .ZN(n8531) );
  ND2D1BWP30P140LVT U12525 ( .A1(n8532), .A2(n8531), .ZN(N3106) );
  AOI22D1BWP30P140LVT U12526 ( .A1(i_data_bus[509]), .A2(n10602), .B1(
        i_data_bus[445]), .B2(n10601), .ZN(n8534) );
  AOI22D1BWP30P140LVT U12527 ( .A1(i_data_bus[413]), .A2(n10603), .B1(
        i_data_bus[477]), .B2(n10604), .ZN(n8533) );
  ND2D1BWP30P140LVT U12528 ( .A1(n8534), .A2(n8533), .ZN(N3122) );
  AOI22D1BWP30P140LVT U12529 ( .A1(i_data_bus[385]), .A2(n10603), .B1(
        i_data_bus[417]), .B2(n10601), .ZN(n8536) );
  AOI22D1BWP30P140LVT U12530 ( .A1(i_data_bus[481]), .A2(n10602), .B1(
        i_data_bus[449]), .B2(n10604), .ZN(n8535) );
  ND2D1BWP30P140LVT U12531 ( .A1(n8536), .A2(n8535), .ZN(N3094) );
  AOI22D1BWP30P140LVT U12532 ( .A1(i_data_bus[498]), .A2(n10602), .B1(
        i_data_bus[402]), .B2(n10603), .ZN(n8538) );
  AOI22D1BWP30P140LVT U12533 ( .A1(i_data_bus[434]), .A2(n10601), .B1(
        i_data_bus[466]), .B2(n10604), .ZN(n8537) );
  ND2D1BWP30P140LVT U12534 ( .A1(n8538), .A2(n8537), .ZN(N3111) );
  AOI22D1BWP30P140LVT U12535 ( .A1(i_data_bus[389]), .A2(n10603), .B1(
        i_data_bus[485]), .B2(n10602), .ZN(n8540) );
  AOI22D1BWP30P140LVT U12536 ( .A1(i_data_bus[421]), .A2(n10601), .B1(
        i_data_bus[453]), .B2(n10604), .ZN(n8539) );
  ND2D1BWP30P140LVT U12537 ( .A1(n8540), .A2(n8539), .ZN(N3098) );
  AOI22D1BWP30P140LVT U12538 ( .A1(i_data_bus[427]), .A2(n10601), .B1(
        i_data_bus[491]), .B2(n10602), .ZN(n8542) );
  AOI22D1BWP30P140LVT U12539 ( .A1(i_data_bus[395]), .A2(n10603), .B1(
        i_data_bus[459]), .B2(n10604), .ZN(n8541) );
  ND2D1BWP30P140LVT U12540 ( .A1(n8542), .A2(n8541), .ZN(N3104) );
  AOI22D1BWP30P140LVT U12541 ( .A1(i_data_bus[414]), .A2(n10603), .B1(
        i_data_bus[510]), .B2(n10602), .ZN(n8544) );
  AOI22D1BWP30P140LVT U12542 ( .A1(i_data_bus[446]), .A2(n10601), .B1(
        i_data_bus[478]), .B2(n10604), .ZN(n8543) );
  ND2D1BWP30P140LVT U12543 ( .A1(n8544), .A2(n8543), .ZN(N3123) );
  AOI22D1BWP30P140LVT U12544 ( .A1(i_data_bus[767]), .A2(n10466), .B1(
        i_data_bus[671]), .B2(n10467), .ZN(n8546) );
  AOI22D1BWP30P140LVT U12545 ( .A1(i_data_bus[703]), .A2(n10468), .B1(
        i_data_bus[735]), .B2(n10465), .ZN(n8545) );
  ND2D1BWP30P140LVT U12546 ( .A1(n8546), .A2(n8545), .ZN(N11052) );
  AOI22D1BWP30P140LVT U12547 ( .A1(i_data_bus[675]), .A2(n10468), .B1(
        i_data_bus[739]), .B2(n10466), .ZN(n8548) );
  AOI22D1BWP30P140LVT U12548 ( .A1(i_data_bus[643]), .A2(n10467), .B1(
        i_data_bus[707]), .B2(n10465), .ZN(n8547) );
  ND2D1BWP30P140LVT U12549 ( .A1(n8548), .A2(n8547), .ZN(N11024) );
  AOI22D1BWP30P140LVT U12550 ( .A1(i_data_bus[746]), .A2(n10466), .B1(
        i_data_bus[682]), .B2(n10468), .ZN(n8550) );
  AOI22D1BWP30P140LVT U12551 ( .A1(i_data_bus[650]), .A2(n10467), .B1(
        i_data_bus[714]), .B2(n10465), .ZN(n8549) );
  ND2D1BWP30P140LVT U12552 ( .A1(n8550), .A2(n8549), .ZN(N11031) );
  AOI22D1BWP30P140LVT U12553 ( .A1(i_data_bus[665]), .A2(n10467), .B1(
        i_data_bus[761]), .B2(n10466), .ZN(n8552) );
  AOI22D1BWP30P140LVT U12554 ( .A1(i_data_bus[697]), .A2(n10468), .B1(
        i_data_bus[729]), .B2(n10465), .ZN(n8551) );
  ND2D1BWP30P140LVT U12555 ( .A1(n8552), .A2(n8551), .ZN(N11046) );
  AOI22D1BWP30P140LVT U12556 ( .A1(i_data_bus[644]), .A2(n10467), .B1(
        i_data_bus[676]), .B2(n10468), .ZN(n8554) );
  AOI22D1BWP30P140LVT U12557 ( .A1(i_data_bus[740]), .A2(n10466), .B1(
        i_data_bus[708]), .B2(n10465), .ZN(n8553) );
  ND2D1BWP30P140LVT U12558 ( .A1(n8554), .A2(n8553), .ZN(N11025) );
  AOI22D1BWP30P140LVT U12559 ( .A1(i_data_bus[763]), .A2(n10466), .B1(
        i_data_bus[699]), .B2(n10468), .ZN(n8556) );
  AOI22D1BWP30P140LVT U12560 ( .A1(i_data_bus[667]), .A2(n10467), .B1(
        i_data_bus[731]), .B2(n10465), .ZN(n8555) );
  ND2D1BWP30P140LVT U12561 ( .A1(n8556), .A2(n8555), .ZN(N11048) );
  AOI22D1BWP30P140LVT U12562 ( .A1(i_data_bus[653]), .A2(n10467), .B1(
        i_data_bus[685]), .B2(n10468), .ZN(n8558) );
  AOI22D1BWP30P140LVT U12563 ( .A1(i_data_bus[749]), .A2(n10466), .B1(
        i_data_bus[717]), .B2(n10465), .ZN(n8557) );
  ND2D1BWP30P140LVT U12564 ( .A1(n8558), .A2(n8557), .ZN(N11034) );
  AOI22D1BWP30P140LVT U12565 ( .A1(i_data_bus[752]), .A2(n10530), .B1(
        i_data_bus[720]), .B2(n10531), .ZN(n8560) );
  AOI22D1BWP30P140LVT U12566 ( .A1(i_data_bus[688]), .A2(n10532), .B1(
        i_data_bus[656]), .B2(n10529), .ZN(n8559) );
  ND2D1BWP30P140LVT U12567 ( .A1(n8560), .A2(n8559), .ZN(N7289) );
  AOI22D1BWP30P140LVT U12568 ( .A1(i_data_bus[703]), .A2(n10532), .B1(
        i_data_bus[735]), .B2(n10531), .ZN(n8562) );
  AOI22D1BWP30P140LVT U12569 ( .A1(i_data_bus[767]), .A2(n10530), .B1(
        i_data_bus[671]), .B2(n10529), .ZN(n8561) );
  ND2D1BWP30P140LVT U12570 ( .A1(n8562), .A2(n8561), .ZN(N7304) );
  AOI22D1BWP30P140LVT U12571 ( .A1(i_data_bus[709]), .A2(n10531), .B1(
        i_data_bus[741]), .B2(n10530), .ZN(n8564) );
  AOI22D1BWP30P140LVT U12572 ( .A1(i_data_bus[677]), .A2(n10532), .B1(
        i_data_bus[645]), .B2(n10529), .ZN(n8563) );
  ND2D1BWP30P140LVT U12573 ( .A1(n8564), .A2(n8563), .ZN(N7278) );
  AOI22D1BWP30P140LVT U12574 ( .A1(i_data_bus[712]), .A2(n10531), .B1(
        i_data_bus[680]), .B2(n10532), .ZN(n8566) );
  AOI22D1BWP30P140LVT U12575 ( .A1(i_data_bus[744]), .A2(n10530), .B1(
        i_data_bus[648]), .B2(n10529), .ZN(n8565) );
  ND2D1BWP30P140LVT U12576 ( .A1(n8566), .A2(n8565), .ZN(N7281) );
  AOI22D1BWP30P140LVT U12577 ( .A1(i_data_bus[740]), .A2(n10530), .B1(
        i_data_bus[676]), .B2(n10532), .ZN(n8568) );
  AOI22D1BWP30P140LVT U12578 ( .A1(i_data_bus[708]), .A2(n10531), .B1(
        i_data_bus[644]), .B2(n10529), .ZN(n8567) );
  ND2D1BWP30P140LVT U12579 ( .A1(n8568), .A2(n8567), .ZN(N7277) );
  AOI22D1BWP30P140LVT U12580 ( .A1(i_data_bus[730]), .A2(n10531), .B1(
        i_data_bus[762]), .B2(n10530), .ZN(n8570) );
  AOI22D1BWP30P140LVT U12581 ( .A1(i_data_bus[698]), .A2(n10532), .B1(
        i_data_bus[666]), .B2(n10529), .ZN(n8569) );
  ND2D1BWP30P140LVT U12582 ( .A1(n8570), .A2(n8569), .ZN(N7299) );
  AOI22D1BWP30P140LVT U12583 ( .A1(i_data_bus[686]), .A2(n10532), .B1(
        i_data_bus[750]), .B2(n10530), .ZN(n8572) );
  AOI22D1BWP30P140LVT U12584 ( .A1(i_data_bus[718]), .A2(n10531), .B1(
        i_data_bus[654]), .B2(n10529), .ZN(n8571) );
  ND2D1BWP30P140LVT U12585 ( .A1(n8572), .A2(n8571), .ZN(N7287) );
  AOI22D1BWP30P140LVT U12586 ( .A1(i_data_bus[679]), .A2(n10532), .B1(
        i_data_bus[743]), .B2(n10530), .ZN(n8574) );
  AOI22D1BWP30P140LVT U12587 ( .A1(i_data_bus[711]), .A2(n10531), .B1(
        i_data_bus[647]), .B2(n10529), .ZN(n8573) );
  ND2D1BWP30P140LVT U12588 ( .A1(n8574), .A2(n8573), .ZN(N7280) );
  AOI22D1BWP30P140LVT U12589 ( .A1(i_data_bus[719]), .A2(n10531), .B1(
        i_data_bus[687]), .B2(n10532), .ZN(n8576) );
  AOI22D1BWP30P140LVT U12590 ( .A1(i_data_bus[751]), .A2(n10530), .B1(
        i_data_bus[655]), .B2(n10529), .ZN(n8575) );
  ND2D1BWP30P140LVT U12591 ( .A1(n8576), .A2(n8575), .ZN(N7288) );
  AOI22D1BWP30P140LVT U12592 ( .A1(i_data_bus[694]), .A2(n10532), .B1(
        i_data_bus[726]), .B2(n10531), .ZN(n8578) );
  AOI22D1BWP30P140LVT U12593 ( .A1(i_data_bus[758]), .A2(n10530), .B1(
        i_data_bus[662]), .B2(n10529), .ZN(n8577) );
  ND2D1BWP30P140LVT U12594 ( .A1(n8578), .A2(n8577), .ZN(N7295) );
  AOI22D1BWP30P140LVT U12595 ( .A1(i_data_bus[587]), .A2(n10565), .B1(
        i_data_bus[523]), .B2(n10566), .ZN(n8580) );
  AOI22D1BWP30P140LVT U12596 ( .A1(i_data_bus[619]), .A2(n10568), .B1(
        i_data_bus[555]), .B2(n10567), .ZN(n8579) );
  ND2D1BWP30P140LVT U12597 ( .A1(n8580), .A2(n8579), .ZN(N5194) );
  AOI22D1BWP30P140LVT U12598 ( .A1(i_data_bus[611]), .A2(n10568), .B1(
        i_data_bus[515]), .B2(n10566), .ZN(n8582) );
  AOI22D1BWP30P140LVT U12599 ( .A1(i_data_bus[579]), .A2(n10565), .B1(
        i_data_bus[547]), .B2(n10567), .ZN(n8581) );
  ND2D1BWP30P140LVT U12600 ( .A1(n8582), .A2(n8581), .ZN(N5186) );
  AOI22D1BWP30P140LVT U12601 ( .A1(i_data_bus[631]), .A2(n10568), .B1(
        i_data_bus[535]), .B2(n10566), .ZN(n8584) );
  AOI22D1BWP30P140LVT U12602 ( .A1(i_data_bus[599]), .A2(n10565), .B1(
        i_data_bus[567]), .B2(n10567), .ZN(n8583) );
  ND2D1BWP30P140LVT U12603 ( .A1(n8584), .A2(n8583), .ZN(N5206) );
  AOI22D1BWP30P140LVT U12604 ( .A1(i_data_bus[577]), .A2(n10565), .B1(
        i_data_bus[609]), .B2(n10568), .ZN(n8586) );
  AOI22D1BWP30P140LVT U12605 ( .A1(i_data_bus[513]), .A2(n10566), .B1(
        i_data_bus[545]), .B2(n10567), .ZN(n8585) );
  ND2D1BWP30P140LVT U12606 ( .A1(n8586), .A2(n8585), .ZN(N5184) );
  AOI22D1BWP30P140LVT U12607 ( .A1(i_data_bus[512]), .A2(n10566), .B1(
        i_data_bus[576]), .B2(n10565), .ZN(n8588) );
  AOI22D1BWP30P140LVT U12608 ( .A1(i_data_bus[608]), .A2(n10568), .B1(
        i_data_bus[544]), .B2(n10567), .ZN(n8587) );
  ND2D1BWP30P140LVT U12609 ( .A1(n8588), .A2(n8587), .ZN(N5183) );
  AOI22D1BWP30P140LVT U12610 ( .A1(i_data_bus[519]), .A2(n10566), .B1(
        i_data_bus[583]), .B2(n10565), .ZN(n8590) );
  AOI22D1BWP30P140LVT U12611 ( .A1(i_data_bus[615]), .A2(n10568), .B1(
        i_data_bus[551]), .B2(n10567), .ZN(n8589) );
  ND2D1BWP30P140LVT U12612 ( .A1(n8590), .A2(n8589), .ZN(N5190) );
  AOI22D1BWP30P140LVT U12613 ( .A1(i_data_bus[597]), .A2(n10565), .B1(
        i_data_bus[629]), .B2(n10568), .ZN(n8592) );
  AOI22D1BWP30P140LVT U12614 ( .A1(i_data_bus[533]), .A2(n10566), .B1(
        i_data_bus[565]), .B2(n10567), .ZN(n8591) );
  ND2D1BWP30P140LVT U12615 ( .A1(n8592), .A2(n8591), .ZN(N5204) );
  AOI22D1BWP30P140LVT U12616 ( .A1(i_data_bus[698]), .A2(n10593), .B1(
        i_data_bus[762]), .B2(n10595), .ZN(n8594) );
  AOI22D1BWP30P140LVT U12617 ( .A1(i_data_bus[666]), .A2(n10596), .B1(
        i_data_bus[730]), .B2(n10594), .ZN(n8593) );
  ND2D1BWP30P140LVT U12618 ( .A1(n8594), .A2(n8593), .ZN(N3551) );
  AOI22D1BWP30P140LVT U12619 ( .A1(i_data_bus[657]), .A2(n10596), .B1(
        i_data_bus[689]), .B2(n10593), .ZN(n8596) );
  AOI22D1BWP30P140LVT U12620 ( .A1(i_data_bus[753]), .A2(n10595), .B1(
        i_data_bus[721]), .B2(n10594), .ZN(n8595) );
  ND2D1BWP30P140LVT U12621 ( .A1(n8596), .A2(n8595), .ZN(N3542) );
  AOI22D1BWP30P140LVT U12622 ( .A1(i_data_bus[665]), .A2(n10596), .B1(
        i_data_bus[761]), .B2(n10595), .ZN(n8598) );
  AOI22D1BWP30P140LVT U12623 ( .A1(i_data_bus[697]), .A2(n10593), .B1(
        i_data_bus[729]), .B2(n10594), .ZN(n8597) );
  ND2D1BWP30P140LVT U12624 ( .A1(n8598), .A2(n8597), .ZN(N3550) );
  AOI22D1BWP30P140LVT U12625 ( .A1(i_data_bus[648]), .A2(n10596), .B1(
        i_data_bus[680]), .B2(n10593), .ZN(n8600) );
  AOI22D1BWP30P140LVT U12626 ( .A1(i_data_bus[744]), .A2(n10595), .B1(
        i_data_bus[712]), .B2(n10594), .ZN(n8599) );
  ND2D1BWP30P140LVT U12627 ( .A1(n8600), .A2(n8599), .ZN(N3533) );
  AOI22D1BWP30P140LVT U12628 ( .A1(i_data_bus[765]), .A2(n10595), .B1(
        i_data_bus[701]), .B2(n10593), .ZN(n8602) );
  AOI22D1BWP30P140LVT U12629 ( .A1(i_data_bus[669]), .A2(n10596), .B1(
        i_data_bus[733]), .B2(n10594), .ZN(n8601) );
  ND2D1BWP30P140LVT U12630 ( .A1(n8602), .A2(n8601), .ZN(N3554) );
  AOI22D1BWP30P140LVT U12631 ( .A1(i_data_bus[653]), .A2(n10596), .B1(
        i_data_bus[685]), .B2(n10593), .ZN(n8604) );
  AOI22D1BWP30P140LVT U12632 ( .A1(i_data_bus[749]), .A2(n10595), .B1(
        i_data_bus[717]), .B2(n10594), .ZN(n8603) );
  ND2D1BWP30P140LVT U12633 ( .A1(n8604), .A2(n8603), .ZN(N3538) );
  AOI22D1BWP30P140LVT U12634 ( .A1(i_data_bus[651]), .A2(n10435), .B1(
        i_data_bus[683]), .B2(n10436), .ZN(n8606) );
  AOI22D1BWP30P140LVT U12635 ( .A1(i_data_bus[715]), .A2(n10434), .B1(
        i_data_bus[747]), .B2(n10433), .ZN(n8605) );
  ND2D1BWP30P140LVT U12636 ( .A1(n8606), .A2(n8605), .ZN(N12906) );
  AOI22D1BWP30P140LVT U12637 ( .A1(i_data_bus[710]), .A2(n10434), .B1(
        i_data_bus[678]), .B2(n10436), .ZN(n8608) );
  AOI22D1BWP30P140LVT U12638 ( .A1(i_data_bus[646]), .A2(n10435), .B1(
        i_data_bus[742]), .B2(n10433), .ZN(n8607) );
  ND2D1BWP30P140LVT U12639 ( .A1(n8608), .A2(n8607), .ZN(N12901) );
  AOI22D1BWP30P140LVT U12640 ( .A1(i_data_bus[726]), .A2(n10434), .B1(
        i_data_bus[662]), .B2(n10435), .ZN(n8610) );
  AOI22D1BWP30P140LVT U12641 ( .A1(i_data_bus[694]), .A2(n10436), .B1(
        i_data_bus[758]), .B2(n10433), .ZN(n8609) );
  ND2D1BWP30P140LVT U12642 ( .A1(n8610), .A2(n8609), .ZN(N12917) );
  AOI22D1BWP30P140LVT U12643 ( .A1(i_data_bus[700]), .A2(n10436), .B1(
        i_data_bus[668]), .B2(n10435), .ZN(n8612) );
  AOI22D1BWP30P140LVT U12644 ( .A1(i_data_bus[732]), .A2(n10434), .B1(
        i_data_bus[764]), .B2(n10433), .ZN(n8611) );
  ND2D1BWP30P140LVT U12645 ( .A1(n8612), .A2(n8611), .ZN(N12923) );
  AOI22D1BWP30P140LVT U12646 ( .A1(i_data_bus[692]), .A2(n10436), .B1(
        i_data_bus[724]), .B2(n10434), .ZN(n8614) );
  AOI22D1BWP30P140LVT U12647 ( .A1(i_data_bus[660]), .A2(n10435), .B1(
        i_data_bus[756]), .B2(n10433), .ZN(n8613) );
  ND2D1BWP30P140LVT U12648 ( .A1(n8614), .A2(n8613), .ZN(N12915) );
  AOI22D1BWP30P140LVT U12649 ( .A1(i_data_bus[666]), .A2(n10435), .B1(
        i_data_bus[730]), .B2(n10434), .ZN(n8616) );
  AOI22D1BWP30P140LVT U12650 ( .A1(i_data_bus[698]), .A2(n10436), .B1(
        i_data_bus[762]), .B2(n10433), .ZN(n8615) );
  ND2D1BWP30P140LVT U12651 ( .A1(n8616), .A2(n8615), .ZN(N12921) );
  AOI22D1BWP30P140LVT U12652 ( .A1(i_data_bus[659]), .A2(n10498), .B1(
        i_data_bus[723]), .B2(n10497), .ZN(n8618) );
  AOI22D1BWP30P140LVT U12653 ( .A1(i_data_bus[755]), .A2(n10500), .B1(
        i_data_bus[691]), .B2(n10499), .ZN(n8617) );
  ND2D1BWP30P140LVT U12654 ( .A1(n8618), .A2(n8617), .ZN(N9166) );
  AOI22D1BWP30P140LVT U12655 ( .A1(i_data_bus[725]), .A2(n10497), .B1(
        i_data_bus[661]), .B2(n10498), .ZN(n8620) );
  AOI22D1BWP30P140LVT U12656 ( .A1(i_data_bus[757]), .A2(n10500), .B1(
        i_data_bus[693]), .B2(n10499), .ZN(n8619) );
  ND2D1BWP30P140LVT U12657 ( .A1(n8620), .A2(n8619), .ZN(N9168) );
  AOI22D1BWP30P140LVT U12658 ( .A1(i_data_bus[652]), .A2(n10498), .B1(
        i_data_bus[748]), .B2(n10500), .ZN(n8622) );
  AOI22D1BWP30P140LVT U12659 ( .A1(i_data_bus[716]), .A2(n10497), .B1(
        i_data_bus[684]), .B2(n10499), .ZN(n8621) );
  ND2D1BWP30P140LVT U12660 ( .A1(n8622), .A2(n8621), .ZN(N9159) );
  AOI22D1BWP30P140LVT U12661 ( .A1(i_data_bus[645]), .A2(n10498), .B1(
        i_data_bus[741]), .B2(n10500), .ZN(n8624) );
  AOI22D1BWP30P140LVT U12662 ( .A1(i_data_bus[709]), .A2(n10497), .B1(
        i_data_bus[677]), .B2(n10499), .ZN(n8623) );
  ND2D1BWP30P140LVT U12663 ( .A1(n8624), .A2(n8623), .ZN(N9152) );
  AOI22D1BWP30P140LVT U12664 ( .A1(i_data_bus[649]), .A2(n10498), .B1(
        i_data_bus[745]), .B2(n10500), .ZN(n8626) );
  AOI22D1BWP30P140LVT U12665 ( .A1(i_data_bus[713]), .A2(n10497), .B1(
        i_data_bus[681]), .B2(n10499), .ZN(n8625) );
  ND2D1BWP30P140LVT U12666 ( .A1(n8626), .A2(n8625), .ZN(N9156) );
  AOI22D1BWP30P140LVT U12667 ( .A1(i_data_bus[707]), .A2(n10497), .B1(
        i_data_bus[739]), .B2(n10500), .ZN(n8628) );
  AOI22D1BWP30P140LVT U12668 ( .A1(i_data_bus[643]), .A2(n10498), .B1(
        i_data_bus[675]), .B2(n10499), .ZN(n8627) );
  ND2D1BWP30P140LVT U12669 ( .A1(n8628), .A2(n8627), .ZN(N9150) );
  AOI22D1BWP30P140LVT U12670 ( .A1(i_data_bus[740]), .A2(n10500), .B1(
        i_data_bus[644]), .B2(n10498), .ZN(n8630) );
  AOI22D1BWP30P140LVT U12671 ( .A1(i_data_bus[708]), .A2(n10497), .B1(
        i_data_bus[676]), .B2(n10499), .ZN(n8629) );
  ND2D1BWP30P140LVT U12672 ( .A1(n8630), .A2(n8629), .ZN(N9151) );
  AOI22D1BWP30P140LVT U12673 ( .A1(i_data_bus[752]), .A2(n10500), .B1(
        i_data_bus[656]), .B2(n10498), .ZN(n8632) );
  AOI22D1BWP30P140LVT U12674 ( .A1(i_data_bus[720]), .A2(n10497), .B1(
        i_data_bus[688]), .B2(n10499), .ZN(n8631) );
  ND2D1BWP30P140LVT U12675 ( .A1(n8632), .A2(n8631), .ZN(N9163) );
  AOI22D1BWP30P140LVT U12676 ( .A1(i_data_bus[669]), .A2(n10498), .B1(
        i_data_bus[733]), .B2(n10497), .ZN(n8634) );
  AOI22D1BWP30P140LVT U12677 ( .A1(i_data_bus[765]), .A2(n10500), .B1(
        i_data_bus[701]), .B2(n10499), .ZN(n8633) );
  ND2D1BWP30P140LVT U12678 ( .A1(n8634), .A2(n8633), .ZN(N9176) );
  AOI22D1BWP30P140LVT U12679 ( .A1(i_data_bus[783]), .A2(n10462), .B1(
        i_data_bus[815]), .B2(n10464), .ZN(n8636) );
  AOI22D1BWP30P140LVT U12680 ( .A1(i_data_bus[879]), .A2(n10461), .B1(
        i_data_bus[847]), .B2(n10463), .ZN(n8635) );
  ND2D1BWP30P140LVT U12681 ( .A1(n8636), .A2(n8635), .ZN(N11252) );
  AOI22D1BWP30P140LVT U12682 ( .A1(i_data_bus[771]), .A2(n10462), .B1(
        i_data_bus[803]), .B2(n10464), .ZN(n8638) );
  AOI22D1BWP30P140LVT U12683 ( .A1(i_data_bus[867]), .A2(n10461), .B1(
        i_data_bus[835]), .B2(n10463), .ZN(n8637) );
  ND2D1BWP30P140LVT U12684 ( .A1(n8638), .A2(n8637), .ZN(N11240) );
  AOI22D1BWP30P140LVT U12685 ( .A1(i_data_bus[801]), .A2(n10464), .B1(
        i_data_bus[865]), .B2(n10461), .ZN(n8640) );
  AOI22D1BWP30P140LVT U12686 ( .A1(i_data_bus[769]), .A2(n10462), .B1(
        i_data_bus[833]), .B2(n10463), .ZN(n8639) );
  ND2D1BWP30P140LVT U12687 ( .A1(n8640), .A2(n8639), .ZN(N11238) );
  AOI22D1BWP30P140LVT U12688 ( .A1(i_data_bus[885]), .A2(n10461), .B1(
        i_data_bus[821]), .B2(n10464), .ZN(n8642) );
  AOI22D1BWP30P140LVT U12689 ( .A1(i_data_bus[789]), .A2(n10462), .B1(
        i_data_bus[853]), .B2(n10463), .ZN(n8641) );
  ND2D1BWP30P140LVT U12690 ( .A1(n8642), .A2(n8641), .ZN(N11258) );
  AOI22D1BWP30P140LVT U12691 ( .A1(i_data_bus[810]), .A2(n10464), .B1(
        i_data_bus[874]), .B2(n10461), .ZN(n8644) );
  AOI22D1BWP30P140LVT U12692 ( .A1(i_data_bus[778]), .A2(n10462), .B1(
        i_data_bus[842]), .B2(n10463), .ZN(n8643) );
  ND2D1BWP30P140LVT U12693 ( .A1(n8644), .A2(n8643), .ZN(N11247) );
  AOI22D1BWP30P140LVT U12694 ( .A1(i_data_bus[805]), .A2(n10464), .B1(
        i_data_bus[773]), .B2(n10462), .ZN(n8646) );
  AOI22D1BWP30P140LVT U12695 ( .A1(i_data_bus[869]), .A2(n10461), .B1(
        i_data_bus[837]), .B2(n10463), .ZN(n8645) );
  ND2D1BWP30P140LVT U12696 ( .A1(n8646), .A2(n8645), .ZN(N11242) );
  AOI22D1BWP30P140LVT U12697 ( .A1(i_data_bus[870]), .A2(n10461), .B1(
        i_data_bus[774]), .B2(n10462), .ZN(n8648) );
  AOI22D1BWP30P140LVT U12698 ( .A1(i_data_bus[806]), .A2(n10464), .B1(
        i_data_bus[838]), .B2(n10463), .ZN(n8647) );
  ND2D1BWP30P140LVT U12699 ( .A1(n8648), .A2(n8647), .ZN(N11243) );
  AOI22D1BWP30P140LVT U12700 ( .A1(i_data_bus[820]), .A2(n10464), .B1(
        i_data_bus[884]), .B2(n10461), .ZN(n8650) );
  AOI22D1BWP30P140LVT U12701 ( .A1(i_data_bus[788]), .A2(n10462), .B1(
        i_data_bus[852]), .B2(n10463), .ZN(n8649) );
  ND2D1BWP30P140LVT U12702 ( .A1(n8650), .A2(n8649), .ZN(N11257) );
  AOI22D1BWP30P140LVT U12703 ( .A1(i_data_bus[807]), .A2(n10464), .B1(
        i_data_bus[775]), .B2(n10462), .ZN(n8652) );
  AOI22D1BWP30P140LVT U12704 ( .A1(i_data_bus[871]), .A2(n10461), .B1(
        i_data_bus[839]), .B2(n10463), .ZN(n8651) );
  ND2D1BWP30P140LVT U12705 ( .A1(n8652), .A2(n8651), .ZN(N11244) );
  AOI22D1BWP30P140LVT U12706 ( .A1(i_data_bus[988]), .A2(n10555), .B1(
        i_data_bus[956]), .B2(n10553), .ZN(n8654) );
  AOI22D1BWP30P140LVT U12707 ( .A1(i_data_bus[924]), .A2(n10554), .B1(
        i_data_bus[1020]), .B2(n10556), .ZN(n8653) );
  ND2D1BWP30P140LVT U12708 ( .A1(n8654), .A2(n8653), .ZN(N5859) );
  AOI22D1BWP30P140LVT U12709 ( .A1(i_data_bus[961]), .A2(n10555), .B1(
        i_data_bus[897]), .B2(n10554), .ZN(n8656) );
  AOI22D1BWP30P140LVT U12710 ( .A1(i_data_bus[929]), .A2(n10553), .B1(
        i_data_bus[993]), .B2(n10556), .ZN(n8655) );
  ND2D1BWP30P140LVT U12711 ( .A1(n8656), .A2(n8655), .ZN(N5832) );
  AOI22D1BWP30P140LVT U12712 ( .A1(i_data_bus[898]), .A2(n10554), .B1(
        i_data_bus[930]), .B2(n10553), .ZN(n8658) );
  AOI22D1BWP30P140LVT U12713 ( .A1(i_data_bus[962]), .A2(n10555), .B1(
        i_data_bus[994]), .B2(n10556), .ZN(n8657) );
  ND2D1BWP30P140LVT U12714 ( .A1(n8658), .A2(n8657), .ZN(N5833) );
  AOI22D1BWP30P140LVT U12715 ( .A1(i_data_bus[971]), .A2(n10555), .B1(
        i_data_bus[907]), .B2(n10554), .ZN(n8660) );
  AOI22D1BWP30P140LVT U12716 ( .A1(i_data_bus[939]), .A2(n10553), .B1(
        i_data_bus[1003]), .B2(n10556), .ZN(n8659) );
  ND2D1BWP30P140LVT U12717 ( .A1(n8660), .A2(n8659), .ZN(N5842) );
  AOI22D1BWP30P140LVT U12718 ( .A1(i_data_bus[946]), .A2(n10553), .B1(
        i_data_bus[914]), .B2(n10554), .ZN(n8662) );
  AOI22D1BWP30P140LVT U12719 ( .A1(i_data_bus[978]), .A2(n10555), .B1(
        i_data_bus[1010]), .B2(n10556), .ZN(n8661) );
  ND2D1BWP30P140LVT U12720 ( .A1(n8662), .A2(n8661), .ZN(N5849) );
  AOI22D1BWP30P140LVT U12721 ( .A1(i_data_bus[951]), .A2(n10553), .B1(
        i_data_bus[983]), .B2(n10555), .ZN(n8664) );
  AOI22D1BWP30P140LVT U12722 ( .A1(i_data_bus[919]), .A2(n10554), .B1(
        i_data_bus[1015]), .B2(n10556), .ZN(n8663) );
  ND2D1BWP30P140LVT U12723 ( .A1(n8664), .A2(n8663), .ZN(N5854) );
  AOI22D1BWP30P140LVT U12724 ( .A1(i_data_bus[985]), .A2(n10555), .B1(
        i_data_bus[921]), .B2(n10554), .ZN(n8666) );
  AOI22D1BWP30P140LVT U12725 ( .A1(i_data_bus[953]), .A2(n10553), .B1(
        i_data_bus[1017]), .B2(n10556), .ZN(n8665) );
  ND2D1BWP30P140LVT U12726 ( .A1(n8666), .A2(n8665), .ZN(N5856) );
  AOI22D1BWP30P140LVT U12727 ( .A1(i_data_bus[955]), .A2(n10553), .B1(
        i_data_bus[923]), .B2(n10554), .ZN(n8668) );
  AOI22D1BWP30P140LVT U12728 ( .A1(i_data_bus[987]), .A2(n10555), .B1(
        i_data_bus[1019]), .B2(n10556), .ZN(n8667) );
  ND2D1BWP30P140LVT U12729 ( .A1(n8668), .A2(n8667), .ZN(N5858) );
  AOI22D1BWP30P140LVT U12730 ( .A1(i_data_bus[925]), .A2(n10554), .B1(
        i_data_bus[957]), .B2(n10553), .ZN(n8670) );
  AOI22D1BWP30P140LVT U12731 ( .A1(i_data_bus[989]), .A2(n10555), .B1(
        i_data_bus[1021]), .B2(n10556), .ZN(n8669) );
  ND2D1BWP30P140LVT U12732 ( .A1(n8670), .A2(n8669), .ZN(N5860) );
  AOI22D1BWP30P140LVT U12733 ( .A1(i_data_bus[482]), .A2(n10412), .B1(
        i_data_bus[386]), .B2(n10409), .ZN(n8672) );
  AOI22D1BWP30P140LVT U12734 ( .A1(i_data_bus[418]), .A2(n10411), .B1(
        i_data_bus[450]), .B2(n10410), .ZN(n8671) );
  ND2D1BWP30P140LVT U12735 ( .A1(n8672), .A2(n8671), .ZN(N14339) );
  AOI22D1BWP30P140LVT U12736 ( .A1(i_data_bus[417]), .A2(n10411), .B1(
        i_data_bus[481]), .B2(n10412), .ZN(n8674) );
  AOI22D1BWP30P140LVT U12737 ( .A1(i_data_bus[385]), .A2(n10409), .B1(
        i_data_bus[449]), .B2(n10410), .ZN(n8673) );
  ND2D1BWP30P140LVT U12738 ( .A1(n8674), .A2(n8673), .ZN(N14338) );
  AOI22D1BWP30P140LVT U12739 ( .A1(i_data_bus[427]), .A2(n10411), .B1(
        i_data_bus[491]), .B2(n10412), .ZN(n8676) );
  AOI22D1BWP30P140LVT U12740 ( .A1(i_data_bus[395]), .A2(n10409), .B1(
        i_data_bus[459]), .B2(n10410), .ZN(n8675) );
  ND2D1BWP30P140LVT U12741 ( .A1(n8676), .A2(n8675), .ZN(N14348) );
  AOI22D1BWP30P140LVT U12742 ( .A1(i_data_bus[392]), .A2(n10409), .B1(
        i_data_bus[424]), .B2(n10411), .ZN(n8678) );
  AOI22D1BWP30P140LVT U12743 ( .A1(i_data_bus[488]), .A2(n10412), .B1(
        i_data_bus[456]), .B2(n10410), .ZN(n8677) );
  ND2D1BWP30P140LVT U12744 ( .A1(n8678), .A2(n8677), .ZN(N14345) );
  AOI22D1BWP30P140LVT U12745 ( .A1(i_data_bus[406]), .A2(n10409), .B1(
        i_data_bus[438]), .B2(n10411), .ZN(n8680) );
  AOI22D1BWP30P140LVT U12746 ( .A1(i_data_bus[502]), .A2(n10412), .B1(
        i_data_bus[470]), .B2(n10410), .ZN(n8679) );
  ND2D1BWP30P140LVT U12747 ( .A1(n8680), .A2(n8679), .ZN(N14359) );
  AOI22D1BWP30P140LVT U12748 ( .A1(i_data_bus[509]), .A2(n10412), .B1(
        i_data_bus[445]), .B2(n10411), .ZN(n8682) );
  AOI22D1BWP30P140LVT U12749 ( .A1(i_data_bus[413]), .A2(n10409), .B1(
        i_data_bus[477]), .B2(n10410), .ZN(n8681) );
  ND2D1BWP30P140LVT U12750 ( .A1(n8682), .A2(n8681), .ZN(N14366) );
  AOI22D1BWP30P140LVT U12751 ( .A1(i_data_bus[404]), .A2(n10409), .B1(
        i_data_bus[500]), .B2(n10412), .ZN(n8684) );
  AOI22D1BWP30P140LVT U12752 ( .A1(i_data_bus[436]), .A2(n10411), .B1(
        i_data_bus[468]), .B2(n10410), .ZN(n8683) );
  ND2D1BWP30P140LVT U12753 ( .A1(n8684), .A2(n8683), .ZN(N14357) );
  AOI22D1BWP30P140LVT U12754 ( .A1(i_data_bus[398]), .A2(n10409), .B1(
        i_data_bus[494]), .B2(n10412), .ZN(n8686) );
  AOI22D1BWP30P140LVT U12755 ( .A1(i_data_bus[430]), .A2(n10411), .B1(
        i_data_bus[462]), .B2(n10410), .ZN(n8685) );
  ND2D1BWP30P140LVT U12756 ( .A1(n8686), .A2(n8685), .ZN(N14351) );
  AOI22D1BWP30P140LVT U12757 ( .A1(i_data_bus[506]), .A2(n10412), .B1(
        i_data_bus[442]), .B2(n10411), .ZN(n8688) );
  AOI22D1BWP30P140LVT U12758 ( .A1(i_data_bus[410]), .A2(n10409), .B1(
        i_data_bus[474]), .B2(n10410), .ZN(n8687) );
  ND2D1BWP30P140LVT U12759 ( .A1(n8688), .A2(n8687), .ZN(N14363) );
  AOI22D1BWP30P140LVT U12760 ( .A1(i_data_bus[498]), .A2(n10412), .B1(
        i_data_bus[434]), .B2(n10411), .ZN(n8690) );
  AOI22D1BWP30P140LVT U12761 ( .A1(i_data_bus[402]), .A2(n10409), .B1(
        i_data_bus[466]), .B2(n10410), .ZN(n8689) );
  ND2D1BWP30P140LVT U12762 ( .A1(n8690), .A2(n8689), .ZN(N14355) );
  AOI22D1BWP30P140LVT U12763 ( .A1(i_data_bus[850]), .A2(n10527), .B1(
        i_data_bus[818]), .B2(n10525), .ZN(n8692) );
  AOI22D1BWP30P140LVT U12764 ( .A1(i_data_bus[882]), .A2(n10526), .B1(
        i_data_bus[786]), .B2(n10528), .ZN(n8691) );
  ND2D1BWP30P140LVT U12765 ( .A1(n8692), .A2(n8691), .ZN(N7507) );
  AOI22D1BWP30P140LVT U12766 ( .A1(i_data_bus[870]), .A2(n10526), .B1(
        i_data_bus[806]), .B2(n10525), .ZN(n8694) );
  AOI22D1BWP30P140LVT U12767 ( .A1(i_data_bus[838]), .A2(n10527), .B1(
        i_data_bus[774]), .B2(n10528), .ZN(n8693) );
  ND2D1BWP30P140LVT U12768 ( .A1(n8694), .A2(n8693), .ZN(N7495) );
  AOI22D1BWP30P140LVT U12769 ( .A1(i_data_bus[853]), .A2(n10527), .B1(
        i_data_bus[821]), .B2(n10525), .ZN(n8696) );
  AOI22D1BWP30P140LVT U12770 ( .A1(i_data_bus[885]), .A2(n10526), .B1(
        i_data_bus[789]), .B2(n10528), .ZN(n8695) );
  ND2D1BWP30P140LVT U12771 ( .A1(n8696), .A2(n8695), .ZN(N7510) );
  AOI22D1BWP30P140LVT U12772 ( .A1(i_data_bus[878]), .A2(n10526), .B1(
        i_data_bus[846]), .B2(n10527), .ZN(n8698) );
  AOI22D1BWP30P140LVT U12773 ( .A1(i_data_bus[814]), .A2(n10525), .B1(
        i_data_bus[782]), .B2(n10528), .ZN(n8697) );
  ND2D1BWP30P140LVT U12774 ( .A1(n8698), .A2(n8697), .ZN(N7503) );
  AOI22D1BWP30P140LVT U12775 ( .A1(i_data_bus[836]), .A2(n10527), .B1(
        i_data_bus[804]), .B2(n10525), .ZN(n8700) );
  AOI22D1BWP30P140LVT U12776 ( .A1(i_data_bus[868]), .A2(n10526), .B1(
        i_data_bus[772]), .B2(n10528), .ZN(n8699) );
  ND2D1BWP30P140LVT U12777 ( .A1(n8700), .A2(n8699), .ZN(N7493) );
  AOI22D1BWP30P140LVT U12778 ( .A1(i_data_bus[801]), .A2(n10525), .B1(
        i_data_bus[833]), .B2(n10527), .ZN(n8702) );
  AOI22D1BWP30P140LVT U12779 ( .A1(i_data_bus[865]), .A2(n10526), .B1(
        i_data_bus[769]), .B2(n10528), .ZN(n8701) );
  ND2D1BWP30P140LVT U12780 ( .A1(n8702), .A2(n8701), .ZN(N7490) );
  AOI22D1BWP30P140LVT U12781 ( .A1(i_data_bus[828]), .A2(n10525), .B1(
        i_data_bus[892]), .B2(n10526), .ZN(n8704) );
  AOI22D1BWP30P140LVT U12782 ( .A1(i_data_bus[860]), .A2(n10527), .B1(
        i_data_bus[796]), .B2(n10528), .ZN(n8703) );
  ND2D1BWP30P140LVT U12783 ( .A1(n8704), .A2(n8703), .ZN(N7517) );
  AOI22D1BWP30P140LVT U12784 ( .A1(i_data_bus[840]), .A2(n10527), .B1(
        i_data_bus[808]), .B2(n10525), .ZN(n8706) );
  AOI22D1BWP30P140LVT U12785 ( .A1(i_data_bus[872]), .A2(n10526), .B1(
        i_data_bus[776]), .B2(n10528), .ZN(n8705) );
  ND2D1BWP30P140LVT U12786 ( .A1(n8706), .A2(n8705), .ZN(N7497) );
  AOI22D1BWP30P140LVT U12787 ( .A1(i_data_bus[800]), .A2(n10525), .B1(
        i_data_bus[864]), .B2(n10526), .ZN(n8708) );
  AOI22D1BWP30P140LVT U12788 ( .A1(i_data_bus[832]), .A2(n10527), .B1(
        i_data_bus[768]), .B2(n10528), .ZN(n8707) );
  ND2D1BWP30P140LVT U12789 ( .A1(n8708), .A2(n8707), .ZN(N7489) );
  AOI22D1BWP30P140LVT U12790 ( .A1(i_data_bus[857]), .A2(n10527), .B1(
        i_data_bus[889]), .B2(n10526), .ZN(n8710) );
  AOI22D1BWP30P140LVT U12791 ( .A1(i_data_bus[825]), .A2(n10525), .B1(
        i_data_bus[793]), .B2(n10528), .ZN(n8709) );
  ND2D1BWP30P140LVT U12792 ( .A1(n8710), .A2(n8709), .ZN(N7514) );
  AOI22D1BWP30P140LVT U12793 ( .A1(i_data_bus[873]), .A2(n10526), .B1(
        i_data_bus[809]), .B2(n10525), .ZN(n8712) );
  AOI22D1BWP30P140LVT U12794 ( .A1(i_data_bus[841]), .A2(n10527), .B1(
        i_data_bus[777]), .B2(n10528), .ZN(n8711) );
  ND2D1BWP30P140LVT U12795 ( .A1(n8712), .A2(n8711), .ZN(N7498) );
  AOI22D1BWP30P140LVT U12796 ( .A1(i_data_bus[866]), .A2(n10526), .B1(
        i_data_bus[834]), .B2(n10527), .ZN(n8714) );
  AOI22D1BWP30P140LVT U12797 ( .A1(i_data_bus[802]), .A2(n10525), .B1(
        i_data_bus[770]), .B2(n10528), .ZN(n8713) );
  ND2D1BWP30P140LVT U12798 ( .A1(n8714), .A2(n8713), .ZN(N7491) );
  AOI22D1BWP30P140LVT U12799 ( .A1(i_data_bus[605]), .A2(n10437), .B1(
        i_data_bus[541]), .B2(n10438), .ZN(n8716) );
  AOI22D1BWP30P140LVT U12800 ( .A1(i_data_bus[637]), .A2(n10440), .B1(
        i_data_bus[573]), .B2(n10439), .ZN(n8715) );
  ND2D1BWP30P140LVT U12801 ( .A1(n8716), .A2(n8715), .ZN(N12708) );
  AOI22D1BWP30P140LVT U12802 ( .A1(i_data_bus[512]), .A2(n10438), .B1(
        i_data_bus[576]), .B2(n10437), .ZN(n8718) );
  AOI22D1BWP30P140LVT U12803 ( .A1(i_data_bus[608]), .A2(n10440), .B1(
        i_data_bus[544]), .B2(n10439), .ZN(n8717) );
  ND2D1BWP30P140LVT U12804 ( .A1(n8718), .A2(n8717), .ZN(N12679) );
  AOI22D1BWP30P140LVT U12805 ( .A1(i_data_bus[513]), .A2(n10438), .B1(
        i_data_bus[577]), .B2(n10437), .ZN(n8720) );
  AOI22D1BWP30P140LVT U12806 ( .A1(i_data_bus[609]), .A2(n10440), .B1(
        i_data_bus[545]), .B2(n10439), .ZN(n8719) );
  ND2D1BWP30P140LVT U12807 ( .A1(n8720), .A2(n8719), .ZN(N12680) );
  AOI22D1BWP30P140LVT U12808 ( .A1(i_data_bus[587]), .A2(n10437), .B1(
        i_data_bus[523]), .B2(n10438), .ZN(n8722) );
  AOI22D1BWP30P140LVT U12809 ( .A1(i_data_bus[619]), .A2(n10440), .B1(
        i_data_bus[555]), .B2(n10439), .ZN(n8721) );
  ND2D1BWP30P140LVT U12810 ( .A1(n8722), .A2(n8721), .ZN(N12690) );
  AOI22D1BWP30P140LVT U12811 ( .A1(i_data_bus[597]), .A2(n10437), .B1(
        i_data_bus[629]), .B2(n10440), .ZN(n8724) );
  AOI22D1BWP30P140LVT U12812 ( .A1(i_data_bus[533]), .A2(n10438), .B1(
        i_data_bus[565]), .B2(n10439), .ZN(n8723) );
  ND2D1BWP30P140LVT U12813 ( .A1(n8724), .A2(n8723), .ZN(N12700) );
  AOI22D1BWP30P140LVT U12814 ( .A1(i_data_bus[531]), .A2(n10438), .B1(
        i_data_bus[627]), .B2(n10440), .ZN(n8726) );
  AOI22D1BWP30P140LVT U12815 ( .A1(i_data_bus[595]), .A2(n10437), .B1(
        i_data_bus[563]), .B2(n10439), .ZN(n8725) );
  ND2D1BWP30P140LVT U12816 ( .A1(n8726), .A2(n8725), .ZN(N12698) );
  AOI22D1BWP30P140LVT U12817 ( .A1(i_data_bus[612]), .A2(n10440), .B1(
        i_data_bus[580]), .B2(n10437), .ZN(n8728) );
  AOI22D1BWP30P140LVT U12818 ( .A1(i_data_bus[516]), .A2(n10438), .B1(
        i_data_bus[548]), .B2(n10439), .ZN(n8727) );
  ND2D1BWP30P140LVT U12819 ( .A1(n8728), .A2(n8727), .ZN(N12683) );
  AOI22D1BWP30P140LVT U12820 ( .A1(i_data_bus[578]), .A2(n10437), .B1(
        i_data_bus[514]), .B2(n10438), .ZN(n8730) );
  AOI22D1BWP30P140LVT U12821 ( .A1(i_data_bus[610]), .A2(n10440), .B1(
        i_data_bus[546]), .B2(n10439), .ZN(n8729) );
  ND2D1BWP30P140LVT U12822 ( .A1(n8730), .A2(n8729), .ZN(N12681) );
  AOI22D1BWP30P140LVT U12823 ( .A1(i_data_bus[600]), .A2(n10437), .B1(
        i_data_bus[632]), .B2(n10440), .ZN(n8732) );
  AOI22D1BWP30P140LVT U12824 ( .A1(i_data_bus[536]), .A2(n10438), .B1(
        i_data_bus[568]), .B2(n10439), .ZN(n8731) );
  ND2D1BWP30P140LVT U12825 ( .A1(n8732), .A2(n8731), .ZN(N12703) );
  AOI22D1BWP30P140LVT U12826 ( .A1(i_data_bus[594]), .A2(n10437), .B1(
        i_data_bus[626]), .B2(n10440), .ZN(n8734) );
  AOI22D1BWP30P140LVT U12827 ( .A1(i_data_bus[530]), .A2(n10438), .B1(
        i_data_bus[562]), .B2(n10439), .ZN(n8733) );
  ND2D1BWP30P140LVT U12828 ( .A1(n8734), .A2(n8733), .ZN(N12697) );
  AOI22D1BWP30P140LVT U12829 ( .A1(i_data_bus[631]), .A2(n10440), .B1(
        i_data_bus[535]), .B2(n10438), .ZN(n8736) );
  AOI22D1BWP30P140LVT U12830 ( .A1(i_data_bus[599]), .A2(n10437), .B1(
        i_data_bus[567]), .B2(n10439), .ZN(n8735) );
  ND2D1BWP30P140LVT U12831 ( .A1(n8736), .A2(n8735), .ZN(N12702) );
  AOI22D1BWP30P140LVT U12832 ( .A1(i_data_bus[687]), .A2(n10593), .B1(
        i_data_bus[751]), .B2(n10595), .ZN(n8738) );
  AOI22D1BWP30P140LVT U12833 ( .A1(i_data_bus[719]), .A2(n10594), .B1(
        i_data_bus[655]), .B2(n10596), .ZN(n8737) );
  ND2D1BWP30P140LVT U12834 ( .A1(n8738), .A2(n8737), .ZN(N3540) );
  AOI22D1BWP30P140LVT U12835 ( .A1(i_data_bus[703]), .A2(n10593), .B1(
        i_data_bus[767]), .B2(n10595), .ZN(n8740) );
  AOI22D1BWP30P140LVT U12836 ( .A1(i_data_bus[735]), .A2(n10594), .B1(
        i_data_bus[671]), .B2(n10596), .ZN(n8739) );
  ND2D1BWP30P140LVT U12837 ( .A1(n8740), .A2(n8739), .ZN(N3556) );
  AOI22D1BWP30P140LVT U12838 ( .A1(i_data_bus[752]), .A2(n10595), .B1(
        i_data_bus[720]), .B2(n10594), .ZN(n8742) );
  AOI22D1BWP30P140LVT U12839 ( .A1(i_data_bus[688]), .A2(n10593), .B1(
        i_data_bus[656]), .B2(n10596), .ZN(n8741) );
  ND2D1BWP30P140LVT U12840 ( .A1(n8742), .A2(n8741), .ZN(N3541) );
  AOI22D1BWP30P140LVT U12841 ( .A1(i_data_bus[714]), .A2(n10594), .B1(
        i_data_bus[682]), .B2(n10593), .ZN(n8744) );
  AOI22D1BWP30P140LVT U12842 ( .A1(i_data_bus[746]), .A2(n10595), .B1(
        i_data_bus[650]), .B2(n10596), .ZN(n8743) );
  ND2D1BWP30P140LVT U12843 ( .A1(n8744), .A2(n8743), .ZN(N3535) );
  AOI22D1BWP30P140LVT U12844 ( .A1(i_data_bus[716]), .A2(n10594), .B1(
        i_data_bus[748]), .B2(n10595), .ZN(n8746) );
  AOI22D1BWP30P140LVT U12845 ( .A1(i_data_bus[684]), .A2(n10593), .B1(
        i_data_bus[652]), .B2(n10596), .ZN(n8745) );
  ND2D1BWP30P140LVT U12846 ( .A1(n8746), .A2(n8745), .ZN(N3537) );
  AOI22D1BWP30P140LVT U12847 ( .A1(i_data_bus[694]), .A2(n10593), .B1(
        i_data_bus[726]), .B2(n10594), .ZN(n8748) );
  AOI22D1BWP30P140LVT U12848 ( .A1(i_data_bus[758]), .A2(n10595), .B1(
        i_data_bus[662]), .B2(n10596), .ZN(n8747) );
  ND2D1BWP30P140LVT U12849 ( .A1(n8748), .A2(n8747), .ZN(N3547) );
  AOI22D1BWP30P140LVT U12850 ( .A1(i_data_bus[732]), .A2(n10594), .B1(
        i_data_bus[700]), .B2(n10593), .ZN(n8750) );
  AOI22D1BWP30P140LVT U12851 ( .A1(i_data_bus[764]), .A2(n10595), .B1(
        i_data_bus[668]), .B2(n10596), .ZN(n8749) );
  ND2D1BWP30P140LVT U12852 ( .A1(n8750), .A2(n8749), .ZN(N3553) );
  AOI22D1BWP30P140LVT U12853 ( .A1(i_data_bus[681]), .A2(n10593), .B1(
        i_data_bus[745]), .B2(n10595), .ZN(n8752) );
  AOI22D1BWP30P140LVT U12854 ( .A1(i_data_bus[713]), .A2(n10594), .B1(
        i_data_bus[649]), .B2(n10596), .ZN(n8751) );
  ND2D1BWP30P140LVT U12855 ( .A1(n8752), .A2(n8751), .ZN(N3534) );
  AOI22D1BWP30P140LVT U12856 ( .A1(i_data_bus[708]), .A2(n10594), .B1(
        i_data_bus[676]), .B2(n10593), .ZN(n8754) );
  AOI22D1BWP30P140LVT U12857 ( .A1(i_data_bus[740]), .A2(n10595), .B1(
        i_data_bus[644]), .B2(n10596), .ZN(n8753) );
  ND2D1BWP30P140LVT U12858 ( .A1(n8754), .A2(n8753), .ZN(N3529) );
  AOI22D1BWP30P140LVT U12859 ( .A1(i_data_bus[611]), .A2(n10470), .B1(
        i_data_bus[515]), .B2(n10471), .ZN(n8756) );
  AOI22D1BWP30P140LVT U12860 ( .A1(i_data_bus[579]), .A2(n10469), .B1(
        i_data_bus[547]), .B2(n10472), .ZN(n8755) );
  ND2D1BWP30P140LVT U12861 ( .A1(n8756), .A2(n8755), .ZN(N10808) );
  AOI22D1BWP30P140LVT U12862 ( .A1(i_data_bus[599]), .A2(n10469), .B1(
        i_data_bus[631]), .B2(n10470), .ZN(n8758) );
  AOI22D1BWP30P140LVT U12863 ( .A1(i_data_bus[535]), .A2(n10471), .B1(
        i_data_bus[567]), .B2(n10472), .ZN(n8757) );
  ND2D1BWP30P140LVT U12864 ( .A1(n8758), .A2(n8757), .ZN(N10828) );
  AOI22D1BWP30P140LVT U12865 ( .A1(i_data_bus[531]), .A2(n10471), .B1(
        i_data_bus[595]), .B2(n10469), .ZN(n8760) );
  AOI22D1BWP30P140LVT U12866 ( .A1(i_data_bus[627]), .A2(n10470), .B1(
        i_data_bus[563]), .B2(n10472), .ZN(n8759) );
  ND2D1BWP30P140LVT U12867 ( .A1(n8760), .A2(n8759), .ZN(N10824) );
  AOI22D1BWP30P140LVT U12868 ( .A1(i_data_bus[513]), .A2(n10471), .B1(
        i_data_bus[577]), .B2(n10469), .ZN(n8762) );
  AOI22D1BWP30P140LVT U12869 ( .A1(i_data_bus[609]), .A2(n10470), .B1(
        i_data_bus[545]), .B2(n10472), .ZN(n8761) );
  ND2D1BWP30P140LVT U12870 ( .A1(n8762), .A2(n8761), .ZN(N10806) );
  AOI22D1BWP30P140LVT U12871 ( .A1(i_data_bus[608]), .A2(n10470), .B1(
        i_data_bus[576]), .B2(n10469), .ZN(n8764) );
  AOI22D1BWP30P140LVT U12872 ( .A1(i_data_bus[512]), .A2(n10471), .B1(
        i_data_bus[544]), .B2(n10472), .ZN(n8763) );
  ND2D1BWP30P140LVT U12873 ( .A1(n8764), .A2(n8763), .ZN(N10805) );
  AOI22D1BWP30P140LVT U12874 ( .A1(i_data_bus[578]), .A2(n10469), .B1(
        i_data_bus[514]), .B2(n10471), .ZN(n8766) );
  AOI22D1BWP30P140LVT U12875 ( .A1(i_data_bus[610]), .A2(n10470), .B1(
        i_data_bus[546]), .B2(n10472), .ZN(n8765) );
  ND2D1BWP30P140LVT U12876 ( .A1(n8766), .A2(n8765), .ZN(N10807) );
  AOI22D1BWP30P140LVT U12877 ( .A1(i_data_bus[533]), .A2(n10471), .B1(
        i_data_bus[629]), .B2(n10470), .ZN(n8768) );
  AOI22D1BWP30P140LVT U12878 ( .A1(i_data_bus[597]), .A2(n10469), .B1(
        i_data_bus[565]), .B2(n10472), .ZN(n8767) );
  ND2D1BWP30P140LVT U12879 ( .A1(n8768), .A2(n8767), .ZN(N10826) );
  AOI22D1BWP30P140LVT U12880 ( .A1(i_data_bus[634]), .A2(n10470), .B1(
        i_data_bus[538]), .B2(n10471), .ZN(n8770) );
  AOI22D1BWP30P140LVT U12881 ( .A1(i_data_bus[602]), .A2(n10469), .B1(
        i_data_bus[570]), .B2(n10472), .ZN(n8769) );
  ND2D1BWP30P140LVT U12882 ( .A1(n8770), .A2(n8769), .ZN(N10831) );
  AOI22D1BWP30P140LVT U12883 ( .A1(i_data_bus[521]), .A2(n10471), .B1(
        i_data_bus[585]), .B2(n10469), .ZN(n8772) );
  AOI22D1BWP30P140LVT U12884 ( .A1(i_data_bus[617]), .A2(n10470), .B1(
        i_data_bus[553]), .B2(n10472), .ZN(n8771) );
  ND2D1BWP30P140LVT U12885 ( .A1(n8772), .A2(n8771), .ZN(N10814) );
  AOI22D1BWP30P140LVT U12886 ( .A1(i_data_bus[802]), .A2(n10430), .B1(
        i_data_bus[770]), .B2(n10429), .ZN(n8774) );
  AOI22D1BWP30P140LVT U12887 ( .A1(i_data_bus[866]), .A2(n10431), .B1(
        i_data_bus[834]), .B2(n10432), .ZN(n8773) );
  ND2D1BWP30P140LVT U12888 ( .A1(n8774), .A2(n8773), .ZN(N13113) );
  AOI22D1BWP30P140LVT U12889 ( .A1(i_data_bus[827]), .A2(n10430), .B1(
        i_data_bus[891]), .B2(n10431), .ZN(n8776) );
  AOI22D1BWP30P140LVT U12890 ( .A1(i_data_bus[795]), .A2(n10429), .B1(
        i_data_bus[859]), .B2(n10432), .ZN(n8775) );
  ND2D1BWP30P140LVT U12891 ( .A1(n8776), .A2(n8775), .ZN(N13138) );
  AOI22D1BWP30P140LVT U12892 ( .A1(i_data_bus[869]), .A2(n10431), .B1(
        i_data_bus[773]), .B2(n10429), .ZN(n8778) );
  AOI22D1BWP30P140LVT U12893 ( .A1(i_data_bus[805]), .A2(n10430), .B1(
        i_data_bus[837]), .B2(n10432), .ZN(n8777) );
  ND2D1BWP30P140LVT U12894 ( .A1(n8778), .A2(n8777), .ZN(N13116) );
  AOI22D1BWP30P140LVT U12895 ( .A1(i_data_bus[783]), .A2(n10429), .B1(
        i_data_bus[815]), .B2(n10430), .ZN(n8780) );
  AOI22D1BWP30P140LVT U12896 ( .A1(i_data_bus[879]), .A2(n10431), .B1(
        i_data_bus[847]), .B2(n10432), .ZN(n8779) );
  ND2D1BWP30P140LVT U12897 ( .A1(n8780), .A2(n8779), .ZN(N13126) );
  AOI22D1BWP30P140LVT U12898 ( .A1(i_data_bus[251]), .A2(n10484), .B1(
        i_data_bus[219]), .B2(n10482), .ZN(n8782) );
  AOI22D1BWP30P140LVT U12899 ( .A1(i_data_bus[187]), .A2(n10483), .B1(
        i_data_bus[155]), .B2(n10481), .ZN(n8781) );
  ND2D1BWP30P140LVT U12900 ( .A1(n8782), .A2(n8781), .ZN(N10184) );
  AOI22D1BWP30P140LVT U12901 ( .A1(i_data_bus[174]), .A2(n10483), .B1(
        i_data_bus[238]), .B2(n10484), .ZN(n8784) );
  AOI22D1BWP30P140LVT U12902 ( .A1(i_data_bus[206]), .A2(n10482), .B1(
        i_data_bus[142]), .B2(n10481), .ZN(n8783) );
  ND2D1BWP30P140LVT U12903 ( .A1(n8784), .A2(n8783), .ZN(N10171) );
  AOI22D1BWP30P140LVT U12904 ( .A1(i_data_bus[168]), .A2(n10483), .B1(
        i_data_bus[232]), .B2(n10484), .ZN(n8786) );
  AOI22D1BWP30P140LVT U12905 ( .A1(i_data_bus[200]), .A2(n10482), .B1(
        i_data_bus[136]), .B2(n10481), .ZN(n8785) );
  ND2D1BWP30P140LVT U12906 ( .A1(n8786), .A2(n8785), .ZN(N10165) );
  AOI22D1BWP30P140LVT U12907 ( .A1(i_data_bus[231]), .A2(n10484), .B1(
        i_data_bus[167]), .B2(n10483), .ZN(n8788) );
  AOI22D1BWP30P140LVT U12908 ( .A1(i_data_bus[199]), .A2(n10482), .B1(
        i_data_bus[135]), .B2(n10481), .ZN(n8787) );
  ND2D1BWP30P140LVT U12909 ( .A1(n8788), .A2(n8787), .ZN(N10164) );
  AOI22D1BWP30P140LVT U12910 ( .A1(i_data_bus[222]), .A2(n10482), .B1(
        i_data_bus[254]), .B2(n10484), .ZN(n8790) );
  AOI22D1BWP30P140LVT U12911 ( .A1(i_data_bus[190]), .A2(n10483), .B1(
        i_data_bus[158]), .B2(n10481), .ZN(n8789) );
  ND2D1BWP30P140LVT U12912 ( .A1(n8790), .A2(n8789), .ZN(N10187) );
  AOI22D1BWP30P140LVT U12913 ( .A1(i_data_bus[194]), .A2(n10482), .B1(
        i_data_bus[226]), .B2(n10484), .ZN(n8792) );
  AOI22D1BWP30P140LVT U12914 ( .A1(i_data_bus[162]), .A2(n10483), .B1(
        i_data_bus[130]), .B2(n10481), .ZN(n8791) );
  ND2D1BWP30P140LVT U12915 ( .A1(n8792), .A2(n8791), .ZN(N10159) );
  AOI22D1BWP30P140LVT U12916 ( .A1(i_data_bus[249]), .A2(n10484), .B1(
        i_data_bus[185]), .B2(n10483), .ZN(n8794) );
  AOI22D1BWP30P140LVT U12917 ( .A1(i_data_bus[217]), .A2(n10482), .B1(
        i_data_bus[153]), .B2(n10481), .ZN(n8793) );
  ND2D1BWP30P140LVT U12918 ( .A1(n8794), .A2(n8793), .ZN(N10182) );
  AOI22D1BWP30P140LVT U12919 ( .A1(i_data_bus[248]), .A2(n10484), .B1(
        i_data_bus[216]), .B2(n10482), .ZN(n8796) );
  AOI22D1BWP30P140LVT U12920 ( .A1(i_data_bus[184]), .A2(n10483), .B1(
        i_data_bus[152]), .B2(n10481), .ZN(n8795) );
  ND2D1BWP30P140LVT U12921 ( .A1(n8796), .A2(n8795), .ZN(N10181) );
  AOI22D1BWP30P140LVT U12922 ( .A1(i_data_bus[210]), .A2(n10482), .B1(
        i_data_bus[242]), .B2(n10484), .ZN(n8798) );
  AOI22D1BWP30P140LVT U12923 ( .A1(i_data_bus[178]), .A2(n10483), .B1(
        i_data_bus[146]), .B2(n10481), .ZN(n8797) );
  ND2D1BWP30P140LVT U12924 ( .A1(n8798), .A2(n8797), .ZN(N10175) );
  AOI22D1BWP30P140LVT U12925 ( .A1(i_data_bus[170]), .A2(n10483), .B1(
        i_data_bus[202]), .B2(n10482), .ZN(n8800) );
  AOI22D1BWP30P140LVT U12926 ( .A1(i_data_bus[234]), .A2(n10484), .B1(
        i_data_bus[138]), .B2(n10481), .ZN(n8799) );
  ND2D1BWP30P140LVT U12927 ( .A1(n8800), .A2(n8799), .ZN(N10167) );
  AOI22D1BWP30P140LVT U12928 ( .A1(i_data_bus[201]), .A2(n10482), .B1(
        i_data_bus[169]), .B2(n10483), .ZN(n8802) );
  AOI22D1BWP30P140LVT U12929 ( .A1(i_data_bus[233]), .A2(n10484), .B1(
        i_data_bus[137]), .B2(n10481), .ZN(n8801) );
  ND2D1BWP30P140LVT U12930 ( .A1(n8802), .A2(n8801), .ZN(N10166) );
  AOI22D1BWP30P140LVT U12931 ( .A1(i_data_bus[54]), .A2(n10453), .B1(
        i_data_bus[22]), .B2(n10456), .ZN(n8804) );
  AOI22D1BWP30P140LVT U12932 ( .A1(i_data_bus[118]), .A2(n10455), .B1(
        i_data_bus[86]), .B2(n10454), .ZN(n8803) );
  ND2D1BWP30P140LVT U12933 ( .A1(n8804), .A2(n8803), .ZN(N11837) );
  AOI22D1BWP30P140LVT U12934 ( .A1(i_data_bus[116]), .A2(n10455), .B1(
        i_data_bus[20]), .B2(n10456), .ZN(n8806) );
  AOI22D1BWP30P140LVT U12935 ( .A1(i_data_bus[52]), .A2(n10453), .B1(
        i_data_bus[84]), .B2(n10454), .ZN(n8805) );
  ND2D1BWP30P140LVT U12936 ( .A1(n8806), .A2(n8805), .ZN(N11835) );
  AOI22D1BWP30P140LVT U12937 ( .A1(i_data_bus[14]), .A2(n10456), .B1(
        i_data_bus[110]), .B2(n10455), .ZN(n8808) );
  AOI22D1BWP30P140LVT U12938 ( .A1(i_data_bus[46]), .A2(n10453), .B1(
        i_data_bus[78]), .B2(n10454), .ZN(n8807) );
  ND2D1BWP30P140LVT U12939 ( .A1(n8808), .A2(n8807), .ZN(N11829) );
  AOI22D1BWP30P140LVT U12940 ( .A1(i_data_bus[120]), .A2(n10455), .B1(
        i_data_bus[56]), .B2(n10453), .ZN(n8810) );
  AOI22D1BWP30P140LVT U12941 ( .A1(i_data_bus[24]), .A2(n10456), .B1(
        i_data_bus[88]), .B2(n10454), .ZN(n8809) );
  ND2D1BWP30P140LVT U12942 ( .A1(n8810), .A2(n8809), .ZN(N11839) );
  AOI22D1BWP30P140LVT U12943 ( .A1(i_data_bus[59]), .A2(n10453), .B1(
        i_data_bus[27]), .B2(n10456), .ZN(n8812) );
  AOI22D1BWP30P140LVT U12944 ( .A1(i_data_bus[123]), .A2(n10455), .B1(
        i_data_bus[91]), .B2(n10454), .ZN(n8811) );
  ND2D1BWP30P140LVT U12945 ( .A1(n8812), .A2(n8811), .ZN(N11842) );
  AOI22D1BWP30P140LVT U12946 ( .A1(i_data_bus[45]), .A2(n10453), .B1(
        i_data_bus[13]), .B2(n10456), .ZN(n8814) );
  AOI22D1BWP30P140LVT U12947 ( .A1(i_data_bus[109]), .A2(n10455), .B1(
        i_data_bus[77]), .B2(n10454), .ZN(n8813) );
  ND2D1BWP30P140LVT U12948 ( .A1(n8814), .A2(n8813), .ZN(N11828) );
  AOI22D1BWP30P140LVT U12949 ( .A1(i_data_bus[462]), .A2(n10538), .B1(
        i_data_bus[494]), .B2(n10539), .ZN(n8816) );
  AOI22D1BWP30P140LVT U12950 ( .A1(i_data_bus[398]), .A2(n10537), .B1(
        i_data_bus[430]), .B2(n10540), .ZN(n8815) );
  ND2D1BWP30P140LVT U12951 ( .A1(n8816), .A2(n8815), .ZN(N6855) );
  AOI22D1BWP30P140LVT U12952 ( .A1(i_data_bus[402]), .A2(n10537), .B1(
        i_data_bus[466]), .B2(n10538), .ZN(n8818) );
  AOI22D1BWP30P140LVT U12953 ( .A1(i_data_bus[498]), .A2(n10539), .B1(
        i_data_bus[434]), .B2(n10540), .ZN(n8817) );
  ND2D1BWP30P140LVT U12954 ( .A1(n8818), .A2(n8817), .ZN(N6859) );
  AOI22D1BWP30P140LVT U12955 ( .A1(i_data_bus[413]), .A2(n10537), .B1(
        i_data_bus[477]), .B2(n10538), .ZN(n8820) );
  AOI22D1BWP30P140LVT U12956 ( .A1(i_data_bus[509]), .A2(n10539), .B1(
        i_data_bus[445]), .B2(n10540), .ZN(n8819) );
  ND2D1BWP30P140LVT U12957 ( .A1(n8820), .A2(n8819), .ZN(N6870) );
  AOI22D1BWP30P140LVT U12958 ( .A1(i_data_bus[469]), .A2(n10538), .B1(
        i_data_bus[501]), .B2(n10539), .ZN(n8822) );
  AOI22D1BWP30P140LVT U12959 ( .A1(i_data_bus[405]), .A2(n10537), .B1(
        i_data_bus[437]), .B2(n10540), .ZN(n8821) );
  ND2D1BWP30P140LVT U12960 ( .A1(n8822), .A2(n8821), .ZN(N6862) );
  AOI22D1BWP30P140LVT U12961 ( .A1(i_data_bus[481]), .A2(n10539), .B1(
        i_data_bus[449]), .B2(n10538), .ZN(n8824) );
  AOI22D1BWP30P140LVT U12962 ( .A1(i_data_bus[385]), .A2(n10537), .B1(
        i_data_bus[417]), .B2(n10540), .ZN(n8823) );
  ND2D1BWP30P140LVT U12963 ( .A1(n8824), .A2(n8823), .ZN(N6842) );
  AOI22D1BWP30P140LVT U12964 ( .A1(i_data_bus[455]), .A2(n10538), .B1(
        i_data_bus[487]), .B2(n10539), .ZN(n8826) );
  AOI22D1BWP30P140LVT U12965 ( .A1(i_data_bus[391]), .A2(n10537), .B1(
        i_data_bus[423]), .B2(n10540), .ZN(n8825) );
  ND2D1BWP30P140LVT U12966 ( .A1(n8826), .A2(n8825), .ZN(N6848) );
  AOI22D1BWP30P140LVT U12967 ( .A1(i_data_bus[489]), .A2(n10539), .B1(
        i_data_bus[393]), .B2(n10537), .ZN(n8828) );
  AOI22D1BWP30P140LVT U12968 ( .A1(i_data_bus[457]), .A2(n10538), .B1(
        i_data_bus[425]), .B2(n10540), .ZN(n8827) );
  ND2D1BWP30P140LVT U12969 ( .A1(n8828), .A2(n8827), .ZN(N6850) );
  AOI22D1BWP30P140LVT U12970 ( .A1(i_data_bus[485]), .A2(n10539), .B1(
        i_data_bus[453]), .B2(n10538), .ZN(n8830) );
  AOI22D1BWP30P140LVT U12971 ( .A1(i_data_bus[389]), .A2(n10537), .B1(
        i_data_bus[421]), .B2(n10540), .ZN(n8829) );
  ND2D1BWP30P140LVT U12972 ( .A1(n8830), .A2(n8829), .ZN(N6846) );
  AOI22D1BWP30P140LVT U12973 ( .A1(i_data_bus[458]), .A2(n10538), .B1(
        i_data_bus[394]), .B2(n10537), .ZN(n8832) );
  AOI22D1BWP30P140LVT U12974 ( .A1(i_data_bus[490]), .A2(n10539), .B1(
        i_data_bus[426]), .B2(n10540), .ZN(n8831) );
  ND2D1BWP30P140LVT U12975 ( .A1(n8832), .A2(n8831), .ZN(N6851) );
  AOI22D1BWP30P140LVT U12976 ( .A1(i_data_bus[488]), .A2(n10539), .B1(
        i_data_bus[392]), .B2(n10537), .ZN(n8834) );
  AOI22D1BWP30P140LVT U12977 ( .A1(i_data_bus[456]), .A2(n10538), .B1(
        i_data_bus[424]), .B2(n10540), .ZN(n8833) );
  ND2D1BWP30P140LVT U12978 ( .A1(n8834), .A2(n8833), .ZN(N6849) );
  AOI22D1BWP30P140LVT U12979 ( .A1(i_data_bus[829]), .A2(n10560), .B1(
        i_data_bus[861]), .B2(n10557), .ZN(n8836) );
  AOI22D1BWP30P140LVT U12980 ( .A1(i_data_bus[893]), .A2(n10559), .B1(
        i_data_bus[797]), .B2(n10558), .ZN(n8835) );
  ND2D1BWP30P140LVT U12981 ( .A1(n8836), .A2(n8835), .ZN(N5644) );
  AOI22D1BWP30P140LVT U12982 ( .A1(i_data_bus[855]), .A2(n10557), .B1(
        i_data_bus[887]), .B2(n10559), .ZN(n8838) );
  AOI22D1BWP30P140LVT U12983 ( .A1(i_data_bus[823]), .A2(n10560), .B1(
        i_data_bus[791]), .B2(n10558), .ZN(n8837) );
  ND2D1BWP30P140LVT U12984 ( .A1(n8838), .A2(n8837), .ZN(N5638) );
  AOI22D1BWP30P140LVT U12985 ( .A1(i_data_bus[807]), .A2(n10560), .B1(
        i_data_bus[839]), .B2(n10557), .ZN(n8840) );
  AOI22D1BWP30P140LVT U12986 ( .A1(i_data_bus[871]), .A2(n10559), .B1(
        i_data_bus[775]), .B2(n10558), .ZN(n8839) );
  ND2D1BWP30P140LVT U12987 ( .A1(n8840), .A2(n8839), .ZN(N5622) );
  AOI22D1BWP30P140LVT U12988 ( .A1(i_data_bus[850]), .A2(n10557), .B1(
        i_data_bus[818]), .B2(n10560), .ZN(n8842) );
  AOI22D1BWP30P140LVT U12989 ( .A1(i_data_bus[882]), .A2(n10559), .B1(
        i_data_bus[786]), .B2(n10558), .ZN(n8841) );
  ND2D1BWP30P140LVT U12990 ( .A1(n8842), .A2(n8841), .ZN(N5633) );
  AOI22D1BWP30P140LVT U12991 ( .A1(i_data_bus[873]), .A2(n10559), .B1(
        i_data_bus[809]), .B2(n10560), .ZN(n8844) );
  AOI22D1BWP30P140LVT U12992 ( .A1(i_data_bus[841]), .A2(n10557), .B1(
        i_data_bus[777]), .B2(n10558), .ZN(n8843) );
  ND2D1BWP30P140LVT U12993 ( .A1(n8844), .A2(n8843), .ZN(N5624) );
  AOI22D1BWP30P140LVT U12994 ( .A1(i_data_bus[888]), .A2(n10559), .B1(
        i_data_bus[824]), .B2(n10560), .ZN(n8846) );
  AOI22D1BWP30P140LVT U12995 ( .A1(i_data_bus[856]), .A2(n10557), .B1(
        i_data_bus[792]), .B2(n10558), .ZN(n8845) );
  ND2D1BWP30P140LVT U12996 ( .A1(n8846), .A2(n8845), .ZN(N5639) );
  AOI22D1BWP30P140LVT U12997 ( .A1(i_data_bus[884]), .A2(n10559), .B1(
        i_data_bus[852]), .B2(n10557), .ZN(n8848) );
  AOI22D1BWP30P140LVT U12998 ( .A1(i_data_bus[820]), .A2(n10560), .B1(
        i_data_bus[788]), .B2(n10558), .ZN(n8847) );
  ND2D1BWP30P140LVT U12999 ( .A1(n8848), .A2(n8847), .ZN(N5635) );
  AOI22D1BWP30P140LVT U13000 ( .A1(i_data_bus[996]), .A2(n10556), .B1(
        i_data_bus[900]), .B2(n10554), .ZN(n8850) );
  AOI22D1BWP30P140LVT U13001 ( .A1(i_data_bus[932]), .A2(n10553), .B1(
        i_data_bus[964]), .B2(n10555), .ZN(n8849) );
  ND2D1BWP30P140LVT U13002 ( .A1(n8850), .A2(n8849), .ZN(N5835) );
  AOI22D1BWP30P140LVT U13003 ( .A1(i_data_bus[952]), .A2(n10553), .B1(
        i_data_bus[920]), .B2(n10554), .ZN(n8852) );
  AOI22D1BWP30P140LVT U13004 ( .A1(i_data_bus[1016]), .A2(n10556), .B1(
        i_data_bus[984]), .B2(n10555), .ZN(n8851) );
  ND2D1BWP30P140LVT U13005 ( .A1(n8852), .A2(n8851), .ZN(N5855) );
  AOI22D1BWP30P140LVT U13006 ( .A1(i_data_bus[940]), .A2(n10553), .B1(
        i_data_bus[1004]), .B2(n10556), .ZN(n8854) );
  AOI22D1BWP30P140LVT U13007 ( .A1(i_data_bus[908]), .A2(n10554), .B1(
        i_data_bus[972]), .B2(n10555), .ZN(n8853) );
  ND2D1BWP30P140LVT U13008 ( .A1(n8854), .A2(n8853), .ZN(N5843) );
  AOI22D1BWP30P140LVT U13009 ( .A1(i_data_bus[896]), .A2(n10554), .B1(
        i_data_bus[928]), .B2(n10553), .ZN(n8856) );
  AOI22D1BWP30P140LVT U13010 ( .A1(i_data_bus[992]), .A2(n10556), .B1(
        i_data_bus[960]), .B2(n10555), .ZN(n8855) );
  ND2D1BWP30P140LVT U13011 ( .A1(n8856), .A2(n8855), .ZN(N5831) );
  AOI22D1BWP30P140LVT U13012 ( .A1(i_data_bus[910]), .A2(n10554), .B1(
        i_data_bus[942]), .B2(n10553), .ZN(n8858) );
  AOI22D1BWP30P140LVT U13013 ( .A1(i_data_bus[1006]), .A2(n10556), .B1(
        i_data_bus[974]), .B2(n10555), .ZN(n8857) );
  ND2D1BWP30P140LVT U13014 ( .A1(n8858), .A2(n8857), .ZN(N5845) );
  AOI22D1BWP30P140LVT U13015 ( .A1(i_data_bus[926]), .A2(n10554), .B1(
        i_data_bus[1022]), .B2(n10556), .ZN(n8860) );
  AOI22D1BWP30P140LVT U13016 ( .A1(i_data_bus[958]), .A2(n10553), .B1(
        i_data_bus[990]), .B2(n10555), .ZN(n8859) );
  ND2D1BWP30P140LVT U13017 ( .A1(n8860), .A2(n8859), .ZN(N5861) );
  AOI22D1BWP30P140LVT U13018 ( .A1(i_data_bus[947]), .A2(n10553), .B1(
        i_data_bus[915]), .B2(n10554), .ZN(n8862) );
  AOI22D1BWP30P140LVT U13019 ( .A1(i_data_bus[1011]), .A2(n10556), .B1(
        i_data_bus[979]), .B2(n10555), .ZN(n8861) );
  ND2D1BWP30P140LVT U13020 ( .A1(n8862), .A2(n8861), .ZN(N5850) );
  AOI22D1BWP30P140LVT U13021 ( .A1(i_data_bus[1016]), .A2(n10523), .B1(
        i_data_bus[984]), .B2(n10522), .ZN(n8864) );
  AOI22D1BWP30P140LVT U13022 ( .A1(i_data_bus[952]), .A2(n10521), .B1(
        i_data_bus[920]), .B2(n10524), .ZN(n8863) );
  ND2D1BWP30P140LVT U13023 ( .A1(n8864), .A2(n8863), .ZN(N7729) );
  AOI22D1BWP30P140LVT U13024 ( .A1(i_data_bus[1014]), .A2(n10523), .B1(
        i_data_bus[982]), .B2(n10522), .ZN(n8866) );
  AOI22D1BWP30P140LVT U13025 ( .A1(i_data_bus[950]), .A2(n10521), .B1(
        i_data_bus[918]), .B2(n10524), .ZN(n8865) );
  ND2D1BWP30P140LVT U13026 ( .A1(n8866), .A2(n8865), .ZN(N7727) );
  AOI22D1BWP30P140LVT U13027 ( .A1(i_data_bus[978]), .A2(n10522), .B1(
        i_data_bus[1010]), .B2(n10523), .ZN(n8868) );
  AOI22D1BWP30P140LVT U13028 ( .A1(i_data_bus[946]), .A2(n10521), .B1(
        i_data_bus[914]), .B2(n10524), .ZN(n8867) );
  ND2D1BWP30P140LVT U13029 ( .A1(n8868), .A2(n8867), .ZN(N7723) );
  AOI22D1BWP30P140LVT U13030 ( .A1(i_data_bus[998]), .A2(n10523), .B1(
        i_data_bus[966]), .B2(n10522), .ZN(n8870) );
  AOI22D1BWP30P140LVT U13031 ( .A1(i_data_bus[934]), .A2(n10521), .B1(
        i_data_bus[902]), .B2(n10524), .ZN(n8869) );
  ND2D1BWP30P140LVT U13032 ( .A1(n8870), .A2(n8869), .ZN(N7711) );
  AOI22D1BWP30P140LVT U13033 ( .A1(i_data_bus[945]), .A2(n10521), .B1(
        i_data_bus[977]), .B2(n10522), .ZN(n8872) );
  AOI22D1BWP30P140LVT U13034 ( .A1(i_data_bus[1009]), .A2(n10523), .B1(
        i_data_bus[913]), .B2(n10524), .ZN(n8871) );
  ND2D1BWP30P140LVT U13035 ( .A1(n8872), .A2(n8871), .ZN(N7722) );
  AOI22D1BWP30P140LVT U13036 ( .A1(i_data_bus[222]), .A2(n10578), .B1(
        i_data_bus[158]), .B2(n10577), .ZN(n8874) );
  AOI22D1BWP30P140LVT U13037 ( .A1(i_data_bus[190]), .A2(n10579), .B1(
        i_data_bus[254]), .B2(n10580), .ZN(n8873) );
  ND2D1BWP30P140LVT U13038 ( .A1(n8874), .A2(n8873), .ZN(N4565) );
  AOI22D1BWP30P140LVT U13039 ( .A1(i_data_bus[147]), .A2(n10577), .B1(
        i_data_bus[211]), .B2(n10578), .ZN(n8876) );
  AOI22D1BWP30P140LVT U13040 ( .A1(i_data_bus[179]), .A2(n10579), .B1(
        i_data_bus[243]), .B2(n10580), .ZN(n8875) );
  ND2D1BWP30P140LVT U13041 ( .A1(n8876), .A2(n8875), .ZN(N4554) );
  AOI22D1BWP30P140LVT U13042 ( .A1(i_data_bus[165]), .A2(n10579), .B1(
        i_data_bus[197]), .B2(n10578), .ZN(n8878) );
  AOI22D1BWP30P140LVT U13043 ( .A1(i_data_bus[133]), .A2(n10577), .B1(
        i_data_bus[229]), .B2(n10580), .ZN(n8877) );
  ND2D1BWP30P140LVT U13044 ( .A1(n8878), .A2(n8877), .ZN(N4540) );
  AOI22D1BWP30P140LVT U13045 ( .A1(i_data_bus[144]), .A2(n10577), .B1(
        i_data_bus[208]), .B2(n10578), .ZN(n8880) );
  AOI22D1BWP30P140LVT U13046 ( .A1(i_data_bus[176]), .A2(n10579), .B1(
        i_data_bus[240]), .B2(n10580), .ZN(n8879) );
  ND2D1BWP30P140LVT U13047 ( .A1(n8880), .A2(n8879), .ZN(N4551) );
  AOI22D1BWP30P140LVT U13048 ( .A1(i_data_bus[161]), .A2(n10579), .B1(
        i_data_bus[129]), .B2(n10577), .ZN(n8882) );
  AOI22D1BWP30P140LVT U13049 ( .A1(i_data_bus[193]), .A2(n10578), .B1(
        i_data_bus[225]), .B2(n10580), .ZN(n8881) );
  ND2D1BWP30P140LVT U13050 ( .A1(n8882), .A2(n8881), .ZN(N4536) );
  AOI22D1BWP30P140LVT U13051 ( .A1(i_data_bus[178]), .A2(n10579), .B1(
        i_data_bus[210]), .B2(n10578), .ZN(n8884) );
  AOI22D1BWP30P140LVT U13052 ( .A1(i_data_bus[146]), .A2(n10577), .B1(
        i_data_bus[242]), .B2(n10580), .ZN(n8883) );
  ND2D1BWP30P140LVT U13053 ( .A1(n8884), .A2(n8883), .ZN(N4553) );
  AOI22D1BWP30P140LVT U13054 ( .A1(i_data_bus[205]), .A2(n10578), .B1(
        i_data_bus[141]), .B2(n10577), .ZN(n8886) );
  AOI22D1BWP30P140LVT U13055 ( .A1(i_data_bus[173]), .A2(n10579), .B1(
        i_data_bus[237]), .B2(n10580), .ZN(n8885) );
  ND2D1BWP30P140LVT U13056 ( .A1(n8886), .A2(n8885), .ZN(N4548) );
  AOI22D1BWP30P140LVT U13057 ( .A1(i_data_bus[220]), .A2(n10578), .B1(
        i_data_bus[188]), .B2(n10579), .ZN(n8888) );
  AOI22D1BWP30P140LVT U13058 ( .A1(i_data_bus[156]), .A2(n10577), .B1(
        i_data_bus[252]), .B2(n10580), .ZN(n8887) );
  ND2D1BWP30P140LVT U13059 ( .A1(n8888), .A2(n8887), .ZN(N4563) );
  AOI22D1BWP30P140LVT U13060 ( .A1(i_data_bus[186]), .A2(n10579), .B1(
        i_data_bus[218]), .B2(n10578), .ZN(n8890) );
  AOI22D1BWP30P140LVT U13061 ( .A1(i_data_bus[154]), .A2(n10577), .B1(
        i_data_bus[250]), .B2(n10580), .ZN(n8889) );
  ND2D1BWP30P140LVT U13062 ( .A1(n8890), .A2(n8889), .ZN(N4561) );
  AOI22D1BWP30P140LVT U13063 ( .A1(i_data_bus[506]), .A2(n10506), .B1(
        i_data_bus[442]), .B2(n10507), .ZN(n8892) );
  AOI22D1BWP30P140LVT U13064 ( .A1(i_data_bus[410]), .A2(n10505), .B1(
        i_data_bus[474]), .B2(n10508), .ZN(n8891) );
  ND2D1BWP30P140LVT U13065 ( .A1(n8892), .A2(n8891), .ZN(N8741) );
  AOI22D1BWP30P140LVT U13066 ( .A1(i_data_bus[398]), .A2(n10505), .B1(
        i_data_bus[494]), .B2(n10506), .ZN(n8894) );
  AOI22D1BWP30P140LVT U13067 ( .A1(i_data_bus[430]), .A2(n10507), .B1(
        i_data_bus[462]), .B2(n10508), .ZN(n8893) );
  ND2D1BWP30P140LVT U13068 ( .A1(n8894), .A2(n8893), .ZN(N8729) );
  AOI22D1BWP30P140LVT U13069 ( .A1(i_data_bus[384]), .A2(n10505), .B1(
        i_data_bus[480]), .B2(n10506), .ZN(n8896) );
  AOI22D1BWP30P140LVT U13070 ( .A1(i_data_bus[416]), .A2(n10507), .B1(
        i_data_bus[448]), .B2(n10508), .ZN(n8895) );
  ND2D1BWP30P140LVT U13071 ( .A1(n8896), .A2(n8895), .ZN(N8715) );
  AOI22D1BWP30P140LVT U13072 ( .A1(i_data_bus[420]), .A2(n10507), .B1(
        i_data_bus[484]), .B2(n10506), .ZN(n8898) );
  AOI22D1BWP30P140LVT U13073 ( .A1(i_data_bus[388]), .A2(n10505), .B1(
        i_data_bus[452]), .B2(n10508), .ZN(n8897) );
  ND2D1BWP30P140LVT U13074 ( .A1(n8898), .A2(n8897), .ZN(N8719) );
  AOI22D1BWP30P140LVT U13075 ( .A1(i_data_bus[508]), .A2(n10506), .B1(
        i_data_bus[412]), .B2(n10505), .ZN(n8900) );
  AOI22D1BWP30P140LVT U13076 ( .A1(i_data_bus[444]), .A2(n10507), .B1(
        i_data_bus[476]), .B2(n10508), .ZN(n8899) );
  ND2D1BWP30P140LVT U13077 ( .A1(n8900), .A2(n8899), .ZN(N8743) );
  AOI22D1BWP30P140LVT U13078 ( .A1(i_data_bus[431]), .A2(n10507), .B1(
        i_data_bus[495]), .B2(n10506), .ZN(n8902) );
  AOI22D1BWP30P140LVT U13079 ( .A1(i_data_bus[399]), .A2(n10505), .B1(
        i_data_bus[463]), .B2(n10508), .ZN(n8901) );
  ND2D1BWP30P140LVT U13080 ( .A1(n8902), .A2(n8901), .ZN(N8730) );
  AOI22D1BWP30P140LVT U13081 ( .A1(i_data_bus[443]), .A2(n10507), .B1(
        i_data_bus[411]), .B2(n10505), .ZN(n8904) );
  AOI22D1BWP30P140LVT U13082 ( .A1(i_data_bus[507]), .A2(n10506), .B1(
        i_data_bus[475]), .B2(n10508), .ZN(n8903) );
  ND2D1BWP30P140LVT U13083 ( .A1(n8904), .A2(n8903), .ZN(N8742) );
  AOI22D1BWP30P140LVT U13084 ( .A1(i_data_bus[433]), .A2(n10507), .B1(
        i_data_bus[497]), .B2(n10506), .ZN(n8906) );
  AOI22D1BWP30P140LVT U13085 ( .A1(i_data_bus[401]), .A2(n10505), .B1(
        i_data_bus[465]), .B2(n10508), .ZN(n8905) );
  ND2D1BWP30P140LVT U13086 ( .A1(n8906), .A2(n8905), .ZN(N8732) );
  AOI22D1BWP30P140LVT U13087 ( .A1(i_data_bus[250]), .A2(n10449), .B1(
        i_data_bus[218]), .B2(n10451), .ZN(n8908) );
  AOI22D1BWP30P140LVT U13088 ( .A1(i_data_bus[186]), .A2(n10450), .B1(
        i_data_bus[154]), .B2(n10452), .ZN(n8907) );
  ND2D1BWP30P140LVT U13089 ( .A1(n8908), .A2(n8907), .ZN(N12057) );
  AOI22D1BWP30P140LVT U13090 ( .A1(i_data_bus[214]), .A2(n10451), .B1(
        i_data_bus[246]), .B2(n10449), .ZN(n8910) );
  AOI22D1BWP30P140LVT U13091 ( .A1(i_data_bus[182]), .A2(n10450), .B1(
        i_data_bus[150]), .B2(n10452), .ZN(n8909) );
  ND2D1BWP30P140LVT U13092 ( .A1(n8910), .A2(n8909), .ZN(N12053) );
  AOI22D1BWP30P140LVT U13093 ( .A1(i_data_bus[236]), .A2(n10449), .B1(
        i_data_bus[204]), .B2(n10451), .ZN(n8912) );
  AOI22D1BWP30P140LVT U13094 ( .A1(i_data_bus[172]), .A2(n10450), .B1(
        i_data_bus[140]), .B2(n10452), .ZN(n8911) );
  ND2D1BWP30P140LVT U13095 ( .A1(n8912), .A2(n8911), .ZN(N12043) );
  AOI22D1BWP30P140LVT U13096 ( .A1(i_data_bus[185]), .A2(n10450), .B1(
        i_data_bus[217]), .B2(n10451), .ZN(n8914) );
  AOI22D1BWP30P140LVT U13097 ( .A1(i_data_bus[249]), .A2(n10449), .B1(
        i_data_bus[153]), .B2(n10452), .ZN(n8913) );
  ND2D1BWP30P140LVT U13098 ( .A1(n8914), .A2(n8913), .ZN(N12056) );
  AOI22D1BWP30P140LVT U13099 ( .A1(i_data_bus[235]), .A2(n10449), .B1(
        i_data_bus[171]), .B2(n10450), .ZN(n8916) );
  AOI22D1BWP30P140LVT U13100 ( .A1(i_data_bus[203]), .A2(n10451), .B1(
        i_data_bus[139]), .B2(n10452), .ZN(n8915) );
  ND2D1BWP30P140LVT U13101 ( .A1(n8916), .A2(n8915), .ZN(N12042) );
  AOI22D1BWP30P140LVT U13102 ( .A1(i_data_bus[198]), .A2(n10451), .B1(
        i_data_bus[166]), .B2(n10450), .ZN(n8918) );
  AOI22D1BWP30P140LVT U13103 ( .A1(i_data_bus[230]), .A2(n10449), .B1(
        i_data_bus[134]), .B2(n10452), .ZN(n8917) );
  ND2D1BWP30P140LVT U13104 ( .A1(n8918), .A2(n8917), .ZN(N12037) );
  AOI22D1BWP30P140LVT U13105 ( .A1(i_data_bus[167]), .A2(n10450), .B1(
        i_data_bus[199]), .B2(n10451), .ZN(n8920) );
  AOI22D1BWP30P140LVT U13106 ( .A1(i_data_bus[231]), .A2(n10449), .B1(
        i_data_bus[135]), .B2(n10452), .ZN(n8919) );
  ND2D1BWP30P140LVT U13107 ( .A1(n8920), .A2(n8919), .ZN(N12038) );
  AOI22D1BWP30P140LVT U13108 ( .A1(i_data_bus[227]), .A2(n10449), .B1(
        i_data_bus[195]), .B2(n10451), .ZN(n8922) );
  AOI22D1BWP30P140LVT U13109 ( .A1(i_data_bus[163]), .A2(n10450), .B1(
        i_data_bus[131]), .B2(n10452), .ZN(n8921) );
  ND2D1BWP30P140LVT U13110 ( .A1(n8922), .A2(n8921), .ZN(N12034) );
  AOI22D1BWP30P140LVT U13111 ( .A1(i_data_bus[201]), .A2(n10451), .B1(
        i_data_bus[169]), .B2(n10450), .ZN(n8924) );
  AOI22D1BWP30P140LVT U13112 ( .A1(i_data_bus[233]), .A2(n10449), .B1(
        i_data_bus[137]), .B2(n10452), .ZN(n8923) );
  ND2D1BWP30P140LVT U13113 ( .A1(n8924), .A2(n8923), .ZN(N12040) );
  AOI22D1BWP30P140LVT U13114 ( .A1(i_data_bus[190]), .A2(n10450), .B1(
        i_data_bus[254]), .B2(n10449), .ZN(n8926) );
  AOI22D1BWP30P140LVT U13115 ( .A1(i_data_bus[222]), .A2(n10451), .B1(
        i_data_bus[158]), .B2(n10452), .ZN(n8925) );
  ND2D1BWP30P140LVT U13116 ( .A1(n8926), .A2(n8925), .ZN(N12061) );
  AOI22D1BWP30P140LVT U13117 ( .A1(i_data_bus[214]), .A2(n10610), .B1(
        i_data_bus[182]), .B2(n10609), .ZN(n8928) );
  AOI22D1BWP30P140LVT U13118 ( .A1(i_data_bus[150]), .A2(n10612), .B1(
        i_data_bus[246]), .B2(n10611), .ZN(n8927) );
  ND2D1BWP30P140LVT U13119 ( .A1(n8928), .A2(n8927), .ZN(N2683) );
  AOI22D1BWP30P140LVT U13120 ( .A1(i_data_bus[160]), .A2(n10609), .B1(
        i_data_bus[192]), .B2(n10610), .ZN(n8930) );
  AOI22D1BWP30P140LVT U13121 ( .A1(i_data_bus[128]), .A2(n10612), .B1(
        i_data_bus[224]), .B2(n10611), .ZN(n8929) );
  ND2D1BWP30P140LVT U13122 ( .A1(n8930), .A2(n8929), .ZN(N2661) );
  AOI22D1BWP30P140LVT U13123 ( .A1(i_data_bus[205]), .A2(n10610), .B1(
        i_data_bus[173]), .B2(n10609), .ZN(n8932) );
  AOI22D1BWP30P140LVT U13124 ( .A1(i_data_bus[141]), .A2(n10612), .B1(
        i_data_bus[237]), .B2(n10611), .ZN(n8931) );
  ND2D1BWP30P140LVT U13125 ( .A1(n8932), .A2(n8931), .ZN(N2674) );
  AOI22D1BWP30P140LVT U13126 ( .A1(i_data_bus[207]), .A2(n10610), .B1(
        i_data_bus[143]), .B2(n10612), .ZN(n8934) );
  AOI22D1BWP30P140LVT U13127 ( .A1(i_data_bus[175]), .A2(n10609), .B1(
        i_data_bus[239]), .B2(n10611), .ZN(n8933) );
  ND2D1BWP30P140LVT U13128 ( .A1(n8934), .A2(n8933), .ZN(N2676) );
  AOI22D1BWP30P140LVT U13129 ( .A1(i_data_bus[181]), .A2(n10609), .B1(
        i_data_bus[213]), .B2(n10610), .ZN(n8936) );
  AOI22D1BWP30P140LVT U13130 ( .A1(i_data_bus[149]), .A2(n10612), .B1(
        i_data_bus[245]), .B2(n10611), .ZN(n8935) );
  ND2D1BWP30P140LVT U13131 ( .A1(n8936), .A2(n8935), .ZN(N2682) );
  AOI22D1BWP30P140LVT U13132 ( .A1(i_data_bus[159]), .A2(n10612), .B1(
        i_data_bus[191]), .B2(n10609), .ZN(n8938) );
  AOI22D1BWP30P140LVT U13133 ( .A1(i_data_bus[223]), .A2(n10610), .B1(
        i_data_bus[255]), .B2(n10611), .ZN(n8937) );
  ND2D1BWP30P140LVT U13134 ( .A1(n8938), .A2(n8937), .ZN(N2692) );
  AOI22D1BWP30P140LVT U13135 ( .A1(i_data_bus[183]), .A2(n10609), .B1(
        i_data_bus[151]), .B2(n10612), .ZN(n8940) );
  AOI22D1BWP30P140LVT U13136 ( .A1(i_data_bus[215]), .A2(n10610), .B1(
        i_data_bus[247]), .B2(n10611), .ZN(n8939) );
  ND2D1BWP30P140LVT U13137 ( .A1(n8940), .A2(n8939), .ZN(N2684) );
  AOI22D1BWP30P140LVT U13138 ( .A1(i_data_bus[848]), .A2(n10432), .B1(
        i_data_bus[880]), .B2(n10431), .ZN(n8942) );
  AOI22D1BWP30P140LVT U13139 ( .A1(i_data_bus[784]), .A2(n10429), .B1(
        i_data_bus[816]), .B2(n10430), .ZN(n8941) );
  ND2D1BWP30P140LVT U13140 ( .A1(n8942), .A2(n8941), .ZN(N13127) );
  AOI22D1BWP30P140LVT U13141 ( .A1(i_data_bus[887]), .A2(n10431), .B1(
        i_data_bus[791]), .B2(n10429), .ZN(n8944) );
  AOI22D1BWP30P140LVT U13142 ( .A1(i_data_bus[855]), .A2(n10432), .B1(
        i_data_bus[823]), .B2(n10430), .ZN(n8943) );
  ND2D1BWP30P140LVT U13143 ( .A1(n8944), .A2(n8943), .ZN(N13134) );
  AOI22D1BWP30P140LVT U13144 ( .A1(i_data_bus[789]), .A2(n10429), .B1(
        i_data_bus[853]), .B2(n10432), .ZN(n8946) );
  AOI22D1BWP30P140LVT U13145 ( .A1(i_data_bus[885]), .A2(n10431), .B1(
        i_data_bus[821]), .B2(n10430), .ZN(n8945) );
  ND2D1BWP30P140LVT U13146 ( .A1(n8946), .A2(n8945), .ZN(N13132) );
  AOI22D1BWP30P140LVT U13147 ( .A1(i_data_bus[841]), .A2(n10432), .B1(
        i_data_bus[777]), .B2(n10429), .ZN(n8948) );
  AOI22D1BWP30P140LVT U13148 ( .A1(i_data_bus[873]), .A2(n10431), .B1(
        i_data_bus[809]), .B2(n10430), .ZN(n8947) );
  ND2D1BWP30P140LVT U13149 ( .A1(n8948), .A2(n8947), .ZN(N13120) );
  AOI22D1BWP30P140LVT U13150 ( .A1(i_data_bus[836]), .A2(n10432), .B1(
        i_data_bus[868]), .B2(n10431), .ZN(n8950) );
  AOI22D1BWP30P140LVT U13151 ( .A1(i_data_bus[772]), .A2(n10429), .B1(
        i_data_bus[804]), .B2(n10430), .ZN(n8949) );
  ND2D1BWP30P140LVT U13152 ( .A1(n8950), .A2(n8949), .ZN(N13115) );
  AOI22D1BWP30P140LVT U13153 ( .A1(i_data_bus[797]), .A2(n10429), .B1(
        i_data_bus[861]), .B2(n10432), .ZN(n8952) );
  AOI22D1BWP30P140LVT U13154 ( .A1(i_data_bus[893]), .A2(n10431), .B1(
        i_data_bus[829]), .B2(n10430), .ZN(n8951) );
  ND2D1BWP30P140LVT U13155 ( .A1(n8952), .A2(n8951), .ZN(N13140) );
  AOI22D1BWP30P140LVT U13156 ( .A1(i_data_bus[895]), .A2(n10431), .B1(
        i_data_bus[799]), .B2(n10429), .ZN(n8954) );
  AOI22D1BWP30P140LVT U13157 ( .A1(i_data_bus[863]), .A2(n10432), .B1(
        i_data_bus[831]), .B2(n10430), .ZN(n8953) );
  ND2D1BWP30P140LVT U13158 ( .A1(n8954), .A2(n8953), .ZN(N13142) );
  AOI22D1BWP30P140LVT U13159 ( .A1(i_data_bus[856]), .A2(n10432), .B1(
        i_data_bus[792]), .B2(n10429), .ZN(n8956) );
  AOI22D1BWP30P140LVT U13160 ( .A1(i_data_bus[888]), .A2(n10431), .B1(
        i_data_bus[824]), .B2(n10430), .ZN(n8955) );
  ND2D1BWP30P140LVT U13161 ( .A1(n8956), .A2(n8955), .ZN(N13135) );
  AOI22D1BWP30P140LVT U13162 ( .A1(i_data_bus[881]), .A2(n10431), .B1(
        i_data_bus[849]), .B2(n10432), .ZN(n8958) );
  AOI22D1BWP30P140LVT U13163 ( .A1(i_data_bus[785]), .A2(n10429), .B1(
        i_data_bus[817]), .B2(n10430), .ZN(n8957) );
  ND2D1BWP30P140LVT U13164 ( .A1(n8958), .A2(n8957), .ZN(N13128) );
  AOI22D1BWP30P140LVT U13165 ( .A1(i_data_bus[771]), .A2(n10429), .B1(
        i_data_bus[867]), .B2(n10431), .ZN(n8960) );
  AOI22D1BWP30P140LVT U13166 ( .A1(i_data_bus[835]), .A2(n10432), .B1(
        i_data_bus[803]), .B2(n10430), .ZN(n8959) );
  ND2D1BWP30P140LVT U13167 ( .A1(n8960), .A2(n8959), .ZN(N13114) );
  AOI22D1BWP30P140LVT U13168 ( .A1(i_data_bus[882]), .A2(n10431), .B1(
        i_data_bus[786]), .B2(n10429), .ZN(n8962) );
  AOI22D1BWP30P140LVT U13169 ( .A1(i_data_bus[850]), .A2(n10432), .B1(
        i_data_bus[818]), .B2(n10430), .ZN(n8961) );
  ND2D1BWP30P140LVT U13170 ( .A1(n8962), .A2(n8961), .ZN(N13129) );
  AOI22D1BWP30P140LVT U13171 ( .A1(i_data_bus[222]), .A2(n10514), .B1(
        i_data_bus[190]), .B2(n10515), .ZN(n8964) );
  AOI22D1BWP30P140LVT U13172 ( .A1(i_data_bus[158]), .A2(n10513), .B1(
        i_data_bus[254]), .B2(n10516), .ZN(n8963) );
  ND2D1BWP30P140LVT U13173 ( .A1(n8964), .A2(n8963), .ZN(N8313) );
  AOI22D1BWP30P140LVT U13174 ( .A1(i_data_bus[214]), .A2(n10514), .B1(
        i_data_bus[150]), .B2(n10513), .ZN(n8966) );
  AOI22D1BWP30P140LVT U13175 ( .A1(i_data_bus[182]), .A2(n10515), .B1(
        i_data_bus[246]), .B2(n10516), .ZN(n8965) );
  ND2D1BWP30P140LVT U13176 ( .A1(n8966), .A2(n8965), .ZN(N8305) );
  AOI22D1BWP30P140LVT U13177 ( .A1(i_data_bus[208]), .A2(n10514), .B1(
        i_data_bus[176]), .B2(n10515), .ZN(n8968) );
  AOI22D1BWP30P140LVT U13178 ( .A1(i_data_bus[144]), .A2(n10513), .B1(
        i_data_bus[240]), .B2(n10516), .ZN(n8967) );
  ND2D1BWP30P140LVT U13179 ( .A1(n8968), .A2(n8967), .ZN(N8299) );
  AOI22D1BWP30P140LVT U13180 ( .A1(i_data_bus[179]), .A2(n10515), .B1(
        i_data_bus[147]), .B2(n10513), .ZN(n8970) );
  AOI22D1BWP30P140LVT U13181 ( .A1(i_data_bus[211]), .A2(n10514), .B1(
        i_data_bus[243]), .B2(n10516), .ZN(n8969) );
  ND2D1BWP30P140LVT U13182 ( .A1(n8970), .A2(n8969), .ZN(N8302) );
  AOI22D1BWP30P140LVT U13183 ( .A1(i_data_bus[181]), .A2(n10515), .B1(
        i_data_bus[213]), .B2(n10514), .ZN(n8972) );
  AOI22D1BWP30P140LVT U13184 ( .A1(i_data_bus[149]), .A2(n10513), .B1(
        i_data_bus[245]), .B2(n10516), .ZN(n8971) );
  ND2D1BWP30P140LVT U13185 ( .A1(n8972), .A2(n8971), .ZN(N8304) );
  AOI22D1BWP30P140LVT U13186 ( .A1(i_data_bus[168]), .A2(n10515), .B1(
        i_data_bus[136]), .B2(n10513), .ZN(n8974) );
  AOI22D1BWP30P140LVT U13187 ( .A1(i_data_bus[200]), .A2(n10514), .B1(
        i_data_bus[232]), .B2(n10516), .ZN(n8973) );
  ND2D1BWP30P140LVT U13188 ( .A1(n8974), .A2(n8973), .ZN(N8291) );
  AOI22D1BWP30P140LVT U13189 ( .A1(i_data_bus[205]), .A2(n10514), .B1(
        i_data_bus[141]), .B2(n10513), .ZN(n8976) );
  AOI22D1BWP30P140LVT U13190 ( .A1(i_data_bus[173]), .A2(n10515), .B1(
        i_data_bus[237]), .B2(n10516), .ZN(n8975) );
  ND2D1BWP30P140LVT U13191 ( .A1(n8976), .A2(n8975), .ZN(N8296) );
  AOI22D1BWP30P140LVT U13192 ( .A1(i_data_bus[178]), .A2(n10515), .B1(
        i_data_bus[146]), .B2(n10513), .ZN(n8978) );
  AOI22D1BWP30P140LVT U13193 ( .A1(i_data_bus[210]), .A2(n10514), .B1(
        i_data_bus[242]), .B2(n10516), .ZN(n8977) );
  ND2D1BWP30P140LVT U13194 ( .A1(n8978), .A2(n8977), .ZN(N8301) );
  AOI22D1BWP30P140LVT U13195 ( .A1(i_data_bus[133]), .A2(n10513), .B1(
        i_data_bus[197]), .B2(n10514), .ZN(n8980) );
  AOI22D1BWP30P140LVT U13196 ( .A1(i_data_bus[165]), .A2(n10515), .B1(
        i_data_bus[229]), .B2(n10516), .ZN(n8979) );
  ND2D1BWP30P140LVT U13197 ( .A1(n8980), .A2(n8979), .ZN(N8288) );
  AOI22D1BWP30P140LVT U13198 ( .A1(i_data_bus[154]), .A2(n10513), .B1(
        i_data_bus[218]), .B2(n10514), .ZN(n8982) );
  AOI22D1BWP30P140LVT U13199 ( .A1(i_data_bus[186]), .A2(n10515), .B1(
        i_data_bus[250]), .B2(n10516), .ZN(n8981) );
  ND2D1BWP30P140LVT U13200 ( .A1(n8982), .A2(n8981), .ZN(N8309) );
  AOI22D1BWP30P140LVT U13201 ( .A1(i_data_bus[168]), .A2(n10545), .B1(
        i_data_bus[232]), .B2(n10547), .ZN(n8984) );
  AOI22D1BWP30P140LVT U13202 ( .A1(i_data_bus[200]), .A2(n10548), .B1(
        i_data_bus[136]), .B2(n10546), .ZN(n8983) );
  ND2D1BWP30P140LVT U13203 ( .A1(n8984), .A2(n8983), .ZN(N6417) );
  AOI22D1BWP30P140LVT U13204 ( .A1(i_data_bus[255]), .A2(n10547), .B1(
        i_data_bus[191]), .B2(n10545), .ZN(n8986) );
  AOI22D1BWP30P140LVT U13205 ( .A1(i_data_bus[223]), .A2(n10548), .B1(
        i_data_bus[159]), .B2(n10546), .ZN(n8985) );
  ND2D1BWP30P140LVT U13206 ( .A1(n8986), .A2(n8985), .ZN(N6440) );
  AOI22D1BWP30P140LVT U13207 ( .A1(i_data_bus[235]), .A2(n10547), .B1(
        i_data_bus[171]), .B2(n10545), .ZN(n8988) );
  AOI22D1BWP30P140LVT U13208 ( .A1(i_data_bus[203]), .A2(n10548), .B1(
        i_data_bus[139]), .B2(n10546), .ZN(n8987) );
  ND2D1BWP30P140LVT U13209 ( .A1(n8988), .A2(n8987), .ZN(N6420) );
  AOI22D1BWP30P140LVT U13210 ( .A1(i_data_bus[185]), .A2(n10545), .B1(
        i_data_bus[217]), .B2(n10548), .ZN(n8990) );
  AOI22D1BWP30P140LVT U13211 ( .A1(i_data_bus[249]), .A2(n10547), .B1(
        i_data_bus[153]), .B2(n10546), .ZN(n8989) );
  ND2D1BWP30P140LVT U13212 ( .A1(n8990), .A2(n8989), .ZN(N6434) );
  AOI22D1BWP30P140LVT U13213 ( .A1(i_data_bus[231]), .A2(n10547), .B1(
        i_data_bus[199]), .B2(n10548), .ZN(n8992) );
  AOI22D1BWP30P140LVT U13214 ( .A1(i_data_bus[167]), .A2(n10545), .B1(
        i_data_bus[135]), .B2(n10546), .ZN(n8991) );
  ND2D1BWP30P140LVT U13215 ( .A1(n8992), .A2(n8991), .ZN(N6416) );
  AOI22D1BWP30P140LVT U13216 ( .A1(i_data_bus[173]), .A2(n10545), .B1(
        i_data_bus[237]), .B2(n10547), .ZN(n8994) );
  AOI22D1BWP30P140LVT U13217 ( .A1(i_data_bus[205]), .A2(n10548), .B1(
        i_data_bus[141]), .B2(n10546), .ZN(n8993) );
  ND2D1BWP30P140LVT U13218 ( .A1(n8994), .A2(n8993), .ZN(N6422) );
  AOI22D1BWP30P140LVT U13219 ( .A1(i_data_bus[204]), .A2(n10548), .B1(
        i_data_bus[172]), .B2(n10545), .ZN(n8996) );
  AOI22D1BWP30P140LVT U13220 ( .A1(i_data_bus[236]), .A2(n10547), .B1(
        i_data_bus[140]), .B2(n10546), .ZN(n8995) );
  ND2D1BWP30P140LVT U13221 ( .A1(n8996), .A2(n8995), .ZN(N6421) );
  AOI22D1BWP30P140LVT U13222 ( .A1(i_data_bus[174]), .A2(n10545), .B1(
        i_data_bus[238]), .B2(n10547), .ZN(n8998) );
  AOI22D1BWP30P140LVT U13223 ( .A1(i_data_bus[206]), .A2(n10548), .B1(
        i_data_bus[142]), .B2(n10546), .ZN(n8997) );
  ND2D1BWP30P140LVT U13224 ( .A1(n8998), .A2(n8997), .ZN(N6423) );
  AOI22D1BWP30P140LVT U13225 ( .A1(i_data_bus[210]), .A2(n10548), .B1(
        i_data_bus[242]), .B2(n10547), .ZN(n9000) );
  AOI22D1BWP30P140LVT U13226 ( .A1(i_data_bus[178]), .A2(n10545), .B1(
        i_data_bus[146]), .B2(n10546), .ZN(n8999) );
  ND2D1BWP30P140LVT U13227 ( .A1(n9000), .A2(n8999), .ZN(N6427) );
  AOI22D1BWP30P140LVT U13228 ( .A1(i_data_bus[258]), .A2(n10575), .B1(
        i_data_bus[290]), .B2(n10573), .ZN(n9002) );
  AOI22D1BWP30P140LVT U13229 ( .A1(i_data_bus[322]), .A2(n10576), .B1(
        i_data_bus[354]), .B2(n10574), .ZN(n9001) );
  ND2D1BWP30P140LVT U13230 ( .A1(n9002), .A2(n9001), .ZN(N4753) );
  AOI22D1BWP30P140LVT U13231 ( .A1(i_data_bus[310]), .A2(n10573), .B1(
        i_data_bus[342]), .B2(n10576), .ZN(n9004) );
  AOI22D1BWP30P140LVT U13232 ( .A1(i_data_bus[278]), .A2(n10575), .B1(
        i_data_bus[374]), .B2(n10574), .ZN(n9003) );
  ND2D1BWP30P140LVT U13233 ( .A1(n9004), .A2(n9003), .ZN(N4773) );
  AOI22D1BWP30P140LVT U13234 ( .A1(i_data_bus[303]), .A2(n10573), .B1(
        i_data_bus[335]), .B2(n10576), .ZN(n9006) );
  AOI22D1BWP30P140LVT U13235 ( .A1(i_data_bus[271]), .A2(n10575), .B1(
        i_data_bus[367]), .B2(n10574), .ZN(n9005) );
  ND2D1BWP30P140LVT U13236 ( .A1(n9006), .A2(n9005), .ZN(N4766) );
  AOI22D1BWP30P140LVT U13237 ( .A1(i_data_bus[313]), .A2(n10573), .B1(
        i_data_bus[281]), .B2(n10575), .ZN(n9008) );
  AOI22D1BWP30P140LVT U13238 ( .A1(i_data_bus[345]), .A2(n10576), .B1(
        i_data_bus[377]), .B2(n10574), .ZN(n9007) );
  ND2D1BWP30P140LVT U13239 ( .A1(n9008), .A2(n9007), .ZN(N4776) );
  AOI22D1BWP30P140LVT U13240 ( .A1(i_data_bus[311]), .A2(n10573), .B1(
        i_data_bus[343]), .B2(n10576), .ZN(n9010) );
  AOI22D1BWP30P140LVT U13241 ( .A1(i_data_bus[279]), .A2(n10575), .B1(
        i_data_bus[375]), .B2(n10574), .ZN(n9009) );
  ND2D1BWP30P140LVT U13242 ( .A1(n9010), .A2(n9009), .ZN(N4774) );
  AOI22D1BWP30P140LVT U13243 ( .A1(i_data_bus[287]), .A2(n10575), .B1(
        i_data_bus[319]), .B2(n10573), .ZN(n9012) );
  AOI22D1BWP30P140LVT U13244 ( .A1(i_data_bus[351]), .A2(n10576), .B1(
        i_data_bus[383]), .B2(n10574), .ZN(n9011) );
  ND2D1BWP30P140LVT U13245 ( .A1(n9012), .A2(n9011), .ZN(N4782) );
  AOI22D1BWP30P140LVT U13246 ( .A1(i_data_bus[341]), .A2(n10576), .B1(
        i_data_bus[277]), .B2(n10575), .ZN(n9014) );
  AOI22D1BWP30P140LVT U13247 ( .A1(i_data_bus[309]), .A2(n10573), .B1(
        i_data_bus[373]), .B2(n10574), .ZN(n9013) );
  ND2D1BWP30P140LVT U13248 ( .A1(n9014), .A2(n9013), .ZN(N4772) );
  AOI22D1BWP30P140LVT U13249 ( .A1(i_data_bus[306]), .A2(n10573), .B1(
        i_data_bus[274]), .B2(n10575), .ZN(n9016) );
  AOI22D1BWP30P140LVT U13250 ( .A1(i_data_bus[338]), .A2(n10576), .B1(
        i_data_bus[370]), .B2(n10574), .ZN(n9015) );
  ND2D1BWP30P140LVT U13251 ( .A1(n9016), .A2(n9015), .ZN(N4769) );
  AOI22D1BWP30P140LVT U13252 ( .A1(i_data_bus[329]), .A2(n10576), .B1(
        i_data_bus[297]), .B2(n10573), .ZN(n9018) );
  AOI22D1BWP30P140LVT U13253 ( .A1(i_data_bus[265]), .A2(n10575), .B1(
        i_data_bus[361]), .B2(n10574), .ZN(n9017) );
  ND2D1BWP30P140LVT U13254 ( .A1(n9018), .A2(n9017), .ZN(N4760) );
  AOI22D1BWP30P140LVT U13255 ( .A1(i_data_bus[282]), .A2(n10575), .B1(
        i_data_bus[314]), .B2(n10573), .ZN(n9020) );
  AOI22D1BWP30P140LVT U13256 ( .A1(i_data_bus[346]), .A2(n10576), .B1(
        i_data_bus[378]), .B2(n10574), .ZN(n9019) );
  ND2D1BWP30P140LVT U13257 ( .A1(n9020), .A2(n9019), .ZN(N4777) );
  AOI22D1BWP30P140LVT U13258 ( .A1(i_data_bus[196]), .A2(n10548), .B1(
        i_data_bus[164]), .B2(n10545), .ZN(n9022) );
  AOI22D1BWP30P140LVT U13259 ( .A1(i_data_bus[132]), .A2(n10546), .B1(
        i_data_bus[228]), .B2(n10547), .ZN(n9021) );
  ND2D1BWP30P140LVT U13260 ( .A1(n9022), .A2(n9021), .ZN(N6413) );
  AOI22D1BWP30P140LVT U13261 ( .A1(i_data_bus[202]), .A2(n10548), .B1(
        i_data_bus[138]), .B2(n10546), .ZN(n9024) );
  AOI22D1BWP30P140LVT U13262 ( .A1(i_data_bus[170]), .A2(n10545), .B1(
        i_data_bus[234]), .B2(n10547), .ZN(n9023) );
  ND2D1BWP30P140LVT U13263 ( .A1(n9024), .A2(n9023), .ZN(N6419) );
  AOI22D1BWP30P140LVT U13264 ( .A1(i_data_bus[137]), .A2(n10546), .B1(
        i_data_bus[169]), .B2(n10545), .ZN(n9026) );
  AOI22D1BWP30P140LVT U13265 ( .A1(i_data_bus[201]), .A2(n10548), .B1(
        i_data_bus[233]), .B2(n10547), .ZN(n9025) );
  ND2D1BWP30P140LVT U13266 ( .A1(n9026), .A2(n9025), .ZN(N6418) );
  AOI22D1BWP30P140LVT U13267 ( .A1(i_data_bus[194]), .A2(n10548), .B1(
        i_data_bus[162]), .B2(n10545), .ZN(n9028) );
  AOI22D1BWP30P140LVT U13268 ( .A1(i_data_bus[130]), .A2(n10546), .B1(
        i_data_bus[226]), .B2(n10547), .ZN(n9027) );
  ND2D1BWP30P140LVT U13269 ( .A1(n9028), .A2(n9027), .ZN(N6411) );
  AOI22D1BWP30P140LVT U13270 ( .A1(i_data_bus[175]), .A2(n10545), .B1(
        i_data_bus[143]), .B2(n10546), .ZN(n9030) );
  AOI22D1BWP30P140LVT U13271 ( .A1(i_data_bus[207]), .A2(n10548), .B1(
        i_data_bus[239]), .B2(n10547), .ZN(n9029) );
  ND2D1BWP30P140LVT U13272 ( .A1(n9030), .A2(n9029), .ZN(N6424) );
  AOI22D1BWP30P140LVT U13273 ( .A1(i_data_bus[220]), .A2(n10548), .B1(
        i_data_bus[188]), .B2(n10545), .ZN(n9032) );
  AOI22D1BWP30P140LVT U13274 ( .A1(i_data_bus[156]), .A2(n10546), .B1(
        i_data_bus[252]), .B2(n10547), .ZN(n9031) );
  ND2D1BWP30P140LVT U13275 ( .A1(n9032), .A2(n9031), .ZN(N6437) );
  AOI22D1BWP30P140LVT U13276 ( .A1(i_data_bus[144]), .A2(n10546), .B1(
        i_data_bus[176]), .B2(n10545), .ZN(n9034) );
  AOI22D1BWP30P140LVT U13277 ( .A1(i_data_bus[208]), .A2(n10548), .B1(
        i_data_bus[240]), .B2(n10547), .ZN(n9033) );
  ND2D1BWP30P140LVT U13278 ( .A1(n9034), .A2(n9033), .ZN(N6425) );
  AOI22D1BWP30P140LVT U13279 ( .A1(i_data_bus[186]), .A2(n10545), .B1(
        i_data_bus[218]), .B2(n10548), .ZN(n9036) );
  AOI22D1BWP30P140LVT U13280 ( .A1(i_data_bus[154]), .A2(n10546), .B1(
        i_data_bus[250]), .B2(n10547), .ZN(n9035) );
  ND2D1BWP30P140LVT U13281 ( .A1(n9036), .A2(n9035), .ZN(N6435) );
  AOI22D1BWP30P140LVT U13282 ( .A1(i_data_bus[190]), .A2(n10545), .B1(
        i_data_bus[158]), .B2(n10546), .ZN(n9038) );
  AOI22D1BWP30P140LVT U13283 ( .A1(i_data_bus[222]), .A2(n10548), .B1(
        i_data_bus[254]), .B2(n10547), .ZN(n9037) );
  ND2D1BWP30P140LVT U13284 ( .A1(n9038), .A2(n9037), .ZN(N6439) );
  AOI22D1BWP30P140LVT U13285 ( .A1(i_data_bus[177]), .A2(n10545), .B1(
        i_data_bus[145]), .B2(n10546), .ZN(n9040) );
  AOI22D1BWP30P140LVT U13286 ( .A1(i_data_bus[209]), .A2(n10548), .B1(
        i_data_bus[241]), .B2(n10547), .ZN(n9039) );
  ND2D1BWP30P140LVT U13287 ( .A1(n9040), .A2(n9039), .ZN(N6426) );
  AOI22D1BWP30P140LVT U13288 ( .A1(i_data_bus[214]), .A2(n10548), .B1(
        i_data_bus[182]), .B2(n10545), .ZN(n9042) );
  AOI22D1BWP30P140LVT U13289 ( .A1(i_data_bus[150]), .A2(n10546), .B1(
        i_data_bus[246]), .B2(n10547), .ZN(n9041) );
  ND2D1BWP30P140LVT U13290 ( .A1(n9042), .A2(n9041), .ZN(N6431) );
  AOI22D1BWP30P140LVT U13291 ( .A1(i_data_bus[151]), .A2(n10546), .B1(
        i_data_bus[215]), .B2(n10548), .ZN(n9044) );
  AOI22D1BWP30P140LVT U13292 ( .A1(i_data_bus[183]), .A2(n10545), .B1(
        i_data_bus[247]), .B2(n10547), .ZN(n9043) );
  ND2D1BWP30P140LVT U13293 ( .A1(n9044), .A2(n9043), .ZN(N6432) );
  AOI22D1BWP30P140LVT U13294 ( .A1(i_data_bus[181]), .A2(n10545), .B1(
        i_data_bus[213]), .B2(n10548), .ZN(n9046) );
  AOI22D1BWP30P140LVT U13295 ( .A1(i_data_bus[149]), .A2(n10546), .B1(
        i_data_bus[245]), .B2(n10547), .ZN(n9045) );
  ND2D1BWP30P140LVT U13296 ( .A1(n9046), .A2(n9045), .ZN(N6430) );
  AOI22D1BWP30P140LVT U13297 ( .A1(i_data_bus[287]), .A2(n10447), .B1(
        i_data_bus[319]), .B2(n10448), .ZN(n9048) );
  AOI22D1BWP30P140LVT U13298 ( .A1(i_data_bus[351]), .A2(n10446), .B1(
        i_data_bus[383]), .B2(n10445), .ZN(n9047) );
  ND2D1BWP30P140LVT U13299 ( .A1(n9048), .A2(n9047), .ZN(N12278) );
  AOI22D1BWP30P140LVT U13300 ( .A1(i_data_bus[258]), .A2(n10447), .B1(
        i_data_bus[290]), .B2(n10448), .ZN(n9050) );
  AOI22D1BWP30P140LVT U13301 ( .A1(i_data_bus[322]), .A2(n10446), .B1(
        i_data_bus[354]), .B2(n10445), .ZN(n9049) );
  ND2D1BWP30P140LVT U13302 ( .A1(n9050), .A2(n9049), .ZN(N12249) );
  AOI22D1BWP30P140LVT U13303 ( .A1(i_data_bus[309]), .A2(n10448), .B1(
        i_data_bus[277]), .B2(n10447), .ZN(n9052) );
  AOI22D1BWP30P140LVT U13304 ( .A1(i_data_bus[341]), .A2(n10446), .B1(
        i_data_bus[373]), .B2(n10445), .ZN(n9051) );
  ND2D1BWP30P140LVT U13305 ( .A1(n9052), .A2(n9051), .ZN(N12268) );
  AOI22D1BWP30P140LVT U13306 ( .A1(i_data_bus[321]), .A2(n10446), .B1(
        i_data_bus[289]), .B2(n10448), .ZN(n9054) );
  AOI22D1BWP30P140LVT U13307 ( .A1(i_data_bus[257]), .A2(n10447), .B1(
        i_data_bus[353]), .B2(n10445), .ZN(n9053) );
  ND2D1BWP30P140LVT U13308 ( .A1(n9054), .A2(n9053), .ZN(N12248) );
  AOI22D1BWP30P140LVT U13309 ( .A1(i_data_bus[312]), .A2(n10448), .B1(
        i_data_bus[344]), .B2(n10446), .ZN(n9056) );
  AOI22D1BWP30P140LVT U13310 ( .A1(i_data_bus[280]), .A2(n10447), .B1(
        i_data_bus[376]), .B2(n10445), .ZN(n9055) );
  ND2D1BWP30P140LVT U13311 ( .A1(n9056), .A2(n9055), .ZN(N12271) );
  AOI22D1BWP30P140LVT U13312 ( .A1(i_data_bus[292]), .A2(n10448), .B1(
        i_data_bus[260]), .B2(n10447), .ZN(n9058) );
  AOI22D1BWP30P140LVT U13313 ( .A1(i_data_bus[324]), .A2(n10446), .B1(
        i_data_bus[356]), .B2(n10445), .ZN(n9057) );
  ND2D1BWP30P140LVT U13314 ( .A1(n9058), .A2(n9057), .ZN(N12251) );
  AOI22D1BWP30P140LVT U13315 ( .A1(i_data_bus[273]), .A2(n10447), .B1(
        i_data_bus[337]), .B2(n10446), .ZN(n9060) );
  AOI22D1BWP30P140LVT U13316 ( .A1(i_data_bus[305]), .A2(n10448), .B1(
        i_data_bus[369]), .B2(n10445), .ZN(n9059) );
  ND2D1BWP30P140LVT U13317 ( .A1(n9060), .A2(n9059), .ZN(N12264) );
  AOI22D1BWP30P140LVT U13318 ( .A1(i_data_bus[329]), .A2(n10446), .B1(
        i_data_bus[297]), .B2(n10448), .ZN(n9062) );
  AOI22D1BWP30P140LVT U13319 ( .A1(i_data_bus[265]), .A2(n10447), .B1(
        i_data_bus[361]), .B2(n10445), .ZN(n9061) );
  ND2D1BWP30P140LVT U13320 ( .A1(n9062), .A2(n9061), .ZN(N12256) );
  AOI22D1BWP30P140LVT U13321 ( .A1(i_data_bus[95]), .A2(n10613), .B1(
        i_data_bus[63]), .B2(n10614), .ZN(n9064) );
  AOI22D1BWP30P140LVT U13322 ( .A1(i_data_bus[127]), .A2(n10616), .B1(
        i_data_bus[31]), .B2(n10615), .ZN(n9063) );
  ND2D1BWP30P140LVT U13323 ( .A1(n9064), .A2(n9063), .ZN(N2476) );
  AOI22D1BWP30P140LVT U13324 ( .A1(i_data_bus[75]), .A2(n10613), .B1(
        i_data_bus[43]), .B2(n10614), .ZN(n9066) );
  AOI22D1BWP30P140LVT U13325 ( .A1(i_data_bus[107]), .A2(n10616), .B1(
        i_data_bus[11]), .B2(n10615), .ZN(n9065) );
  ND2D1BWP30P140LVT U13326 ( .A1(n9066), .A2(n9065), .ZN(N2456) );
  AOI22D1BWP30P140LVT U13327 ( .A1(i_data_bus[39]), .A2(n10614), .B1(
        i_data_bus[71]), .B2(n10613), .ZN(n9068) );
  AOI22D1BWP30P140LVT U13328 ( .A1(i_data_bus[103]), .A2(n10616), .B1(
        i_data_bus[7]), .B2(n10615), .ZN(n9067) );
  ND2D1BWP30P140LVT U13329 ( .A1(n9068), .A2(n9067), .ZN(N2452) );
  AOI22D1BWP30P140LVT U13330 ( .A1(i_data_bus[104]), .A2(n10616), .B1(
        i_data_bus[72]), .B2(n10613), .ZN(n9070) );
  AOI22D1BWP30P140LVT U13331 ( .A1(i_data_bus[40]), .A2(n10614), .B1(
        i_data_bus[8]), .B2(n10615), .ZN(n9069) );
  ND2D1BWP30P140LVT U13332 ( .A1(n9070), .A2(n9069), .ZN(N2453) );
  AOI22D1BWP30P140LVT U13333 ( .A1(i_data_bus[83]), .A2(n10613), .B1(
        i_data_bus[115]), .B2(n10616), .ZN(n9072) );
  AOI22D1BWP30P140LVT U13334 ( .A1(i_data_bus[51]), .A2(n10614), .B1(
        i_data_bus[19]), .B2(n10615), .ZN(n9071) );
  ND2D1BWP30P140LVT U13335 ( .A1(n9072), .A2(n9071), .ZN(N2464) );
  AOI22D1BWP30P140LVT U13336 ( .A1(i_data_bus[52]), .A2(n10614), .B1(
        i_data_bus[116]), .B2(n10616), .ZN(n9074) );
  AOI22D1BWP30P140LVT U13337 ( .A1(i_data_bus[84]), .A2(n10613), .B1(
        i_data_bus[20]), .B2(n10615), .ZN(n9073) );
  ND2D1BWP30P140LVT U13338 ( .A1(n9074), .A2(n9073), .ZN(N2465) );
  AOI22D1BWP30P140LVT U13339 ( .A1(i_data_bus[32]), .A2(n10614), .B1(
        i_data_bus[64]), .B2(n10613), .ZN(n9076) );
  AOI22D1BWP30P140LVT U13340 ( .A1(i_data_bus[96]), .A2(n10616), .B1(
        i_data_bus[0]), .B2(n10615), .ZN(n9075) );
  ND2D1BWP30P140LVT U13341 ( .A1(n9076), .A2(n9075), .ZN(N2445) );
  AOI22D1BWP30P140LVT U13342 ( .A1(i_data_bus[89]), .A2(n10613), .B1(
        i_data_bus[57]), .B2(n10614), .ZN(n9078) );
  AOI22D1BWP30P140LVT U13343 ( .A1(i_data_bus[121]), .A2(n10616), .B1(
        i_data_bus[25]), .B2(n10615), .ZN(n9077) );
  ND2D1BWP30P140LVT U13344 ( .A1(n9078), .A2(n9077), .ZN(N2470) );
  AOI22D1BWP30P140LVT U13345 ( .A1(i_data_bus[122]), .A2(n10616), .B1(
        i_data_bus[58]), .B2(n10614), .ZN(n9080) );
  AOI22D1BWP30P140LVT U13346 ( .A1(i_data_bus[90]), .A2(n10613), .B1(
        i_data_bus[26]), .B2(n10615), .ZN(n9079) );
  ND2D1BWP30P140LVT U13347 ( .A1(n9080), .A2(n9079), .ZN(N2471) );
  AOI22D1BWP30P140LVT U13348 ( .A1(i_data_bus[59]), .A2(n10614), .B1(
        i_data_bus[91]), .B2(n10613), .ZN(n9082) );
  AOI22D1BWP30P140LVT U13349 ( .A1(i_data_bus[123]), .A2(n10616), .B1(
        i_data_bus[27]), .B2(n10615), .ZN(n9081) );
  ND2D1BWP30P140LVT U13350 ( .A1(n9082), .A2(n9081), .ZN(N2472) );
  AOI22D1BWP30P140LVT U13351 ( .A1(i_data_bus[76]), .A2(n10613), .B1(
        i_data_bus[108]), .B2(n10616), .ZN(n9084) );
  AOI22D1BWP30P140LVT U13352 ( .A1(i_data_bus[44]), .A2(n10614), .B1(
        i_data_bus[12]), .B2(n10615), .ZN(n9083) );
  ND2D1BWP30P140LVT U13353 ( .A1(n9084), .A2(n9083), .ZN(N2457) );
  AOI22D1BWP30P140LVT U13354 ( .A1(i_data_bus[77]), .A2(n10613), .B1(
        i_data_bus[45]), .B2(n10614), .ZN(n9086) );
  AOI22D1BWP30P140LVT U13355 ( .A1(i_data_bus[109]), .A2(n10616), .B1(
        i_data_bus[13]), .B2(n10615), .ZN(n9085) );
  ND2D1BWP30P140LVT U13356 ( .A1(n9086), .A2(n9085), .ZN(N2458) );
  AOI22D1BWP30P140LVT U13357 ( .A1(i_data_bus[451]), .A2(n10476), .B1(
        i_data_bus[387]), .B2(n10473), .ZN(n9088) );
  AOI22D1BWP30P140LVT U13358 ( .A1(i_data_bus[483]), .A2(n10475), .B1(
        i_data_bus[419]), .B2(n10474), .ZN(n9087) );
  ND2D1BWP30P140LVT U13359 ( .A1(n9088), .A2(n9087), .ZN(N10592) );
  AOI22D1BWP30P140LVT U13360 ( .A1(i_data_bus[388]), .A2(n10473), .B1(
        i_data_bus[484]), .B2(n10475), .ZN(n9090) );
  AOI22D1BWP30P140LVT U13361 ( .A1(i_data_bus[452]), .A2(n10476), .B1(
        i_data_bus[420]), .B2(n10474), .ZN(n9089) );
  ND2D1BWP30P140LVT U13362 ( .A1(n9090), .A2(n9089), .ZN(N10593) );
  AOI22D1BWP30P140LVT U13363 ( .A1(i_data_bus[389]), .A2(n10473), .B1(
        i_data_bus[453]), .B2(n10476), .ZN(n9092) );
  AOI22D1BWP30P140LVT U13364 ( .A1(i_data_bus[485]), .A2(n10475), .B1(
        i_data_bus[421]), .B2(n10474), .ZN(n9091) );
  ND2D1BWP30P140LVT U13365 ( .A1(n9092), .A2(n9091), .ZN(N10594) );
  AOI22D1BWP30P140LVT U13366 ( .A1(i_data_bus[455]), .A2(n10476), .B1(
        i_data_bus[391]), .B2(n10473), .ZN(n9094) );
  AOI22D1BWP30P140LVT U13367 ( .A1(i_data_bus[487]), .A2(n10475), .B1(
        i_data_bus[423]), .B2(n10474), .ZN(n9093) );
  ND2D1BWP30P140LVT U13368 ( .A1(n9094), .A2(n9093), .ZN(N10596) );
  AOI22D1BWP30P140LVT U13369 ( .A1(i_data_bus[489]), .A2(n10475), .B1(
        i_data_bus[393]), .B2(n10473), .ZN(n9096) );
  AOI22D1BWP30P140LVT U13370 ( .A1(i_data_bus[457]), .A2(n10476), .B1(
        i_data_bus[425]), .B2(n10474), .ZN(n9095) );
  ND2D1BWP30P140LVT U13371 ( .A1(n9096), .A2(n9095), .ZN(N10598) );
  AOI22D1BWP30P140LVT U13372 ( .A1(i_data_bus[415]), .A2(n10473), .B1(
        i_data_bus[511]), .B2(n10475), .ZN(n9098) );
  AOI22D1BWP30P140LVT U13373 ( .A1(i_data_bus[479]), .A2(n10476), .B1(
        i_data_bus[447]), .B2(n10474), .ZN(n9097) );
  ND2D1BWP30P140LVT U13374 ( .A1(n9098), .A2(n9097), .ZN(N10620) );
  AOI22D1BWP30P140LVT U13375 ( .A1(i_data_bus[458]), .A2(n10476), .B1(
        i_data_bus[394]), .B2(n10473), .ZN(n9100) );
  AOI22D1BWP30P140LVT U13376 ( .A1(i_data_bus[490]), .A2(n10475), .B1(
        i_data_bus[426]), .B2(n10474), .ZN(n9099) );
  ND2D1BWP30P140LVT U13377 ( .A1(n9100), .A2(n9099), .ZN(N10599) );
  AOI22D1BWP30P140LVT U13378 ( .A1(i_data_bus[509]), .A2(n10475), .B1(
        i_data_bus[477]), .B2(n10476), .ZN(n9102) );
  AOI22D1BWP30P140LVT U13379 ( .A1(i_data_bus[413]), .A2(n10473), .B1(
        i_data_bus[445]), .B2(n10474), .ZN(n9101) );
  ND2D1BWP30P140LVT U13380 ( .A1(n9102), .A2(n9101), .ZN(N10618) );
  AOI22D1BWP30P140LVT U13381 ( .A1(i_data_bus[410]), .A2(n10473), .B1(
        i_data_bus[474]), .B2(n10476), .ZN(n9104) );
  AOI22D1BWP30P140LVT U13382 ( .A1(i_data_bus[506]), .A2(n10475), .B1(
        i_data_bus[442]), .B2(n10474), .ZN(n9103) );
  ND2D1BWP30P140LVT U13383 ( .A1(n9104), .A2(n9103), .ZN(N10615) );
  AOI22D1BWP30P140LVT U13384 ( .A1(i_data_bus[492]), .A2(n10475), .B1(
        i_data_bus[396]), .B2(n10473), .ZN(n9106) );
  AOI22D1BWP30P140LVT U13385 ( .A1(i_data_bus[460]), .A2(n10476), .B1(
        i_data_bus[428]), .B2(n10474), .ZN(n9105) );
  ND2D1BWP30P140LVT U13386 ( .A1(n9106), .A2(n9105), .ZN(N10601) );
  AOI22D1BWP30P140LVT U13387 ( .A1(i_data_bus[467]), .A2(n10476), .B1(
        i_data_bus[403]), .B2(n10473), .ZN(n9108) );
  AOI22D1BWP30P140LVT U13388 ( .A1(i_data_bus[499]), .A2(n10475), .B1(
        i_data_bus[435]), .B2(n10474), .ZN(n9107) );
  ND2D1BWP30P140LVT U13389 ( .A1(n9108), .A2(n9107), .ZN(N10608) );
  AOI22D1BWP30P140LVT U13390 ( .A1(i_data_bus[468]), .A2(n10476), .B1(
        i_data_bus[500]), .B2(n10475), .ZN(n9110) );
  AOI22D1BWP30P140LVT U13391 ( .A1(i_data_bus[404]), .A2(n10473), .B1(
        i_data_bus[436]), .B2(n10474), .ZN(n9109) );
  ND2D1BWP30P140LVT U13392 ( .A1(n9110), .A2(n9109), .ZN(N10609) );
  AOI22D1BWP30P140LVT U13393 ( .A1(i_data_bus[856]), .A2(n10527), .B1(
        i_data_bus[888]), .B2(n10526), .ZN(n9112) );
  AOI22D1BWP30P140LVT U13394 ( .A1(i_data_bus[792]), .A2(n10528), .B1(
        i_data_bus[824]), .B2(n10525), .ZN(n9111) );
  ND2D1BWP30P140LVT U13395 ( .A1(n9112), .A2(n9111), .ZN(N7513) );
  AOI22D1BWP30P140LVT U13396 ( .A1(i_data_bus[843]), .A2(n10527), .B1(
        i_data_bus[875]), .B2(n10526), .ZN(n9114) );
  AOI22D1BWP30P140LVT U13397 ( .A1(i_data_bus[779]), .A2(n10528), .B1(
        i_data_bus[811]), .B2(n10525), .ZN(n9113) );
  ND2D1BWP30P140LVT U13398 ( .A1(n9114), .A2(n9113), .ZN(N7500) );
  AOI22D1BWP30P140LVT U13399 ( .A1(i_data_bus[858]), .A2(n10527), .B1(
        i_data_bus[794]), .B2(n10528), .ZN(n9116) );
  AOI22D1BWP30P140LVT U13400 ( .A1(i_data_bus[890]), .A2(n10526), .B1(
        i_data_bus[826]), .B2(n10525), .ZN(n9115) );
  ND2D1BWP30P140LVT U13401 ( .A1(n9116), .A2(n9115), .ZN(N7515) );
  AOI22D1BWP30P140LVT U13402 ( .A1(i_data_bus[887]), .A2(n10526), .B1(
        i_data_bus[791]), .B2(n10528), .ZN(n9118) );
  AOI22D1BWP30P140LVT U13403 ( .A1(i_data_bus[855]), .A2(n10527), .B1(
        i_data_bus[823]), .B2(n10525), .ZN(n9117) );
  ND2D1BWP30P140LVT U13404 ( .A1(n9118), .A2(n9117), .ZN(N7512) );
  AOI22D1BWP30P140LVT U13405 ( .A1(i_data_bus[787]), .A2(n10528), .B1(
        i_data_bus[851]), .B2(n10527), .ZN(n9120) );
  AOI22D1BWP30P140LVT U13406 ( .A1(i_data_bus[883]), .A2(n10526), .B1(
        i_data_bus[819]), .B2(n10525), .ZN(n9119) );
  ND2D1BWP30P140LVT U13407 ( .A1(n9120), .A2(n9119), .ZN(N7508) );
  AOI22D1BWP30P140LVT U13408 ( .A1(i_data_bus[778]), .A2(n10528), .B1(
        i_data_bus[874]), .B2(n10526), .ZN(n9122) );
  AOI22D1BWP30P140LVT U13409 ( .A1(i_data_bus[842]), .A2(n10527), .B1(
        i_data_bus[810]), .B2(n10525), .ZN(n9121) );
  ND2D1BWP30P140LVT U13410 ( .A1(n9122), .A2(n9121), .ZN(N7499) );
  AOI22D1BWP30P140LVT U13411 ( .A1(i_data_bus[844]), .A2(n10527), .B1(
        i_data_bus[876]), .B2(n10526), .ZN(n9124) );
  AOI22D1BWP30P140LVT U13412 ( .A1(i_data_bus[780]), .A2(n10528), .B1(
        i_data_bus[812]), .B2(n10525), .ZN(n9123) );
  ND2D1BWP30P140LVT U13413 ( .A1(n9124), .A2(n9123), .ZN(N7501) );
  AOI22D1BWP30P140LVT U13414 ( .A1(i_data_bus[863]), .A2(n10527), .B1(
        i_data_bus[895]), .B2(n10526), .ZN(n9126) );
  AOI22D1BWP30P140LVT U13415 ( .A1(i_data_bus[799]), .A2(n10528), .B1(
        i_data_bus[831]), .B2(n10525), .ZN(n9125) );
  ND2D1BWP30P140LVT U13416 ( .A1(n9126), .A2(n9125), .ZN(N7520) );
  AOI22D1BWP30P140LVT U13417 ( .A1(i_data_bus[797]), .A2(n10528), .B1(
        i_data_bus[861]), .B2(n10527), .ZN(n9128) );
  AOI22D1BWP30P140LVT U13418 ( .A1(i_data_bus[893]), .A2(n10526), .B1(
        i_data_bus[829]), .B2(n10525), .ZN(n9127) );
  ND2D1BWP30P140LVT U13419 ( .A1(n9128), .A2(n9127), .ZN(N7518) );
  AOI22D1BWP30P140LVT U13420 ( .A1(i_data_bus[771]), .A2(n10528), .B1(
        i_data_bus[867]), .B2(n10526), .ZN(n9130) );
  AOI22D1BWP30P140LVT U13421 ( .A1(i_data_bus[835]), .A2(n10527), .B1(
        i_data_bus[803]), .B2(n10525), .ZN(n9129) );
  ND2D1BWP30P140LVT U13422 ( .A1(n9130), .A2(n9129), .ZN(N7492) );
  AOI22D1BWP30P140LVT U13423 ( .A1(i_data_bus[775]), .A2(n10528), .B1(
        i_data_bus[839]), .B2(n10527), .ZN(n9132) );
  AOI22D1BWP30P140LVT U13424 ( .A1(i_data_bus[871]), .A2(n10526), .B1(
        i_data_bus[807]), .B2(n10525), .ZN(n9131) );
  ND2D1BWP30P140LVT U13425 ( .A1(n9132), .A2(n9131), .ZN(N7496) );
  AOI22D1BWP30P140LVT U13426 ( .A1(i_data_bus[271]), .A2(n10605), .B1(
        i_data_bus[335]), .B2(n10607), .ZN(n9134) );
  AOI22D1BWP30P140LVT U13427 ( .A1(i_data_bus[303]), .A2(n10606), .B1(
        i_data_bus[367]), .B2(n10608), .ZN(n9133) );
  ND2D1BWP30P140LVT U13428 ( .A1(n9134), .A2(n9133), .ZN(N2892) );
  AOI22D1BWP30P140LVT U13429 ( .A1(i_data_bus[307]), .A2(n10606), .B1(
        i_data_bus[339]), .B2(n10607), .ZN(n9136) );
  AOI22D1BWP30P140LVT U13430 ( .A1(i_data_bus[275]), .A2(n10605), .B1(
        i_data_bus[371]), .B2(n10608), .ZN(n9135) );
  ND2D1BWP30P140LVT U13431 ( .A1(n9136), .A2(n9135), .ZN(N2896) );
  AOI22D1BWP30P140LVT U13432 ( .A1(i_data_bus[282]), .A2(n10605), .B1(
        i_data_bus[346]), .B2(n10607), .ZN(n9138) );
  AOI22D1BWP30P140LVT U13433 ( .A1(i_data_bus[314]), .A2(n10606), .B1(
        i_data_bus[378]), .B2(n10608), .ZN(n9137) );
  ND2D1BWP30P140LVT U13434 ( .A1(n9138), .A2(n9137), .ZN(N2903) );
  AOI22D1BWP30P140LVT U13435 ( .A1(i_data_bus[327]), .A2(n10607), .B1(
        i_data_bus[263]), .B2(n10605), .ZN(n9140) );
  AOI22D1BWP30P140LVT U13436 ( .A1(i_data_bus[295]), .A2(n10606), .B1(
        i_data_bus[359]), .B2(n10608), .ZN(n9139) );
  ND2D1BWP30P140LVT U13437 ( .A1(n9140), .A2(n9139), .ZN(N2884) );
  AOI22D1BWP30P140LVT U13438 ( .A1(i_data_bus[258]), .A2(n10605), .B1(
        i_data_bus[322]), .B2(n10607), .ZN(n9142) );
  AOI22D1BWP30P140LVT U13439 ( .A1(i_data_bus[290]), .A2(n10606), .B1(
        i_data_bus[354]), .B2(n10608), .ZN(n9141) );
  ND2D1BWP30P140LVT U13440 ( .A1(n9142), .A2(n9141), .ZN(N2879) );
  AOI22D1BWP30P140LVT U13441 ( .A1(i_data_bus[292]), .A2(n10606), .B1(
        i_data_bus[260]), .B2(n10605), .ZN(n9144) );
  AOI22D1BWP30P140LVT U13442 ( .A1(i_data_bus[324]), .A2(n10607), .B1(
        i_data_bus[356]), .B2(n10608), .ZN(n9143) );
  ND2D1BWP30P140LVT U13443 ( .A1(n9144), .A2(n9143), .ZN(N2881) );
  AOI22D1BWP30P140LVT U13444 ( .A1(i_data_bus[265]), .A2(n10605), .B1(
        i_data_bus[297]), .B2(n10606), .ZN(n9146) );
  AOI22D1BWP30P140LVT U13445 ( .A1(i_data_bus[329]), .A2(n10607), .B1(
        i_data_bus[361]), .B2(n10608), .ZN(n9145) );
  ND2D1BWP30P140LVT U13446 ( .A1(n9146), .A2(n9145), .ZN(N2886) );
  AOI22D1BWP30P140LVT U13447 ( .A1(i_data_bus[161]), .A2(n10483), .B1(
        i_data_bus[193]), .B2(n10482), .ZN(n9148) );
  AOI22D1BWP30P140LVT U13448 ( .A1(i_data_bus[129]), .A2(n10481), .B1(
        i_data_bus[225]), .B2(n10484), .ZN(n9147) );
  ND2D1BWP30P140LVT U13449 ( .A1(n9148), .A2(n9147), .ZN(N10158) );
  AOI22D1BWP30P140LVT U13450 ( .A1(i_data_bus[148]), .A2(n10481), .B1(
        i_data_bus[212]), .B2(n10482), .ZN(n9150) );
  AOI22D1BWP30P140LVT U13451 ( .A1(i_data_bus[180]), .A2(n10483), .B1(
        i_data_bus[244]), .B2(n10484), .ZN(n9149) );
  ND2D1BWP30P140LVT U13452 ( .A1(n9150), .A2(n9149), .ZN(N10177) );
  AOI22D1BWP30P140LVT U13453 ( .A1(i_data_bus[182]), .A2(n10483), .B1(
        i_data_bus[150]), .B2(n10481), .ZN(n9152) );
  AOI22D1BWP30P140LVT U13454 ( .A1(i_data_bus[214]), .A2(n10482), .B1(
        i_data_bus[246]), .B2(n10484), .ZN(n9151) );
  ND2D1BWP30P140LVT U13455 ( .A1(n9152), .A2(n9151), .ZN(N10179) );
  AOI22D1BWP30P140LVT U13456 ( .A1(i_data_bus[175]), .A2(n10483), .B1(
        i_data_bus[143]), .B2(n10481), .ZN(n9154) );
  AOI22D1BWP30P140LVT U13457 ( .A1(i_data_bus[207]), .A2(n10482), .B1(
        i_data_bus[239]), .B2(n10484), .ZN(n9153) );
  ND2D1BWP30P140LVT U13458 ( .A1(n9154), .A2(n9153), .ZN(N10172) );
  AOI22D1BWP30P140LVT U13459 ( .A1(i_data_bus[208]), .A2(n10482), .B1(
        i_data_bus[176]), .B2(n10483), .ZN(n9156) );
  AOI22D1BWP30P140LVT U13460 ( .A1(i_data_bus[144]), .A2(n10481), .B1(
        i_data_bus[240]), .B2(n10484), .ZN(n9155) );
  ND2D1BWP30P140LVT U13461 ( .A1(n9156), .A2(n9155), .ZN(N10173) );
  AOI22D1BWP30P140LVT U13462 ( .A1(i_data_bus[159]), .A2(n10481), .B1(
        i_data_bus[191]), .B2(n10483), .ZN(n9158) );
  AOI22D1BWP30P140LVT U13463 ( .A1(i_data_bus[223]), .A2(n10482), .B1(
        i_data_bus[255]), .B2(n10484), .ZN(n9157) );
  ND2D1BWP30P140LVT U13464 ( .A1(n9158), .A2(n9157), .ZN(N10188) );
  AOI22D1BWP30P140LVT U13465 ( .A1(i_data_bus[177]), .A2(n10483), .B1(
        i_data_bus[145]), .B2(n10481), .ZN(n9160) );
  AOI22D1BWP30P140LVT U13466 ( .A1(i_data_bus[209]), .A2(n10482), .B1(
        i_data_bus[241]), .B2(n10484), .ZN(n9159) );
  ND2D1BWP30P140LVT U13467 ( .A1(n9160), .A2(n9159), .ZN(N10174) );
  AOI22D1BWP30P140LVT U13468 ( .A1(i_data_bus[38]), .A2(n10550), .B1(
        i_data_bus[102]), .B2(n10549), .ZN(n9162) );
  AOI22D1BWP30P140LVT U13469 ( .A1(i_data_bus[6]), .A2(n10552), .B1(
        i_data_bus[70]), .B2(n10551), .ZN(n9161) );
  ND2D1BWP30P140LVT U13470 ( .A1(n9162), .A2(n9161), .ZN(N6199) );
  AOI22D1BWP30P140LVT U13471 ( .A1(i_data_bus[45]), .A2(n10550), .B1(
        i_data_bus[13]), .B2(n10552), .ZN(n9164) );
  AOI22D1BWP30P140LVT U13472 ( .A1(i_data_bus[109]), .A2(n10549), .B1(
        i_data_bus[77]), .B2(n10551), .ZN(n9163) );
  ND2D1BWP30P140LVT U13473 ( .A1(n9164), .A2(n9163), .ZN(N6206) );
  AOI22D1BWP30P140LVT U13474 ( .A1(i_data_bus[32]), .A2(n10550), .B1(
        i_data_bus[96]), .B2(n10549), .ZN(n9166) );
  AOI22D1BWP30P140LVT U13475 ( .A1(i_data_bus[0]), .A2(n10552), .B1(
        i_data_bus[64]), .B2(n10551), .ZN(n9165) );
  ND2D1BWP30P140LVT U13476 ( .A1(n9166), .A2(n9165), .ZN(N6193) );
  AOI22D1BWP30P140LVT U13477 ( .A1(i_data_bus[116]), .A2(n10549), .B1(
        i_data_bus[20]), .B2(n10552), .ZN(n9168) );
  AOI22D1BWP30P140LVT U13478 ( .A1(i_data_bus[52]), .A2(n10550), .B1(
        i_data_bus[84]), .B2(n10551), .ZN(n9167) );
  ND2D1BWP30P140LVT U13479 ( .A1(n9168), .A2(n9167), .ZN(N6213) );
  AOI22D1BWP30P140LVT U13480 ( .A1(i_data_bus[17]), .A2(n10552), .B1(
        i_data_bus[113]), .B2(n10549), .ZN(n9170) );
  AOI22D1BWP30P140LVT U13481 ( .A1(i_data_bus[49]), .A2(n10550), .B1(
        i_data_bus[81]), .B2(n10551), .ZN(n9169) );
  ND2D1BWP30P140LVT U13482 ( .A1(n9170), .A2(n9169), .ZN(N6210) );
  AOI22D1BWP30P140LVT U13483 ( .A1(i_data_bus[100]), .A2(n10549), .B1(
        i_data_bus[36]), .B2(n10550), .ZN(n9172) );
  AOI22D1BWP30P140LVT U13484 ( .A1(i_data_bus[4]), .A2(n10552), .B1(
        i_data_bus[68]), .B2(n10551), .ZN(n9171) );
  ND2D1BWP30P140LVT U13485 ( .A1(n9172), .A2(n9171), .ZN(N6197) );
  AOI22D1BWP30P140LVT U13486 ( .A1(i_data_bus[14]), .A2(n10552), .B1(
        i_data_bus[46]), .B2(n10550), .ZN(n9174) );
  AOI22D1BWP30P140LVT U13487 ( .A1(i_data_bus[110]), .A2(n10549), .B1(
        i_data_bus[78]), .B2(n10551), .ZN(n9173) );
  ND2D1BWP30P140LVT U13488 ( .A1(n9174), .A2(n9173), .ZN(N6207) );
  AOI22D1BWP30P140LVT U13489 ( .A1(i_data_bus[123]), .A2(n10549), .B1(
        i_data_bus[59]), .B2(n10550), .ZN(n9176) );
  AOI22D1BWP30P140LVT U13490 ( .A1(i_data_bus[27]), .A2(n10552), .B1(
        i_data_bus[91]), .B2(n10551), .ZN(n9175) );
  ND2D1BWP30P140LVT U13491 ( .A1(n9176), .A2(n9175), .ZN(N6220) );
  AOI22D1BWP30P140LVT U13492 ( .A1(i_data_bus[117]), .A2(n10549), .B1(
        i_data_bus[21]), .B2(n10552), .ZN(n9178) );
  AOI22D1BWP30P140LVT U13493 ( .A1(i_data_bus[53]), .A2(n10550), .B1(
        i_data_bus[85]), .B2(n10551), .ZN(n9177) );
  ND2D1BWP30P140LVT U13494 ( .A1(n9178), .A2(n9177), .ZN(N6214) );
  AOI22D1BWP30P140LVT U13495 ( .A1(i_data_bus[30]), .A2(n10552), .B1(
        i_data_bus[62]), .B2(n10550), .ZN(n9180) );
  AOI22D1BWP30P140LVT U13496 ( .A1(i_data_bus[126]), .A2(n10549), .B1(
        i_data_bus[94]), .B2(n10551), .ZN(n9179) );
  ND2D1BWP30P140LVT U13497 ( .A1(n9180), .A2(n9179), .ZN(N6223) );
  AOI22D1BWP30P140LVT U13498 ( .A1(i_data_bus[33]), .A2(n10550), .B1(
        i_data_bus[1]), .B2(n10552), .ZN(n9182) );
  AOI22D1BWP30P140LVT U13499 ( .A1(i_data_bus[97]), .A2(n10549), .B1(
        i_data_bus[65]), .B2(n10551), .ZN(n9181) );
  ND2D1BWP30P140LVT U13500 ( .A1(n9182), .A2(n9181), .ZN(N6194) );
  AOI22D1BWP30P140LVT U13501 ( .A1(i_data_bus[265]), .A2(n10510), .B1(
        i_data_bus[329]), .B2(n10509), .ZN(n9184) );
  AOI22D1BWP30P140LVT U13502 ( .A1(i_data_bus[297]), .A2(n10512), .B1(
        i_data_bus[361]), .B2(n10511), .ZN(n9183) );
  ND2D1BWP30P140LVT U13503 ( .A1(n9184), .A2(n9183), .ZN(N8508) );
  AOI22D1BWP30P140LVT U13504 ( .A1(i_data_bus[295]), .A2(n10512), .B1(
        i_data_bus[263]), .B2(n10510), .ZN(n9186) );
  AOI22D1BWP30P140LVT U13505 ( .A1(i_data_bus[327]), .A2(n10509), .B1(
        i_data_bus[359]), .B2(n10511), .ZN(n9185) );
  ND2D1BWP30P140LVT U13506 ( .A1(n9186), .A2(n9185), .ZN(N8506) );
  AOI22D1BWP30P140LVT U13507 ( .A1(i_data_bus[305]), .A2(n10512), .B1(
        i_data_bus[337]), .B2(n10509), .ZN(n9188) );
  AOI22D1BWP30P140LVT U13508 ( .A1(i_data_bus[273]), .A2(n10510), .B1(
        i_data_bus[369]), .B2(n10511), .ZN(n9187) );
  ND2D1BWP30P140LVT U13509 ( .A1(n9188), .A2(n9187), .ZN(N8516) );
  AOI22D1BWP30P140LVT U13510 ( .A1(i_data_bus[347]), .A2(n10509), .B1(
        i_data_bus[283]), .B2(n10510), .ZN(n9190) );
  AOI22D1BWP30P140LVT U13511 ( .A1(i_data_bus[315]), .A2(n10512), .B1(
        i_data_bus[379]), .B2(n10511), .ZN(n9189) );
  ND2D1BWP30P140LVT U13512 ( .A1(n9190), .A2(n9189), .ZN(N8526) );
  AOI22D1BWP30P140LVT U13513 ( .A1(i_data_bus[266]), .A2(n10510), .B1(
        i_data_bus[330]), .B2(n10509), .ZN(n9192) );
  AOI22D1BWP30P140LVT U13514 ( .A1(i_data_bus[298]), .A2(n10512), .B1(
        i_data_bus[362]), .B2(n10511), .ZN(n9191) );
  ND2D1BWP30P140LVT U13515 ( .A1(n9192), .A2(n9191), .ZN(N8509) );
  AOI22D1BWP30P140LVT U13516 ( .A1(i_data_bus[292]), .A2(n10512), .B1(
        i_data_bus[260]), .B2(n10510), .ZN(n9194) );
  AOI22D1BWP30P140LVT U13517 ( .A1(i_data_bus[324]), .A2(n10509), .B1(
        i_data_bus[356]), .B2(n10511), .ZN(n9193) );
  ND2D1BWP30P140LVT U13518 ( .A1(n9194), .A2(n9193), .ZN(N8503) );
  AOI22D1BWP30P140LVT U13519 ( .A1(i_data_bus[351]), .A2(n10509), .B1(
        i_data_bus[319]), .B2(n10512), .ZN(n9196) );
  AOI22D1BWP30P140LVT U13520 ( .A1(i_data_bus[287]), .A2(n10510), .B1(
        i_data_bus[383]), .B2(n10511), .ZN(n9195) );
  ND2D1BWP30P140LVT U13521 ( .A1(n9196), .A2(n9195), .ZN(N8530) );
  AOI22D1BWP30P140LVT U13522 ( .A1(i_data_bus[310]), .A2(n10512), .B1(
        i_data_bus[342]), .B2(n10509), .ZN(n9198) );
  AOI22D1BWP30P140LVT U13523 ( .A1(i_data_bus[278]), .A2(n10510), .B1(
        i_data_bus[374]), .B2(n10511), .ZN(n9197) );
  ND2D1BWP30P140LVT U13524 ( .A1(n9198), .A2(n9197), .ZN(N8521) );
  AOI22D1BWP30P140LVT U13525 ( .A1(i_data_bus[48]), .A2(n10583), .B1(
        i_data_bus[112]), .B2(n10584), .ZN(n9200) );
  AOI22D1BWP30P140LVT U13526 ( .A1(i_data_bus[80]), .A2(n10582), .B1(
        i_data_bus[16]), .B2(n10581), .ZN(n9199) );
  ND2D1BWP30P140LVT U13527 ( .A1(n9200), .A2(n9199), .ZN(N4335) );
  AOI22D1BWP30P140LVT U13528 ( .A1(i_data_bus[127]), .A2(n10584), .B1(
        i_data_bus[63]), .B2(n10583), .ZN(n9202) );
  AOI22D1BWP30P140LVT U13529 ( .A1(i_data_bus[95]), .A2(n10582), .B1(
        i_data_bus[31]), .B2(n10581), .ZN(n9201) );
  ND2D1BWP30P140LVT U13530 ( .A1(n9202), .A2(n9201), .ZN(N4350) );
  AOI22D1BWP30P140LVT U13531 ( .A1(i_data_bus[118]), .A2(n10584), .B1(
        i_data_bus[86]), .B2(n10582), .ZN(n9204) );
  AOI22D1BWP30P140LVT U13532 ( .A1(i_data_bus[54]), .A2(n10583), .B1(
        i_data_bus[22]), .B2(n10581), .ZN(n9203) );
  ND2D1BWP30P140LVT U13533 ( .A1(n9204), .A2(n9203), .ZN(N4341) );
  AOI22D1BWP30P140LVT U13534 ( .A1(i_data_bus[90]), .A2(n10582), .B1(
        i_data_bus[58]), .B2(n10583), .ZN(n9206) );
  AOI22D1BWP30P140LVT U13535 ( .A1(i_data_bus[122]), .A2(n10584), .B1(
        i_data_bus[26]), .B2(n10581), .ZN(n9205) );
  ND2D1BWP30P140LVT U13536 ( .A1(n9206), .A2(n9205), .ZN(N4345) );
  AOI22D1BWP30P140LVT U13537 ( .A1(i_data_bus[52]), .A2(n10583), .B1(
        i_data_bus[116]), .B2(n10584), .ZN(n9208) );
  AOI22D1BWP30P140LVT U13538 ( .A1(i_data_bus[84]), .A2(n10582), .B1(
        i_data_bus[20]), .B2(n10581), .ZN(n9207) );
  ND2D1BWP30P140LVT U13539 ( .A1(n9208), .A2(n9207), .ZN(N4339) );
  AOI22D1BWP30P140LVT U13540 ( .A1(i_data_bus[104]), .A2(n10584), .B1(
        i_data_bus[72]), .B2(n10582), .ZN(n9210) );
  AOI22D1BWP30P140LVT U13541 ( .A1(i_data_bus[40]), .A2(n10583), .B1(
        i_data_bus[8]), .B2(n10581), .ZN(n9209) );
  ND2D1BWP30P140LVT U13542 ( .A1(n9210), .A2(n9209), .ZN(N4327) );
  AOI22D1BWP30P140LVT U13543 ( .A1(i_data_bus[44]), .A2(n10583), .B1(
        i_data_bus[108]), .B2(n10584), .ZN(n9212) );
  AOI22D1BWP30P140LVT U13544 ( .A1(i_data_bus[76]), .A2(n10582), .B1(
        i_data_bus[12]), .B2(n10581), .ZN(n9211) );
  ND2D1BWP30P140LVT U13545 ( .A1(n9212), .A2(n9211), .ZN(N4331) );
  AOI22D1BWP30P140LVT U13546 ( .A1(i_data_bus[51]), .A2(n10583), .B1(
        i_data_bus[115]), .B2(n10584), .ZN(n9214) );
  AOI22D1BWP30P140LVT U13547 ( .A1(i_data_bus[83]), .A2(n10582), .B1(
        i_data_bus[19]), .B2(n10581), .ZN(n9213) );
  ND2D1BWP30P140LVT U13548 ( .A1(n9214), .A2(n9213), .ZN(N4338) );
  AOI22D1BWP30P140LVT U13549 ( .A1(i_data_bus[98]), .A2(n10584), .B1(
        i_data_bus[34]), .B2(n10583), .ZN(n9216) );
  AOI22D1BWP30P140LVT U13550 ( .A1(i_data_bus[66]), .A2(n10582), .B1(
        i_data_bus[2]), .B2(n10581), .ZN(n9215) );
  ND2D1BWP30P140LVT U13551 ( .A1(n9216), .A2(n9215), .ZN(N4321) );
  AOI22D1BWP30P140LVT U13552 ( .A1(i_data_bus[75]), .A2(n10582), .B1(
        i_data_bus[107]), .B2(n10584), .ZN(n9218) );
  AOI22D1BWP30P140LVT U13553 ( .A1(i_data_bus[43]), .A2(n10583), .B1(
        i_data_bus[11]), .B2(n10581), .ZN(n9217) );
  ND2D1BWP30P140LVT U13554 ( .A1(n9218), .A2(n9217), .ZN(N4330) );
  AOI22D1BWP30P140LVT U13555 ( .A1(i_data_bus[862]), .A2(n10399), .B1(
        i_data_bus[894]), .B2(n10398), .ZN(n9220) );
  AOI22D1BWP30P140LVT U13556 ( .A1(i_data_bus[798]), .A2(n10397), .B1(
        i_data_bus[830]), .B2(n10400), .ZN(n9219) );
  ND2D1BWP30P140LVT U13557 ( .A1(n9220), .A2(n9219), .ZN(N15015) );
  AOI22D1BWP30P140LVT U13558 ( .A1(i_data_bus[796]), .A2(n10397), .B1(
        i_data_bus[892]), .B2(n10398), .ZN(n9222) );
  AOI22D1BWP30P140LVT U13559 ( .A1(i_data_bus[860]), .A2(n10399), .B1(
        i_data_bus[828]), .B2(n10400), .ZN(n9221) );
  ND2D1BWP30P140LVT U13560 ( .A1(n9222), .A2(n9221), .ZN(N15013) );
  AOI22D1BWP30P140LVT U13561 ( .A1(i_data_bus[889]), .A2(n10398), .B1(
        i_data_bus[793]), .B2(n10397), .ZN(n9224) );
  AOI22D1BWP30P140LVT U13562 ( .A1(i_data_bus[857]), .A2(n10399), .B1(
        i_data_bus[825]), .B2(n10400), .ZN(n9223) );
  ND2D1BWP30P140LVT U13563 ( .A1(n9224), .A2(n9223), .ZN(N15010) );
  AOI22D1BWP30P140LVT U13564 ( .A1(i_data_bus[841]), .A2(n10399), .B1(
        i_data_bus[873]), .B2(n10398), .ZN(n9226) );
  AOI22D1BWP30P140LVT U13565 ( .A1(i_data_bus[777]), .A2(n10397), .B1(
        i_data_bus[809]), .B2(n10400), .ZN(n9225) );
  ND2D1BWP30P140LVT U13566 ( .A1(n9226), .A2(n9225), .ZN(N14994) );
  AOI22D1BWP30P140LVT U13567 ( .A1(i_data_bus[855]), .A2(n10399), .B1(
        i_data_bus[791]), .B2(n10397), .ZN(n9228) );
  AOI22D1BWP30P140LVT U13568 ( .A1(i_data_bus[887]), .A2(n10398), .B1(
        i_data_bus[823]), .B2(n10400), .ZN(n9227) );
  ND2D1BWP30P140LVT U13569 ( .A1(n9228), .A2(n9227), .ZN(N15008) );
  AOI22D1BWP30P140LVT U13570 ( .A1(i_data_bus[849]), .A2(n10399), .B1(
        i_data_bus[785]), .B2(n10397), .ZN(n9230) );
  AOI22D1BWP30P140LVT U13571 ( .A1(i_data_bus[881]), .A2(n10398), .B1(
        i_data_bus[817]), .B2(n10400), .ZN(n9229) );
  ND2D1BWP30P140LVT U13572 ( .A1(n9230), .A2(n9229), .ZN(N15002) );
  AOI22D1BWP30P140LVT U13573 ( .A1(i_data_bus[768]), .A2(n10397), .B1(
        i_data_bus[864]), .B2(n10398), .ZN(n9232) );
  AOI22D1BWP30P140LVT U13574 ( .A1(i_data_bus[832]), .A2(n10399), .B1(
        i_data_bus[800]), .B2(n10400), .ZN(n9231) );
  ND2D1BWP30P140LVT U13575 ( .A1(n9232), .A2(n9231), .ZN(N14985) );
  AOI22D1BWP30P140LVT U13576 ( .A1(i_data_bus[834]), .A2(n10399), .B1(
        i_data_bus[770]), .B2(n10397), .ZN(n9234) );
  AOI22D1BWP30P140LVT U13577 ( .A1(i_data_bus[866]), .A2(n10398), .B1(
        i_data_bus[802]), .B2(n10400), .ZN(n9233) );
  ND2D1BWP30P140LVT U13578 ( .A1(n9234), .A2(n9233), .ZN(N14987) );
  AOI22D1BWP30P140LVT U13579 ( .A1(i_data_bus[553]), .A2(n10406), .B1(
        i_data_bus[585]), .B2(n10408), .ZN(n9236) );
  AOI22D1BWP30P140LVT U13580 ( .A1(i_data_bus[521]), .A2(n10405), .B1(
        i_data_bus[617]), .B2(n10407), .ZN(n9235) );
  ND2D1BWP30P140LVT U13581 ( .A1(n9236), .A2(n9235), .ZN(N14562) );
  AOI22D1BWP30P140LVT U13582 ( .A1(i_data_bus[548]), .A2(n10406), .B1(
        i_data_bus[580]), .B2(n10408), .ZN(n9238) );
  AOI22D1BWP30P140LVT U13583 ( .A1(i_data_bus[516]), .A2(n10405), .B1(
        i_data_bus[612]), .B2(n10407), .ZN(n9237) );
  ND2D1BWP30P140LVT U13584 ( .A1(n9238), .A2(n9237), .ZN(N14557) );
  AOI22D1BWP30P140LVT U13585 ( .A1(i_data_bus[551]), .A2(n10406), .B1(
        i_data_bus[583]), .B2(n10408), .ZN(n9240) );
  AOI22D1BWP30P140LVT U13586 ( .A1(i_data_bus[519]), .A2(n10405), .B1(
        i_data_bus[615]), .B2(n10407), .ZN(n9239) );
  ND2D1BWP30P140LVT U13587 ( .A1(n9240), .A2(n9239), .ZN(N14560) );
  AOI22D1BWP30P140LVT U13588 ( .A1(i_data_bus[543]), .A2(n10405), .B1(
        i_data_bus[575]), .B2(n10406), .ZN(n9242) );
  AOI22D1BWP30P140LVT U13589 ( .A1(i_data_bus[607]), .A2(n10408), .B1(
        i_data_bus[639]), .B2(n10407), .ZN(n9241) );
  ND2D1BWP30P140LVT U13590 ( .A1(n9242), .A2(n9241), .ZN(N14584) );
  AOI22D1BWP30P140LVT U13591 ( .A1(i_data_bus[587]), .A2(n10408), .B1(
        i_data_bus[555]), .B2(n10406), .ZN(n9244) );
  AOI22D1BWP30P140LVT U13592 ( .A1(i_data_bus[523]), .A2(n10405), .B1(
        i_data_bus[619]), .B2(n10407), .ZN(n9243) );
  ND2D1BWP30P140LVT U13593 ( .A1(n9244), .A2(n9243), .ZN(N14564) );
  AOI22D1BWP30P140LVT U13594 ( .A1(i_data_bus[601]), .A2(n10408), .B1(
        i_data_bus[569]), .B2(n10406), .ZN(n9246) );
  AOI22D1BWP30P140LVT U13595 ( .A1(i_data_bus[537]), .A2(n10405), .B1(
        i_data_bus[633]), .B2(n10407), .ZN(n9245) );
  ND2D1BWP30P140LVT U13596 ( .A1(n9246), .A2(n9245), .ZN(N14578) );
  AOI22D1BWP30P140LVT U13597 ( .A1(i_data_bus[722]), .A2(n10497), .B1(
        i_data_bus[690]), .B2(n10499), .ZN(n9248) );
  AOI22D1BWP30P140LVT U13598 ( .A1(i_data_bus[658]), .A2(n10498), .B1(
        i_data_bus[754]), .B2(n10500), .ZN(n9247) );
  ND2D1BWP30P140LVT U13599 ( .A1(n9248), .A2(n9247), .ZN(N9165) );
  AOI22D1BWP30P140LVT U13600 ( .A1(i_data_bus[679]), .A2(n10499), .B1(
        i_data_bus[647]), .B2(n10498), .ZN(n9250) );
  AOI22D1BWP30P140LVT U13601 ( .A1(i_data_bus[711]), .A2(n10497), .B1(
        i_data_bus[743]), .B2(n10500), .ZN(n9249) );
  ND2D1BWP30P140LVT U13602 ( .A1(n9250), .A2(n9249), .ZN(N9154) );
  AOI22D1BWP30P140LVT U13603 ( .A1(i_data_bus[686]), .A2(n10499), .B1(
        i_data_bus[654]), .B2(n10498), .ZN(n9252) );
  AOI22D1BWP30P140LVT U13604 ( .A1(i_data_bus[718]), .A2(n10497), .B1(
        i_data_bus[750]), .B2(n10500), .ZN(n9251) );
  ND2D1BWP30P140LVT U13605 ( .A1(n9252), .A2(n9251), .ZN(N9161) );
  AOI22D1BWP30P140LVT U13606 ( .A1(i_data_bus[700]), .A2(n10499), .B1(
        i_data_bus[668]), .B2(n10498), .ZN(n9254) );
  AOI22D1BWP30P140LVT U13607 ( .A1(i_data_bus[732]), .A2(n10497), .B1(
        i_data_bus[764]), .B2(n10500), .ZN(n9253) );
  ND2D1BWP30P140LVT U13608 ( .A1(n9254), .A2(n9253), .ZN(N9175) );
  AOI22D1BWP30P140LVT U13609 ( .A1(i_data_bus[728]), .A2(n10497), .B1(
        i_data_bus[664]), .B2(n10498), .ZN(n9256) );
  AOI22D1BWP30P140LVT U13610 ( .A1(i_data_bus[696]), .A2(n10499), .B1(
        i_data_bus[760]), .B2(n10500), .ZN(n9255) );
  ND2D1BWP30P140LVT U13611 ( .A1(n9256), .A2(n9255), .ZN(N9171) );
  AOI22D1BWP30P140LVT U13612 ( .A1(i_data_bus[715]), .A2(n10497), .B1(
        i_data_bus[683]), .B2(n10499), .ZN(n9258) );
  AOI22D1BWP30P140LVT U13613 ( .A1(i_data_bus[651]), .A2(n10498), .B1(
        i_data_bus[747]), .B2(n10500), .ZN(n9257) );
  ND2D1BWP30P140LVT U13614 ( .A1(n9258), .A2(n9257), .ZN(N9158) );
  AOI22D1BWP30P140LVT U13615 ( .A1(i_data_bus[726]), .A2(n10497), .B1(
        i_data_bus[662]), .B2(n10498), .ZN(n9260) );
  AOI22D1BWP30P140LVT U13616 ( .A1(i_data_bus[694]), .A2(n10499), .B1(
        i_data_bus[758]), .B2(n10500), .ZN(n9259) );
  ND2D1BWP30P140LVT U13617 ( .A1(n9260), .A2(n9259), .ZN(N9169) );
  AOI22D1BWP30P140LVT U13618 ( .A1(i_data_bus[704]), .A2(n10497), .B1(
        i_data_bus[640]), .B2(n10498), .ZN(n9262) );
  AOI22D1BWP30P140LVT U13619 ( .A1(i_data_bus[672]), .A2(n10499), .B1(
        i_data_bus[736]), .B2(n10500), .ZN(n9261) );
  ND2D1BWP30P140LVT U13620 ( .A1(n9262), .A2(n9261), .ZN(N9147) );
  AOI22D1BWP30P140LVT U13621 ( .A1(i_data_bus[642]), .A2(n10498), .B1(
        i_data_bus[674]), .B2(n10499), .ZN(n9264) );
  AOI22D1BWP30P140LVT U13622 ( .A1(i_data_bus[706]), .A2(n10497), .B1(
        i_data_bus[738]), .B2(n10500), .ZN(n9263) );
  ND2D1BWP30P140LVT U13623 ( .A1(n9264), .A2(n9263), .ZN(N9149) );
  AOI22D1BWP30P140LVT U13624 ( .A1(i_data_bus[673]), .A2(n10499), .B1(
        i_data_bus[705]), .B2(n10497), .ZN(n9266) );
  AOI22D1BWP30P140LVT U13625 ( .A1(i_data_bus[641]), .A2(n10498), .B1(
        i_data_bus[737]), .B2(n10500), .ZN(n9265) );
  ND2D1BWP30P140LVT U13626 ( .A1(n9266), .A2(n9265), .ZN(N9148) );
  AOI22D1BWP30P140LVT U13627 ( .A1(i_data_bus[253]), .A2(n10516), .B1(
        i_data_bus[221]), .B2(n10514), .ZN(n9268) );
  AOI22D1BWP30P140LVT U13628 ( .A1(i_data_bus[189]), .A2(n10515), .B1(
        i_data_bus[157]), .B2(n10513), .ZN(n9267) );
  ND2D1BWP30P140LVT U13629 ( .A1(n9268), .A2(n9267), .ZN(N8312) );
  AOI22D1BWP30P140LVT U13630 ( .A1(i_data_bus[216]), .A2(n10514), .B1(
        i_data_bus[184]), .B2(n10515), .ZN(n9270) );
  AOI22D1BWP30P140LVT U13631 ( .A1(i_data_bus[248]), .A2(n10516), .B1(
        i_data_bus[152]), .B2(n10513), .ZN(n9269) );
  ND2D1BWP30P140LVT U13632 ( .A1(n9270), .A2(n9269), .ZN(N8307) );
  AOI22D1BWP30P140LVT U13633 ( .A1(i_data_bus[204]), .A2(n10578), .B1(
        i_data_bus[172]), .B2(n10579), .ZN(n9272) );
  AOI22D1BWP30P140LVT U13634 ( .A1(i_data_bus[236]), .A2(n10580), .B1(
        i_data_bus[140]), .B2(n10577), .ZN(n9271) );
  ND2D1BWP30P140LVT U13635 ( .A1(n9272), .A2(n9271), .ZN(N4547) );
  AOI22D1BWP30P140LVT U13636 ( .A1(i_data_bus[207]), .A2(n10514), .B1(
        i_data_bus[239]), .B2(n10516), .ZN(n9274) );
  AOI22D1BWP30P140LVT U13637 ( .A1(i_data_bus[175]), .A2(n10515), .B1(
        i_data_bus[143]), .B2(n10513), .ZN(n9273) );
  ND2D1BWP30P140LVT U13638 ( .A1(n9274), .A2(n9273), .ZN(N8298) );
  AOI22D1BWP30P140LVT U13639 ( .A1(i_data_bus[198]), .A2(n10578), .B1(
        i_data_bus[166]), .B2(n10579), .ZN(n9276) );
  AOI22D1BWP30P140LVT U13640 ( .A1(i_data_bus[230]), .A2(n10580), .B1(
        i_data_bus[134]), .B2(n10577), .ZN(n9275) );
  ND2D1BWP30P140LVT U13641 ( .A1(n9276), .A2(n9275), .ZN(N4541) );
  AOI22D1BWP30P140LVT U13642 ( .A1(i_data_bus[255]), .A2(n10580), .B1(
        i_data_bus[191]), .B2(n10579), .ZN(n9278) );
  AOI22D1BWP30P140LVT U13643 ( .A1(i_data_bus[223]), .A2(n10578), .B1(
        i_data_bus[159]), .B2(n10577), .ZN(n9277) );
  ND2D1BWP30P140LVT U13644 ( .A1(n9278), .A2(n9277), .ZN(N4566) );
  AOI22D1BWP30P140LVT U13645 ( .A1(i_data_bus[163]), .A2(n10515), .B1(
        i_data_bus[195]), .B2(n10514), .ZN(n9280) );
  AOI22D1BWP30P140LVT U13646 ( .A1(i_data_bus[227]), .A2(n10516), .B1(
        i_data_bus[131]), .B2(n10513), .ZN(n9279) );
  ND2D1BWP30P140LVT U13647 ( .A1(n9280), .A2(n9279), .ZN(N8286) );
  AOI22D1BWP30P140LVT U13648 ( .A1(i_data_bus[215]), .A2(n10578), .B1(
        i_data_bus[247]), .B2(n10580), .ZN(n9282) );
  AOI22D1BWP30P140LVT U13649 ( .A1(i_data_bus[183]), .A2(n10579), .B1(
        i_data_bus[151]), .B2(n10577), .ZN(n9281) );
  ND2D1BWP30P140LVT U13650 ( .A1(n9282), .A2(n9281), .ZN(N4558) );
  AOI22D1BWP30P140LVT U13651 ( .A1(i_data_bus[170]), .A2(n10515), .B1(
        i_data_bus[202]), .B2(n10514), .ZN(n9284) );
  AOI22D1BWP30P140LVT U13652 ( .A1(i_data_bus[234]), .A2(n10516), .B1(
        i_data_bus[138]), .B2(n10513), .ZN(n9283) );
  ND2D1BWP30P140LVT U13653 ( .A1(n9284), .A2(n9283), .ZN(N8293) );
  AOI22D1BWP30P140LVT U13654 ( .A1(i_data_bus[251]), .A2(n10516), .B1(
        i_data_bus[219]), .B2(n10514), .ZN(n9286) );
  AOI22D1BWP30P140LVT U13655 ( .A1(i_data_bus[187]), .A2(n10515), .B1(
        i_data_bus[155]), .B2(n10513), .ZN(n9285) );
  ND2D1BWP30P140LVT U13656 ( .A1(n9286), .A2(n9285), .ZN(N8310) );
  AOI22D1BWP30P140LVT U13657 ( .A1(i_data_bus[177]), .A2(n10579), .B1(
        i_data_bus[241]), .B2(n10580), .ZN(n9288) );
  AOI22D1BWP30P140LVT U13658 ( .A1(i_data_bus[209]), .A2(n10578), .B1(
        i_data_bus[145]), .B2(n10577), .ZN(n9287) );
  ND2D1BWP30P140LVT U13659 ( .A1(n9288), .A2(n9287), .ZN(N4552) );
  AOI22D1BWP30P140LVT U13660 ( .A1(i_data_bus[235]), .A2(n10516), .B1(
        i_data_bus[171]), .B2(n10515), .ZN(n9290) );
  AOI22D1BWP30P140LVT U13661 ( .A1(i_data_bus[203]), .A2(n10514), .B1(
        i_data_bus[139]), .B2(n10513), .ZN(n9289) );
  ND2D1BWP30P140LVT U13662 ( .A1(n9290), .A2(n9289), .ZN(N8294) );
  AOI22D1BWP30P140LVT U13663 ( .A1(i_data_bus[177]), .A2(n10515), .B1(
        i_data_bus[241]), .B2(n10516), .ZN(n9292) );
  AOI22D1BWP30P140LVT U13664 ( .A1(i_data_bus[209]), .A2(n10514), .B1(
        i_data_bus[145]), .B2(n10513), .ZN(n9291) );
  ND2D1BWP30P140LVT U13665 ( .A1(n9292), .A2(n9291), .ZN(N8300) );
  AOI22D1BWP30P140LVT U13666 ( .A1(i_data_bus[234]), .A2(n10580), .B1(
        i_data_bus[202]), .B2(n10578), .ZN(n9294) );
  AOI22D1BWP30P140LVT U13667 ( .A1(i_data_bus[170]), .A2(n10579), .B1(
        i_data_bus[138]), .B2(n10577), .ZN(n9293) );
  ND2D1BWP30P140LVT U13668 ( .A1(n9294), .A2(n9293), .ZN(N4545) );
  AOI22D1BWP30P140LVT U13669 ( .A1(i_data_bus[194]), .A2(n10514), .B1(
        i_data_bus[226]), .B2(n10516), .ZN(n9296) );
  AOI22D1BWP30P140LVT U13670 ( .A1(i_data_bus[162]), .A2(n10515), .B1(
        i_data_bus[130]), .B2(n10513), .ZN(n9295) );
  ND2D1BWP30P140LVT U13671 ( .A1(n9296), .A2(n9295), .ZN(N8285) );
  AOI22D1BWP30P140LVT U13672 ( .A1(i_data_bus[175]), .A2(n10579), .B1(
        i_data_bus[239]), .B2(n10580), .ZN(n9298) );
  AOI22D1BWP30P140LVT U13673 ( .A1(i_data_bus[207]), .A2(n10578), .B1(
        i_data_bus[143]), .B2(n10577), .ZN(n9297) );
  ND2D1BWP30P140LVT U13674 ( .A1(n9298), .A2(n9297), .ZN(N4550) );
  AOI22D1BWP30P140LVT U13675 ( .A1(i_data_bus[238]), .A2(n10580), .B1(
        i_data_bus[206]), .B2(n10578), .ZN(n9300) );
  AOI22D1BWP30P140LVT U13676 ( .A1(i_data_bus[174]), .A2(n10579), .B1(
        i_data_bus[142]), .B2(n10577), .ZN(n9299) );
  ND2D1BWP30P140LVT U13677 ( .A1(n9300), .A2(n9299), .ZN(N4549) );
  AOI22D1BWP30P140LVT U13678 ( .A1(i_data_bus[201]), .A2(n10578), .B1(
        i_data_bus[169]), .B2(n10579), .ZN(n9302) );
  AOI22D1BWP30P140LVT U13679 ( .A1(i_data_bus[233]), .A2(n10580), .B1(
        i_data_bus[137]), .B2(n10577), .ZN(n9301) );
  ND2D1BWP30P140LVT U13680 ( .A1(n9302), .A2(n9301), .ZN(N4544) );
  AOI22D1BWP30P140LVT U13681 ( .A1(i_data_bus[198]), .A2(n10514), .B1(
        i_data_bus[230]), .B2(n10516), .ZN(n9304) );
  AOI22D1BWP30P140LVT U13682 ( .A1(i_data_bus[166]), .A2(n10515), .B1(
        i_data_bus[134]), .B2(n10513), .ZN(n9303) );
  ND2D1BWP30P140LVT U13683 ( .A1(n9304), .A2(n9303), .ZN(N8289) );
  AOI22D1BWP30P140LVT U13684 ( .A1(i_data_bus[162]), .A2(n10579), .B1(
        i_data_bus[226]), .B2(n10580), .ZN(n9306) );
  AOI22D1BWP30P140LVT U13685 ( .A1(i_data_bus[194]), .A2(n10578), .B1(
        i_data_bus[130]), .B2(n10577), .ZN(n9305) );
  ND2D1BWP30P140LVT U13686 ( .A1(n9306), .A2(n9305), .ZN(N4537) );
  AOI22D1BWP30P140LVT U13687 ( .A1(i_data_bus[227]), .A2(n10580), .B1(
        i_data_bus[195]), .B2(n10578), .ZN(n9308) );
  AOI22D1BWP30P140LVT U13688 ( .A1(i_data_bus[163]), .A2(n10579), .B1(
        i_data_bus[131]), .B2(n10577), .ZN(n9307) );
  ND2D1BWP30P140LVT U13689 ( .A1(n9308), .A2(n9307), .ZN(N4538) );
  AOI22D1BWP30P140LVT U13690 ( .A1(i_data_bus[214]), .A2(n10578), .B1(
        i_data_bus[246]), .B2(n10580), .ZN(n9310) );
  AOI22D1BWP30P140LVT U13691 ( .A1(i_data_bus[182]), .A2(n10579), .B1(
        i_data_bus[150]), .B2(n10577), .ZN(n9309) );
  ND2D1BWP30P140LVT U13692 ( .A1(n9310), .A2(n9309), .ZN(N4557) );
  AOI22D1BWP30P140LVT U13693 ( .A1(i_data_bus[255]), .A2(n10516), .B1(
        i_data_bus[191]), .B2(n10515), .ZN(n9312) );
  AOI22D1BWP30P140LVT U13694 ( .A1(i_data_bus[223]), .A2(n10514), .B1(
        i_data_bus[159]), .B2(n10513), .ZN(n9311) );
  ND2D1BWP30P140LVT U13695 ( .A1(n9312), .A2(n9311), .ZN(N8314) );
  AOI22D1BWP30P140LVT U13696 ( .A1(i_data_bus[952]), .A2(n10428), .B1(
        i_data_bus[920]), .B2(n10425), .ZN(n9314) );
  AOI22D1BWP30P140LVT U13697 ( .A1(i_data_bus[1016]), .A2(n10427), .B1(
        i_data_bus[984]), .B2(n10426), .ZN(n9313) );
  ND2D1BWP30P140LVT U13698 ( .A1(n9314), .A2(n9313), .ZN(N13351) );
  AOI22D1BWP30P140LVT U13699 ( .A1(i_data_bus[929]), .A2(n10428), .B1(
        i_data_bus[897]), .B2(n10425), .ZN(n9316) );
  AOI22D1BWP30P140LVT U13700 ( .A1(i_data_bus[993]), .A2(n10427), .B1(
        i_data_bus[961]), .B2(n10426), .ZN(n9315) );
  ND2D1BWP30P140LVT U13701 ( .A1(n9316), .A2(n9315), .ZN(N13328) );
  AOI22D1BWP30P140LVT U13702 ( .A1(i_data_bus[919]), .A2(n10425), .B1(
        i_data_bus[1015]), .B2(n10427), .ZN(n9318) );
  AOI22D1BWP30P140LVT U13703 ( .A1(i_data_bus[951]), .A2(n10428), .B1(
        i_data_bus[983]), .B2(n10426), .ZN(n9317) );
  ND2D1BWP30P140LVT U13704 ( .A1(n9318), .A2(n9317), .ZN(N13350) );
  AOI22D1BWP30P140LVT U13705 ( .A1(i_data_bus[923]), .A2(n10425), .B1(
        i_data_bus[1019]), .B2(n10427), .ZN(n9320) );
  AOI22D1BWP30P140LVT U13706 ( .A1(i_data_bus[955]), .A2(n10428), .B1(
        i_data_bus[987]), .B2(n10426), .ZN(n9319) );
  ND2D1BWP30P140LVT U13707 ( .A1(n9320), .A2(n9319), .ZN(N13354) );
  AOI22D1BWP30P140LVT U13708 ( .A1(i_data_bus[1011]), .A2(n10427), .B1(
        i_data_bus[915]), .B2(n10425), .ZN(n9322) );
  AOI22D1BWP30P140LVT U13709 ( .A1(i_data_bus[947]), .A2(n10428), .B1(
        i_data_bus[979]), .B2(n10426), .ZN(n9321) );
  ND2D1BWP30P140LVT U13710 ( .A1(n9322), .A2(n9321), .ZN(N13346) );
  AOI22D1BWP30P140LVT U13711 ( .A1(i_data_bus[17]), .A2(n10486), .B1(
        i_data_bus[113]), .B2(n10488), .ZN(n9324) );
  AOI22D1BWP30P140LVT U13712 ( .A1(i_data_bus[49]), .A2(n10485), .B1(
        i_data_bus[81]), .B2(n10487), .ZN(n9323) );
  ND2D1BWP30P140LVT U13713 ( .A1(n9324), .A2(n9323), .ZN(N9958) );
  AOI22D1BWP30P140LVT U13714 ( .A1(i_data_bus[124]), .A2(n10488), .B1(
        i_data_bus[28]), .B2(n10486), .ZN(n9326) );
  AOI22D1BWP30P140LVT U13715 ( .A1(i_data_bus[60]), .A2(n10485), .B1(
        i_data_bus[92]), .B2(n10487), .ZN(n9325) );
  ND2D1BWP30P140LVT U13716 ( .A1(n9326), .A2(n9325), .ZN(N9969) );
  AOI22D1BWP30P140LVT U13717 ( .A1(i_data_bus[100]), .A2(n10488), .B1(
        i_data_bus[36]), .B2(n10485), .ZN(n9328) );
  AOI22D1BWP30P140LVT U13718 ( .A1(i_data_bus[4]), .A2(n10486), .B1(
        i_data_bus[68]), .B2(n10487), .ZN(n9327) );
  ND2D1BWP30P140LVT U13719 ( .A1(n9328), .A2(n9327), .ZN(N9945) );
  AOI22D1BWP30P140LVT U13720 ( .A1(i_data_bus[115]), .A2(n10488), .B1(
        i_data_bus[19]), .B2(n10486), .ZN(n9330) );
  AOI22D1BWP30P140LVT U13721 ( .A1(i_data_bus[51]), .A2(n10485), .B1(
        i_data_bus[83]), .B2(n10487), .ZN(n9329) );
  ND2D1BWP30P140LVT U13722 ( .A1(n9330), .A2(n9329), .ZN(N9960) );
  AOI22D1BWP30P140LVT U13723 ( .A1(i_data_bus[38]), .A2(n10485), .B1(
        i_data_bus[102]), .B2(n10488), .ZN(n9332) );
  AOI22D1BWP30P140LVT U13724 ( .A1(i_data_bus[6]), .A2(n10486), .B1(
        i_data_bus[70]), .B2(n10487), .ZN(n9331) );
  ND2D1BWP30P140LVT U13725 ( .A1(n9332), .A2(n9331), .ZN(N9947) );
  AOI22D1BWP30P140LVT U13726 ( .A1(i_data_bus[45]), .A2(n10485), .B1(
        i_data_bus[13]), .B2(n10486), .ZN(n9334) );
  AOI22D1BWP30P140LVT U13727 ( .A1(i_data_bus[109]), .A2(n10488), .B1(
        i_data_bus[77]), .B2(n10487), .ZN(n9333) );
  ND2D1BWP30P140LVT U13728 ( .A1(n9334), .A2(n9333), .ZN(N9954) );
  AOI22D1BWP30P140LVT U13729 ( .A1(i_data_bus[32]), .A2(n10485), .B1(
        i_data_bus[0]), .B2(n10486), .ZN(n9336) );
  AOI22D1BWP30P140LVT U13730 ( .A1(i_data_bus[96]), .A2(n10488), .B1(
        i_data_bus[64]), .B2(n10487), .ZN(n9335) );
  ND2D1BWP30P140LVT U13731 ( .A1(n9336), .A2(n9335), .ZN(N9941) );
  AOI22D1BWP30P140LVT U13732 ( .A1(i_data_bus[123]), .A2(n10488), .B1(
        i_data_bus[59]), .B2(n10485), .ZN(n9338) );
  AOI22D1BWP30P140LVT U13733 ( .A1(i_data_bus[27]), .A2(n10486), .B1(
        i_data_bus[91]), .B2(n10487), .ZN(n9337) );
  ND2D1BWP30P140LVT U13734 ( .A1(n9338), .A2(n9337), .ZN(N9968) );
  AOI22D1BWP30P140LVT U13735 ( .A1(i_data_bus[14]), .A2(n10486), .B1(
        i_data_bus[110]), .B2(n10488), .ZN(n9340) );
  AOI22D1BWP30P140LVT U13736 ( .A1(i_data_bus[46]), .A2(n10485), .B1(
        i_data_bus[78]), .B2(n10487), .ZN(n9339) );
  ND2D1BWP30P140LVT U13737 ( .A1(n9340), .A2(n9339), .ZN(N9955) );
  AOI22D1BWP30P140LVT U13738 ( .A1(i_data_bus[30]), .A2(n10486), .B1(
        i_data_bus[62]), .B2(n10485), .ZN(n9342) );
  AOI22D1BWP30P140LVT U13739 ( .A1(i_data_bus[126]), .A2(n10488), .B1(
        i_data_bus[94]), .B2(n10487), .ZN(n9341) );
  ND2D1BWP30P140LVT U13740 ( .A1(n9342), .A2(n9341), .ZN(N9971) );
  AOI22D1BWP30P140LVT U13741 ( .A1(i_data_bus[116]), .A2(n10488), .B1(
        i_data_bus[20]), .B2(n10486), .ZN(n9344) );
  AOI22D1BWP30P140LVT U13742 ( .A1(i_data_bus[52]), .A2(n10485), .B1(
        i_data_bus[84]), .B2(n10487), .ZN(n9343) );
  ND2D1BWP30P140LVT U13743 ( .A1(n9344), .A2(n9343), .ZN(N9961) );
  AOI22D1BWP30P140LVT U13744 ( .A1(i_data_bus[838]), .A2(n10557), .B1(
        i_data_bus[774]), .B2(n10558), .ZN(n9346) );
  AOI22D1BWP30P140LVT U13745 ( .A1(i_data_bus[870]), .A2(n10559), .B1(
        i_data_bus[806]), .B2(n10560), .ZN(n9345) );
  ND2D1BWP30P140LVT U13746 ( .A1(n9346), .A2(n9345), .ZN(N5621) );
  AOI22D1BWP30P140LVT U13747 ( .A1(i_data_bus[889]), .A2(n10591), .B1(
        i_data_bus[793]), .B2(n10589), .ZN(n9348) );
  AOI22D1BWP30P140LVT U13748 ( .A1(i_data_bus[857]), .A2(n10590), .B1(
        i_data_bus[825]), .B2(n10592), .ZN(n9347) );
  ND2D1BWP30P140LVT U13749 ( .A1(n9348), .A2(n9347), .ZN(N3766) );
  AOI22D1BWP30P140LVT U13750 ( .A1(i_data_bus[840]), .A2(n10590), .B1(
        i_data_bus[776]), .B2(n10589), .ZN(n9350) );
  AOI22D1BWP30P140LVT U13751 ( .A1(i_data_bus[872]), .A2(n10591), .B1(
        i_data_bus[808]), .B2(n10592), .ZN(n9349) );
  ND2D1BWP30P140LVT U13752 ( .A1(n9350), .A2(n9349), .ZN(N3749) );
  AOI22D1BWP30P140LVT U13753 ( .A1(i_data_bus[771]), .A2(n10558), .B1(
        i_data_bus[835]), .B2(n10557), .ZN(n9352) );
  AOI22D1BWP30P140LVT U13754 ( .A1(i_data_bus[867]), .A2(n10559), .B1(
        i_data_bus[803]), .B2(n10560), .ZN(n9351) );
  ND2D1BWP30P140LVT U13755 ( .A1(n9352), .A2(n9351), .ZN(N5618) );
  AOI22D1BWP30P140LVT U13756 ( .A1(i_data_bus[783]), .A2(n10558), .B1(
        i_data_bus[879]), .B2(n10559), .ZN(n9354) );
  AOI22D1BWP30P140LVT U13757 ( .A1(i_data_bus[847]), .A2(n10557), .B1(
        i_data_bus[815]), .B2(n10560), .ZN(n9353) );
  ND2D1BWP30P140LVT U13758 ( .A1(n9354), .A2(n9353), .ZN(N5630) );
  AOI22D1BWP30P140LVT U13759 ( .A1(i_data_bus[866]), .A2(n10559), .B1(
        i_data_bus[770]), .B2(n10558), .ZN(n9356) );
  AOI22D1BWP30P140LVT U13760 ( .A1(i_data_bus[834]), .A2(n10557), .B1(
        i_data_bus[802]), .B2(n10560), .ZN(n9355) );
  ND2D1BWP30P140LVT U13761 ( .A1(n9356), .A2(n9355), .ZN(N5617) );
  AOI22D1BWP30P140LVT U13762 ( .A1(i_data_bus[843]), .A2(n10590), .B1(
        i_data_bus[875]), .B2(n10591), .ZN(n9358) );
  AOI22D1BWP30P140LVT U13763 ( .A1(i_data_bus[779]), .A2(n10589), .B1(
        i_data_bus[811]), .B2(n10592), .ZN(n9357) );
  ND2D1BWP30P140LVT U13764 ( .A1(n9358), .A2(n9357), .ZN(N3752) );
  AOI22D1BWP30P140LVT U13765 ( .A1(i_data_bus[841]), .A2(n10590), .B1(
        i_data_bus[873]), .B2(n10591), .ZN(n9360) );
  AOI22D1BWP30P140LVT U13766 ( .A1(i_data_bus[777]), .A2(n10589), .B1(
        i_data_bus[809]), .B2(n10592), .ZN(n9359) );
  ND2D1BWP30P140LVT U13767 ( .A1(n9360), .A2(n9359), .ZN(N3750) );
  AOI22D1BWP30P140LVT U13768 ( .A1(i_data_bus[771]), .A2(n10493), .B1(
        i_data_bus[835]), .B2(n10495), .ZN(n9362) );
  AOI22D1BWP30P140LVT U13769 ( .A1(i_data_bus[867]), .A2(n10494), .B1(
        i_data_bus[803]), .B2(n10496), .ZN(n9361) );
  ND2D1BWP30P140LVT U13770 ( .A1(n9362), .A2(n9361), .ZN(N9366) );
  AOI22D1BWP30P140LVT U13771 ( .A1(i_data_bus[860]), .A2(n10590), .B1(
        i_data_bus[892]), .B2(n10591), .ZN(n9364) );
  AOI22D1BWP30P140LVT U13772 ( .A1(i_data_bus[796]), .A2(n10589), .B1(
        i_data_bus[828]), .B2(n10592), .ZN(n9363) );
  ND2D1BWP30P140LVT U13773 ( .A1(n9364), .A2(n9363), .ZN(N3769) );
  AOI22D1BWP30P140LVT U13774 ( .A1(i_data_bus[778]), .A2(n10558), .B1(
        i_data_bus[874]), .B2(n10559), .ZN(n9366) );
  AOI22D1BWP30P140LVT U13775 ( .A1(i_data_bus[842]), .A2(n10557), .B1(
        i_data_bus[810]), .B2(n10560), .ZN(n9365) );
  ND2D1BWP30P140LVT U13776 ( .A1(n9366), .A2(n9365), .ZN(N5625) );
  AOI22D1BWP30P140LVT U13777 ( .A1(i_data_bus[848]), .A2(n10495), .B1(
        i_data_bus[880]), .B2(n10494), .ZN(n9368) );
  AOI22D1BWP30P140LVT U13778 ( .A1(i_data_bus[784]), .A2(n10493), .B1(
        i_data_bus[816]), .B2(n10496), .ZN(n9367) );
  ND2D1BWP30P140LVT U13779 ( .A1(n9368), .A2(n9367), .ZN(N9379) );
  AOI22D1BWP30P140LVT U13780 ( .A1(i_data_bus[775]), .A2(n10493), .B1(
        i_data_bus[839]), .B2(n10495), .ZN(n9370) );
  AOI22D1BWP30P140LVT U13781 ( .A1(i_data_bus[871]), .A2(n10494), .B1(
        i_data_bus[807]), .B2(n10496), .ZN(n9369) );
  ND2D1BWP30P140LVT U13782 ( .A1(n9370), .A2(n9369), .ZN(N9370) );
  AOI22D1BWP30P140LVT U13783 ( .A1(i_data_bus[779]), .A2(n10493), .B1(
        i_data_bus[875]), .B2(n10494), .ZN(n9372) );
  AOI22D1BWP30P140LVT U13784 ( .A1(i_data_bus[843]), .A2(n10495), .B1(
        i_data_bus[811]), .B2(n10496), .ZN(n9371) );
  ND2D1BWP30P140LVT U13785 ( .A1(n9372), .A2(n9371), .ZN(N9374) );
  AOI22D1BWP30P140LVT U13786 ( .A1(i_data_bus[881]), .A2(n10559), .B1(
        i_data_bus[849]), .B2(n10557), .ZN(n9374) );
  AOI22D1BWP30P140LVT U13787 ( .A1(i_data_bus[785]), .A2(n10558), .B1(
        i_data_bus[817]), .B2(n10560), .ZN(n9373) );
  ND2D1BWP30P140LVT U13788 ( .A1(n9374), .A2(n9373), .ZN(N5632) );
  AOI22D1BWP30P140LVT U13789 ( .A1(i_data_bus[858]), .A2(n10557), .B1(
        i_data_bus[890]), .B2(n10559), .ZN(n9376) );
  AOI22D1BWP30P140LVT U13790 ( .A1(i_data_bus[794]), .A2(n10558), .B1(
        i_data_bus[826]), .B2(n10560), .ZN(n9375) );
  ND2D1BWP30P140LVT U13791 ( .A1(n9376), .A2(n9375), .ZN(N5641) );
  AOI22D1BWP30P140LVT U13792 ( .A1(i_data_bus[783]), .A2(n10493), .B1(
        i_data_bus[847]), .B2(n10495), .ZN(n9378) );
  AOI22D1BWP30P140LVT U13793 ( .A1(i_data_bus[879]), .A2(n10494), .B1(
        i_data_bus[815]), .B2(n10496), .ZN(n9377) );
  ND2D1BWP30P140LVT U13794 ( .A1(n9378), .A2(n9377), .ZN(N9378) );
  AOI22D1BWP30P140LVT U13795 ( .A1(i_data_bus[862]), .A2(n10557), .B1(
        i_data_bus[798]), .B2(n10558), .ZN(n9380) );
  AOI22D1BWP30P140LVT U13796 ( .A1(i_data_bus[894]), .A2(n10559), .B1(
        i_data_bus[830]), .B2(n10560), .ZN(n9379) );
  ND2D1BWP30P140LVT U13797 ( .A1(n9380), .A2(n9379), .ZN(N5645) );
  AOI22D1BWP30P140LVT U13798 ( .A1(i_data_bus[863]), .A2(n10557), .B1(
        i_data_bus[799]), .B2(n10558), .ZN(n9382) );
  AOI22D1BWP30P140LVT U13799 ( .A1(i_data_bus[895]), .A2(n10559), .B1(
        i_data_bus[831]), .B2(n10560), .ZN(n9381) );
  ND2D1BWP30P140LVT U13800 ( .A1(n9382), .A2(n9381), .ZN(N5646) );
  AOI22D1BWP30P140LVT U13801 ( .A1(i_data_bus[863]), .A2(n10590), .B1(
        i_data_bus[799]), .B2(n10589), .ZN(n9384) );
  AOI22D1BWP30P140LVT U13802 ( .A1(i_data_bus[895]), .A2(n10591), .B1(
        i_data_bus[831]), .B2(n10592), .ZN(n9383) );
  ND2D1BWP30P140LVT U13803 ( .A1(n9384), .A2(n9383), .ZN(N3772) );
  AOI22D1BWP30P140LVT U13804 ( .A1(i_data_bus[794]), .A2(n10589), .B1(
        i_data_bus[890]), .B2(n10591), .ZN(n9386) );
  AOI22D1BWP30P140LVT U13805 ( .A1(i_data_bus[858]), .A2(n10590), .B1(
        i_data_bus[826]), .B2(n10592), .ZN(n9385) );
  ND2D1BWP30P140LVT U13806 ( .A1(n9386), .A2(n9385), .ZN(N3767) );
  AOI22D1BWP30P140LVT U13807 ( .A1(i_data_bus[789]), .A2(n10493), .B1(
        i_data_bus[853]), .B2(n10495), .ZN(n9388) );
  AOI22D1BWP30P140LVT U13808 ( .A1(i_data_bus[885]), .A2(n10494), .B1(
        i_data_bus[821]), .B2(n10496), .ZN(n9387) );
  ND2D1BWP30P140LVT U13809 ( .A1(n9388), .A2(n9387), .ZN(N9384) );
  AOI22D1BWP30P140LVT U13810 ( .A1(i_data_bus[789]), .A2(n10589), .B1(
        i_data_bus[853]), .B2(n10590), .ZN(n9390) );
  AOI22D1BWP30P140LVT U13811 ( .A1(i_data_bus[885]), .A2(n10591), .B1(
        i_data_bus[821]), .B2(n10592), .ZN(n9389) );
  ND2D1BWP30P140LVT U13812 ( .A1(n9390), .A2(n9389), .ZN(N3762) );
  AOI22D1BWP30P140LVT U13813 ( .A1(i_data_bus[768]), .A2(n10493), .B1(
        i_data_bus[864]), .B2(n10494), .ZN(n9392) );
  AOI22D1BWP30P140LVT U13814 ( .A1(i_data_bus[832]), .A2(n10495), .B1(
        i_data_bus[800]), .B2(n10496), .ZN(n9391) );
  ND2D1BWP30P140LVT U13815 ( .A1(n9392), .A2(n9391), .ZN(N9363) );
  AOI22D1BWP30P140LVT U13816 ( .A1(i_data_bus[840]), .A2(n10557), .B1(
        i_data_bus[776]), .B2(n10558), .ZN(n9394) );
  AOI22D1BWP30P140LVT U13817 ( .A1(i_data_bus[872]), .A2(n10559), .B1(
        i_data_bus[808]), .B2(n10560), .ZN(n9393) );
  ND2D1BWP30P140LVT U13818 ( .A1(n9394), .A2(n9393), .ZN(N5623) );
  AOI22D1BWP30P140LVT U13819 ( .A1(i_data_bus[879]), .A2(n10591), .B1(
        i_data_bus[847]), .B2(n10590), .ZN(n9396) );
  AOI22D1BWP30P140LVT U13820 ( .A1(i_data_bus[783]), .A2(n10589), .B1(
        i_data_bus[815]), .B2(n10592), .ZN(n9395) );
  ND2D1BWP30P140LVT U13821 ( .A1(n9396), .A2(n9395), .ZN(N3756) );
  AOI22D1BWP30P140LVT U13822 ( .A1(i_data_bus[866]), .A2(n10494), .B1(
        i_data_bus[770]), .B2(n10493), .ZN(n9398) );
  AOI22D1BWP30P140LVT U13823 ( .A1(i_data_bus[834]), .A2(n10495), .B1(
        i_data_bus[802]), .B2(n10496), .ZN(n9397) );
  ND2D1BWP30P140LVT U13824 ( .A1(n9398), .A2(n9397), .ZN(N9365) );
  AOI22D1BWP30P140LVT U13825 ( .A1(i_data_bus[797]), .A2(n10493), .B1(
        i_data_bus[861]), .B2(n10495), .ZN(n9400) );
  AOI22D1BWP30P140LVT U13826 ( .A1(i_data_bus[893]), .A2(n10494), .B1(
        i_data_bus[829]), .B2(n10496), .ZN(n9399) );
  ND2D1BWP30P140LVT U13827 ( .A1(n9400), .A2(n9399), .ZN(N9392) );
  AOI22D1BWP30P140LVT U13828 ( .A1(i_data_bus[867]), .A2(n10591), .B1(
        i_data_bus[835]), .B2(n10590), .ZN(n9402) );
  AOI22D1BWP30P140LVT U13829 ( .A1(i_data_bus[771]), .A2(n10589), .B1(
        i_data_bus[803]), .B2(n10592), .ZN(n9401) );
  ND2D1BWP30P140LVT U13830 ( .A1(n9402), .A2(n9401), .ZN(N3744) );
  AOI22D1BWP30P140LVT U13831 ( .A1(i_data_bus[858]), .A2(n10495), .B1(
        i_data_bus[890]), .B2(n10494), .ZN(n9404) );
  AOI22D1BWP30P140LVT U13832 ( .A1(i_data_bus[794]), .A2(n10493), .B1(
        i_data_bus[826]), .B2(n10496), .ZN(n9403) );
  ND2D1BWP30P140LVT U13833 ( .A1(n9404), .A2(n9403), .ZN(N9389) );
  AOI22D1BWP30P140LVT U13834 ( .A1(i_data_bus[888]), .A2(n10494), .B1(
        i_data_bus[792]), .B2(n10493), .ZN(n9406) );
  AOI22D1BWP30P140LVT U13835 ( .A1(i_data_bus[856]), .A2(n10495), .B1(
        i_data_bus[824]), .B2(n10496), .ZN(n9405) );
  ND2D1BWP30P140LVT U13836 ( .A1(n9406), .A2(n9405), .ZN(N9387) );
  AOI22D1BWP30P140LVT U13837 ( .A1(i_data_bus[994]), .A2(n10489), .B1(
        i_data_bus[930]), .B2(n10491), .ZN(n9408) );
  AOI22D1BWP30P140LVT U13838 ( .A1(i_data_bus[898]), .A2(n10492), .B1(
        i_data_bus[962]), .B2(n10490), .ZN(n9407) );
  ND2D1BWP30P140LVT U13839 ( .A1(n9408), .A2(n9407), .ZN(N9581) );
  AOI22D1BWP30P140LVT U13840 ( .A1(i_data_bus[941]), .A2(n10491), .B1(
        i_data_bus[909]), .B2(n10492), .ZN(n9410) );
  AOI22D1BWP30P140LVT U13841 ( .A1(i_data_bus[1005]), .A2(n10489), .B1(
        i_data_bus[973]), .B2(n10490), .ZN(n9409) );
  ND2D1BWP30P140LVT U13842 ( .A1(n9410), .A2(n9409), .ZN(N9592) );
  AOI22D1BWP30P140LVT U13843 ( .A1(i_data_bus[1014]), .A2(n10489), .B1(
        i_data_bus[918]), .B2(n10492), .ZN(n9412) );
  AOI22D1BWP30P140LVT U13844 ( .A1(i_data_bus[950]), .A2(n10491), .B1(
        i_data_bus[982]), .B2(n10490), .ZN(n9411) );
  ND2D1BWP30P140LVT U13845 ( .A1(n9412), .A2(n9411), .ZN(N9601) );
  AOI22D1BWP30P140LVT U13846 ( .A1(i_data_bus[912]), .A2(n10492), .B1(
        i_data_bus[944]), .B2(n10491), .ZN(n9414) );
  AOI22D1BWP30P140LVT U13847 ( .A1(i_data_bus[1008]), .A2(n10489), .B1(
        i_data_bus[976]), .B2(n10490), .ZN(n9413) );
  ND2D1BWP30P140LVT U13848 ( .A1(n9414), .A2(n9413), .ZN(N9595) );
  AOI22D1BWP30P140LVT U13849 ( .A1(i_data_bus[1009]), .A2(n10489), .B1(
        i_data_bus[945]), .B2(n10491), .ZN(n9416) );
  AOI22D1BWP30P140LVT U13850 ( .A1(i_data_bus[913]), .A2(n10492), .B1(
        i_data_bus[977]), .B2(n10490), .ZN(n9415) );
  ND2D1BWP30P140LVT U13851 ( .A1(n9416), .A2(n9415), .ZN(N9596) );
  AOI22D1BWP30P140LVT U13852 ( .A1(i_data_bus[1018]), .A2(n10489), .B1(
        i_data_bus[922]), .B2(n10492), .ZN(n9418) );
  AOI22D1BWP30P140LVT U13853 ( .A1(i_data_bus[954]), .A2(n10491), .B1(
        i_data_bus[986]), .B2(n10490), .ZN(n9417) );
  ND2D1BWP30P140LVT U13854 ( .A1(n9418), .A2(n9417), .ZN(N9605) );
  AOI22D1BWP30P140LVT U13855 ( .A1(i_data_bus[943]), .A2(n10491), .B1(
        i_data_bus[911]), .B2(n10492), .ZN(n9420) );
  AOI22D1BWP30P140LVT U13856 ( .A1(i_data_bus[1007]), .A2(n10489), .B1(
        i_data_bus[975]), .B2(n10490), .ZN(n9419) );
  ND2D1BWP30P140LVT U13857 ( .A1(n9420), .A2(n9419), .ZN(N9594) );
  AOI22D1BWP30P140LVT U13858 ( .A1(i_data_bus[903]), .A2(n10492), .B1(
        i_data_bus[999]), .B2(n10489), .ZN(n9422) );
  AOI22D1BWP30P140LVT U13859 ( .A1(i_data_bus[935]), .A2(n10491), .B1(
        i_data_bus[967]), .B2(n10490), .ZN(n9421) );
  ND2D1BWP30P140LVT U13860 ( .A1(n9422), .A2(n9421), .ZN(N9586) );
  AOI22D1BWP30P140LVT U13861 ( .A1(i_data_bus[32]), .A2(n10453), .B1(
        i_data_bus[64]), .B2(n10454), .ZN(n9424) );
  AOI22D1BWP30P140LVT U13862 ( .A1(i_data_bus[96]), .A2(n10455), .B1(
        i_data_bus[0]), .B2(n10456), .ZN(n9423) );
  ND2D1BWP30P140LVT U13863 ( .A1(n9424), .A2(n9423), .ZN(N11815) );
  AOI22D1BWP30P140LVT U13864 ( .A1(i_data_bus[51]), .A2(n10453), .B1(
        i_data_bus[83]), .B2(n10454), .ZN(n9426) );
  AOI22D1BWP30P140LVT U13865 ( .A1(i_data_bus[115]), .A2(n10455), .B1(
        i_data_bus[19]), .B2(n10456), .ZN(n9425) );
  ND2D1BWP30P140LVT U13866 ( .A1(n9426), .A2(n9425), .ZN(N11834) );
  AOI22D1BWP30P140LVT U13867 ( .A1(i_data_bus[61]), .A2(n10453), .B1(
        i_data_bus[125]), .B2(n10455), .ZN(n9428) );
  AOI22D1BWP30P140LVT U13868 ( .A1(i_data_bus[93]), .A2(n10454), .B1(
        i_data_bus[29]), .B2(n10456), .ZN(n9427) );
  ND2D1BWP30P140LVT U13869 ( .A1(n9428), .A2(n9427), .ZN(N11844) );
  AOI22D1BWP30P140LVT U13870 ( .A1(i_data_bus[89]), .A2(n10454), .B1(
        i_data_bus[57]), .B2(n10453), .ZN(n9430) );
  AOI22D1BWP30P140LVT U13871 ( .A1(i_data_bus[121]), .A2(n10455), .B1(
        i_data_bus[25]), .B2(n10456), .ZN(n9429) );
  ND2D1BWP30P140LVT U13872 ( .A1(n9430), .A2(n9429), .ZN(N11840) );
  AOI22D1BWP30P140LVT U13873 ( .A1(i_data_bus[90]), .A2(n10454), .B1(
        i_data_bus[122]), .B2(n10455), .ZN(n9432) );
  AOI22D1BWP30P140LVT U13874 ( .A1(i_data_bus[58]), .A2(n10453), .B1(
        i_data_bus[26]), .B2(n10456), .ZN(n9431) );
  ND2D1BWP30P140LVT U13875 ( .A1(n9432), .A2(n9431), .ZN(N11841) );
  AOI22D1BWP30P140LVT U13876 ( .A1(i_data_bus[98]), .A2(n10455), .B1(
        i_data_bus[34]), .B2(n10453), .ZN(n9434) );
  AOI22D1BWP30P140LVT U13877 ( .A1(i_data_bus[66]), .A2(n10454), .B1(
        i_data_bus[2]), .B2(n10456), .ZN(n9433) );
  ND2D1BWP30P140LVT U13878 ( .A1(n9434), .A2(n9433), .ZN(N11817) );
  AOI22D1BWP30P140LVT U13879 ( .A1(i_data_bus[104]), .A2(n10455), .B1(
        i_data_bus[72]), .B2(n10454), .ZN(n9436) );
  AOI22D1BWP30P140LVT U13880 ( .A1(i_data_bus[40]), .A2(n10453), .B1(
        i_data_bus[8]), .B2(n10456), .ZN(n9435) );
  ND2D1BWP30P140LVT U13881 ( .A1(n9436), .A2(n9435), .ZN(N11823) );
  AOI22D1BWP30P140LVT U13882 ( .A1(i_data_bus[53]), .A2(n10453), .B1(
        i_data_bus[85]), .B2(n10454), .ZN(n9438) );
  AOI22D1BWP30P140LVT U13883 ( .A1(i_data_bus[117]), .A2(n10455), .B1(
        i_data_bus[21]), .B2(n10456), .ZN(n9437) );
  ND2D1BWP30P140LVT U13884 ( .A1(n9438), .A2(n9437), .ZN(N11836) );
  AOI22D1BWP30P140LVT U13885 ( .A1(i_data_bus[67]), .A2(n10454), .B1(
        i_data_bus[99]), .B2(n10455), .ZN(n9440) );
  AOI22D1BWP30P140LVT U13886 ( .A1(i_data_bus[35]), .A2(n10453), .B1(
        i_data_bus[3]), .B2(n10456), .ZN(n9439) );
  ND2D1BWP30P140LVT U13887 ( .A1(n9440), .A2(n9439), .ZN(N11818) );
  AOI22D1BWP30P140LVT U13888 ( .A1(i_data_bus[48]), .A2(n10453), .B1(
        i_data_bus[80]), .B2(n10454), .ZN(n9442) );
  AOI22D1BWP30P140LVT U13889 ( .A1(i_data_bus[112]), .A2(n10455), .B1(
        i_data_bus[16]), .B2(n10456), .ZN(n9441) );
  ND2D1BWP30P140LVT U13890 ( .A1(n9442), .A2(n9441), .ZN(N11831) );
  AOI22D1BWP30P140LVT U13891 ( .A1(i_data_bus[60]), .A2(n10453), .B1(
        i_data_bus[92]), .B2(n10454), .ZN(n9444) );
  AOI22D1BWP30P140LVT U13892 ( .A1(i_data_bus[124]), .A2(n10455), .B1(
        i_data_bus[28]), .B2(n10456), .ZN(n9443) );
  ND2D1BWP30P140LVT U13893 ( .A1(n9444), .A2(n9443), .ZN(N11843) );
  AOI22D1BWP30P140LVT U13894 ( .A1(i_data_bus[94]), .A2(n10454), .B1(
        i_data_bus[62]), .B2(n10453), .ZN(n9446) );
  AOI22D1BWP30P140LVT U13895 ( .A1(i_data_bus[126]), .A2(n10455), .B1(
        i_data_bus[30]), .B2(n10456), .ZN(n9445) );
  ND2D1BWP30P140LVT U13896 ( .A1(n9446), .A2(n9445), .ZN(N11845) );
  AOI22D1BWP30P140LVT U13897 ( .A1(i_data_bus[76]), .A2(n10454), .B1(
        i_data_bus[108]), .B2(n10455), .ZN(n9448) );
  AOI22D1BWP30P140LVT U13898 ( .A1(i_data_bus[44]), .A2(n10453), .B1(
        i_data_bus[12]), .B2(n10456), .ZN(n9447) );
  ND2D1BWP30P140LVT U13899 ( .A1(n9448), .A2(n9447), .ZN(N11827) );
  AOI22D1BWP30P140LVT U13900 ( .A1(i_data_bus[222]), .A2(n10419), .B1(
        i_data_bus[254]), .B2(n10418), .ZN(n9450) );
  AOI22D1BWP30P140LVT U13901 ( .A1(i_data_bus[190]), .A2(n10420), .B1(
        i_data_bus[158]), .B2(n10417), .ZN(n9449) );
  ND2D1BWP30P140LVT U13902 ( .A1(n9450), .A2(n9449), .ZN(N13935) );
  AOI22D1BWP30P140LVT U13903 ( .A1(i_data_bus[193]), .A2(n10419), .B1(
        i_data_bus[225]), .B2(n10418), .ZN(n9452) );
  AOI22D1BWP30P140LVT U13904 ( .A1(i_data_bus[161]), .A2(n10420), .B1(
        i_data_bus[129]), .B2(n10417), .ZN(n9451) );
  ND2D1BWP30P140LVT U13905 ( .A1(n9452), .A2(n9451), .ZN(N13906) );
  AOI22D1BWP30P140LVT U13906 ( .A1(i_data_bus[177]), .A2(n10420), .B1(
        i_data_bus[241]), .B2(n10418), .ZN(n9454) );
  AOI22D1BWP30P140LVT U13907 ( .A1(i_data_bus[209]), .A2(n10419), .B1(
        i_data_bus[145]), .B2(n10417), .ZN(n9453) );
  ND2D1BWP30P140LVT U13908 ( .A1(n9454), .A2(n9453), .ZN(N13922) );
  AOI22D1BWP30P140LVT U13909 ( .A1(i_data_bus[255]), .A2(n10418), .B1(
        i_data_bus[191]), .B2(n10420), .ZN(n9456) );
  AOI22D1BWP30P140LVT U13910 ( .A1(i_data_bus[223]), .A2(n10419), .B1(
        i_data_bus[159]), .B2(n10417), .ZN(n9455) );
  ND2D1BWP30P140LVT U13911 ( .A1(n9456), .A2(n9455), .ZN(N13936) );
  AOI22D1BWP30P140LVT U13912 ( .A1(i_data_bus[170]), .A2(n10420), .B1(
        i_data_bus[202]), .B2(n10419), .ZN(n9458) );
  AOI22D1BWP30P140LVT U13913 ( .A1(i_data_bus[234]), .A2(n10418), .B1(
        i_data_bus[138]), .B2(n10417), .ZN(n9457) );
  ND2D1BWP30P140LVT U13914 ( .A1(n9458), .A2(n9457), .ZN(N13915) );
  AOI22D1BWP30P140LVT U13915 ( .A1(i_data_bus[168]), .A2(n10420), .B1(
        i_data_bus[232]), .B2(n10418), .ZN(n9460) );
  AOI22D1BWP30P140LVT U13916 ( .A1(i_data_bus[200]), .A2(n10419), .B1(
        i_data_bus[136]), .B2(n10417), .ZN(n9459) );
  ND2D1BWP30P140LVT U13917 ( .A1(n9460), .A2(n9459), .ZN(N13913) );
  AOI22D1BWP30P140LVT U13918 ( .A1(i_data_bus[235]), .A2(n10418), .B1(
        i_data_bus[171]), .B2(n10420), .ZN(n9462) );
  AOI22D1BWP30P140LVT U13919 ( .A1(i_data_bus[203]), .A2(n10419), .B1(
        i_data_bus[139]), .B2(n10417), .ZN(n9461) );
  ND2D1BWP30P140LVT U13920 ( .A1(n9462), .A2(n9461), .ZN(N13916) );
  AOI22D1BWP30P140LVT U13921 ( .A1(i_data_bus[231]), .A2(n10418), .B1(
        i_data_bus[167]), .B2(n10420), .ZN(n9464) );
  AOI22D1BWP30P140LVT U13922 ( .A1(i_data_bus[199]), .A2(n10419), .B1(
        i_data_bus[135]), .B2(n10417), .ZN(n9463) );
  ND2D1BWP30P140LVT U13923 ( .A1(n9464), .A2(n9463), .ZN(N13912) );
  AOI22D1BWP30P140LVT U13924 ( .A1(i_data_bus[211]), .A2(n10419), .B1(
        i_data_bus[243]), .B2(n10418), .ZN(n9466) );
  AOI22D1BWP30P140LVT U13925 ( .A1(i_data_bus[179]), .A2(n10420), .B1(
        i_data_bus[147]), .B2(n10417), .ZN(n9465) );
  ND2D1BWP30P140LVT U13926 ( .A1(n9466), .A2(n9465), .ZN(N13924) );
  AOI22D1BWP30P140LVT U13927 ( .A1(i_data_bus[162]), .A2(n10420), .B1(
        i_data_bus[226]), .B2(n10418), .ZN(n9468) );
  AOI22D1BWP30P140LVT U13928 ( .A1(i_data_bus[194]), .A2(n10419), .B1(
        i_data_bus[130]), .B2(n10417), .ZN(n9467) );
  ND2D1BWP30P140LVT U13929 ( .A1(n9468), .A2(n9467), .ZN(N13907) );
  AOI22D1BWP30P140LVT U13930 ( .A1(i_data_bus[932]), .A2(n10521), .B1(
        i_data_bus[900]), .B2(n10524), .ZN(n9470) );
  AOI22D1BWP30P140LVT U13931 ( .A1(i_data_bus[996]), .A2(n10523), .B1(
        i_data_bus[964]), .B2(n10522), .ZN(n9469) );
  ND2D1BWP30P140LVT U13932 ( .A1(n9470), .A2(n9469), .ZN(N7709) );
  AOI22D1BWP30P140LVT U13933 ( .A1(i_data_bus[951]), .A2(n10521), .B1(
        i_data_bus[1015]), .B2(n10523), .ZN(n9472) );
  AOI22D1BWP30P140LVT U13934 ( .A1(i_data_bus[919]), .A2(n10524), .B1(
        i_data_bus[983]), .B2(n10522), .ZN(n9471) );
  ND2D1BWP30P140LVT U13935 ( .A1(n9472), .A2(n9471), .ZN(N7728) );
  AOI22D1BWP30P140LVT U13936 ( .A1(i_data_bus[935]), .A2(n10521), .B1(
        i_data_bus[999]), .B2(n10523), .ZN(n9474) );
  AOI22D1BWP30P140LVT U13937 ( .A1(i_data_bus[903]), .A2(n10524), .B1(
        i_data_bus[967]), .B2(n10522), .ZN(n9473) );
  ND2D1BWP30P140LVT U13938 ( .A1(n9474), .A2(n9473), .ZN(N7712) );
  AOI22D1BWP30P140LVT U13939 ( .A1(i_data_bus[1023]), .A2(n10523), .B1(
        i_data_bus[959]), .B2(n10521), .ZN(n9476) );
  AOI22D1BWP30P140LVT U13940 ( .A1(i_data_bus[927]), .A2(n10524), .B1(
        i_data_bus[991]), .B2(n10522), .ZN(n9475) );
  ND2D1BWP30P140LVT U13941 ( .A1(n9476), .A2(n9475), .ZN(N7736) );
  AOI22D1BWP30P140LVT U13942 ( .A1(i_data_bus[929]), .A2(n10521), .B1(
        i_data_bus[897]), .B2(n10524), .ZN(n9478) );
  AOI22D1BWP30P140LVT U13943 ( .A1(i_data_bus[993]), .A2(n10523), .B1(
        i_data_bus[961]), .B2(n10522), .ZN(n9477) );
  ND2D1BWP30P140LVT U13944 ( .A1(n9478), .A2(n9477), .ZN(N7706) );
  AOI22D1BWP30P140LVT U13945 ( .A1(i_data_bus[941]), .A2(n10521), .B1(
        i_data_bus[909]), .B2(n10524), .ZN(n9480) );
  AOI22D1BWP30P140LVT U13946 ( .A1(i_data_bus[1005]), .A2(n10523), .B1(
        i_data_bus[973]), .B2(n10522), .ZN(n9479) );
  ND2D1BWP30P140LVT U13947 ( .A1(n9480), .A2(n9479), .ZN(N7718) );
  AOI22D1BWP30P140LVT U13948 ( .A1(i_data_bus[910]), .A2(n10524), .B1(
        i_data_bus[942]), .B2(n10521), .ZN(n9482) );
  AOI22D1BWP30P140LVT U13949 ( .A1(i_data_bus[1006]), .A2(n10523), .B1(
        i_data_bus[974]), .B2(n10522), .ZN(n9481) );
  ND2D1BWP30P140LVT U13950 ( .A1(n9482), .A2(n9481), .ZN(N7719) );
  AOI22D1BWP30P140LVT U13951 ( .A1(i_data_bus[939]), .A2(n10521), .B1(
        i_data_bus[907]), .B2(n10524), .ZN(n9484) );
  AOI22D1BWP30P140LVT U13952 ( .A1(i_data_bus[1003]), .A2(n10523), .B1(
        i_data_bus[971]), .B2(n10522), .ZN(n9483) );
  ND2D1BWP30P140LVT U13953 ( .A1(n9484), .A2(n9483), .ZN(N7716) );
  AOI22D1BWP30P140LVT U13954 ( .A1(i_data_bus[1008]), .A2(n10523), .B1(
        i_data_bus[944]), .B2(n10521), .ZN(n9486) );
  AOI22D1BWP30P140LVT U13955 ( .A1(i_data_bus[912]), .A2(n10524), .B1(
        i_data_bus[976]), .B2(n10522), .ZN(n9485) );
  ND2D1BWP30P140LVT U13956 ( .A1(n9486), .A2(n9485), .ZN(N7721) );
  AOI22D1BWP30P140LVT U13957 ( .A1(i_data_bus[1007]), .A2(n10523), .B1(
        i_data_bus[911]), .B2(n10524), .ZN(n9488) );
  AOI22D1BWP30P140LVT U13958 ( .A1(i_data_bus[943]), .A2(n10521), .B1(
        i_data_bus[975]), .B2(n10522), .ZN(n9487) );
  ND2D1BWP30P140LVT U13959 ( .A1(n9488), .A2(n9487), .ZN(N7720) );
  AOI22D1BWP30P140LVT U13960 ( .A1(i_data_bus[533]), .A2(n10533), .B1(
        i_data_bus[565]), .B2(n10535), .ZN(n9490) );
  AOI22D1BWP30P140LVT U13961 ( .A1(i_data_bus[597]), .A2(n10536), .B1(
        i_data_bus[629]), .B2(n10534), .ZN(n9489) );
  ND2D1BWP30P140LVT U13962 ( .A1(n9490), .A2(n9489), .ZN(N7078) );
  AOI22D1BWP30P140LVT U13963 ( .A1(i_data_bus[558]), .A2(n10472), .B1(
        i_data_bus[526]), .B2(n10471), .ZN(n9492) );
  AOI22D1BWP30P140LVT U13964 ( .A1(i_data_bus[590]), .A2(n10469), .B1(
        i_data_bus[622]), .B2(n10470), .ZN(n9491) );
  ND2D1BWP30P140LVT U13965 ( .A1(n9492), .A2(n9491), .ZN(N10819) );
  AOI22D1BWP30P140LVT U13966 ( .A1(i_data_bus[592]), .A2(n10536), .B1(
        i_data_bus[528]), .B2(n10533), .ZN(n9494) );
  AOI22D1BWP30P140LVT U13967 ( .A1(i_data_bus[560]), .A2(n10535), .B1(
        i_data_bus[624]), .B2(n10534), .ZN(n9493) );
  ND2D1BWP30P140LVT U13968 ( .A1(n9494), .A2(n9493), .ZN(N7073) );
  AOI22D1BWP30P140LVT U13969 ( .A1(i_data_bus[554]), .A2(n10472), .B1(
        i_data_bus[522]), .B2(n10471), .ZN(n9496) );
  AOI22D1BWP30P140LVT U13970 ( .A1(i_data_bus[586]), .A2(n10469), .B1(
        i_data_bus[618]), .B2(n10470), .ZN(n9495) );
  ND2D1BWP30P140LVT U13971 ( .A1(n9496), .A2(n9495), .ZN(N10815) );
  AOI22D1BWP30P140LVT U13972 ( .A1(i_data_bus[556]), .A2(n10535), .B1(
        i_data_bus[588]), .B2(n10536), .ZN(n9498) );
  AOI22D1BWP30P140LVT U13973 ( .A1(i_data_bus[524]), .A2(n10533), .B1(
        i_data_bus[620]), .B2(n10534), .ZN(n9497) );
  ND2D1BWP30P140LVT U13974 ( .A1(n9498), .A2(n9497), .ZN(N7069) );
  AOI22D1BWP30P140LVT U13975 ( .A1(i_data_bus[553]), .A2(n10535), .B1(
        i_data_bus[585]), .B2(n10536), .ZN(n9500) );
  AOI22D1BWP30P140LVT U13976 ( .A1(i_data_bus[521]), .A2(n10533), .B1(
        i_data_bus[617]), .B2(n10534), .ZN(n9499) );
  ND2D1BWP30P140LVT U13977 ( .A1(n9500), .A2(n9499), .ZN(N7066) );
  AOI22D1BWP30P140LVT U13978 ( .A1(i_data_bus[596]), .A2(n10469), .B1(
        i_data_bus[532]), .B2(n10471), .ZN(n9502) );
  AOI22D1BWP30P140LVT U13979 ( .A1(i_data_bus[564]), .A2(n10472), .B1(
        i_data_bus[628]), .B2(n10470), .ZN(n9501) );
  ND2D1BWP30P140LVT U13980 ( .A1(n9502), .A2(n9501), .ZN(N10825) );
  AOI22D1BWP30P140LVT U13981 ( .A1(i_data_bus[601]), .A2(n10536), .B1(
        i_data_bus[569]), .B2(n10535), .ZN(n9504) );
  AOI22D1BWP30P140LVT U13982 ( .A1(i_data_bus[537]), .A2(n10533), .B1(
        i_data_bus[633]), .B2(n10534), .ZN(n9503) );
  ND2D1BWP30P140LVT U13983 ( .A1(n9504), .A2(n9503), .ZN(N7082) );
  AOI22D1BWP30P140LVT U13984 ( .A1(i_data_bus[586]), .A2(n10536), .B1(
        i_data_bus[522]), .B2(n10533), .ZN(n9506) );
  AOI22D1BWP30P140LVT U13985 ( .A1(i_data_bus[554]), .A2(n10535), .B1(
        i_data_bus[618]), .B2(n10534), .ZN(n9505) );
  ND2D1BWP30P140LVT U13986 ( .A1(n9506), .A2(n9505), .ZN(N7067) );
  AOI22D1BWP30P140LVT U13987 ( .A1(i_data_bus[548]), .A2(n10472), .B1(
        i_data_bus[580]), .B2(n10469), .ZN(n9508) );
  AOI22D1BWP30P140LVT U13988 ( .A1(i_data_bus[516]), .A2(n10471), .B1(
        i_data_bus[612]), .B2(n10470), .ZN(n9507) );
  ND2D1BWP30P140LVT U13989 ( .A1(n9508), .A2(n9507), .ZN(N10809) );
  AOI22D1BWP30P140LVT U13990 ( .A1(i_data_bus[556]), .A2(n10472), .B1(
        i_data_bus[524]), .B2(n10471), .ZN(n9510) );
  AOI22D1BWP30P140LVT U13991 ( .A1(i_data_bus[588]), .A2(n10469), .B1(
        i_data_bus[620]), .B2(n10470), .ZN(n9509) );
  ND2D1BWP30P140LVT U13992 ( .A1(n9510), .A2(n9509), .ZN(N10817) );
  AOI22D1BWP30P140LVT U13993 ( .A1(i_data_bus[598]), .A2(n10469), .B1(
        i_data_bus[534]), .B2(n10471), .ZN(n9512) );
  AOI22D1BWP30P140LVT U13994 ( .A1(i_data_bus[566]), .A2(n10472), .B1(
        i_data_bus[630]), .B2(n10470), .ZN(n9511) );
  ND2D1BWP30P140LVT U13995 ( .A1(n9512), .A2(n9511), .ZN(N10827) );
  AOI22D1BWP30P140LVT U13996 ( .A1(i_data_bus[600]), .A2(n10536), .B1(
        i_data_bus[568]), .B2(n10535), .ZN(n9514) );
  AOI22D1BWP30P140LVT U13997 ( .A1(i_data_bus[536]), .A2(n10533), .B1(
        i_data_bus[632]), .B2(n10534), .ZN(n9513) );
  ND2D1BWP30P140LVT U13998 ( .A1(n9514), .A2(n9513), .ZN(N7081) );
  AOI22D1BWP30P140LVT U13999 ( .A1(i_data_bus[559]), .A2(n10472), .B1(
        i_data_bus[527]), .B2(n10471), .ZN(n9516) );
  AOI22D1BWP30P140LVT U14000 ( .A1(i_data_bus[591]), .A2(n10469), .B1(
        i_data_bus[623]), .B2(n10470), .ZN(n9515) );
  ND2D1BWP30P140LVT U14001 ( .A1(n9516), .A2(n9515), .ZN(N10820) );
  AOI22D1BWP30P140LVT U14002 ( .A1(i_data_bus[572]), .A2(n10535), .B1(
        i_data_bus[540]), .B2(n10533), .ZN(n9518) );
  AOI22D1BWP30P140LVT U14003 ( .A1(i_data_bus[604]), .A2(n10536), .B1(
        i_data_bus[636]), .B2(n10534), .ZN(n9517) );
  ND2D1BWP30P140LVT U14004 ( .A1(n9518), .A2(n9517), .ZN(N7085) );
  AOI22D1BWP30P140LVT U14005 ( .A1(i_data_bus[539]), .A2(n10471), .B1(
        i_data_bus[603]), .B2(n10469), .ZN(n9520) );
  AOI22D1BWP30P140LVT U14006 ( .A1(i_data_bus[571]), .A2(n10472), .B1(
        i_data_bus[635]), .B2(n10470), .ZN(n9519) );
  ND2D1BWP30P140LVT U14007 ( .A1(n9520), .A2(n9519), .ZN(N10832) );
  AOI22D1BWP30P140LVT U14008 ( .A1(i_data_bus[530]), .A2(n10471), .B1(
        i_data_bus[562]), .B2(n10472), .ZN(n9522) );
  AOI22D1BWP30P140LVT U14009 ( .A1(i_data_bus[594]), .A2(n10469), .B1(
        i_data_bus[626]), .B2(n10470), .ZN(n9521) );
  ND2D1BWP30P140LVT U14010 ( .A1(n9522), .A2(n9521), .ZN(N10823) );
  AOI22D1BWP30P140LVT U14011 ( .A1(i_data_bus[551]), .A2(n10535), .B1(
        i_data_bus[583]), .B2(n10536), .ZN(n9524) );
  AOI22D1BWP30P140LVT U14012 ( .A1(i_data_bus[519]), .A2(n10533), .B1(
        i_data_bus[615]), .B2(n10534), .ZN(n9523) );
  ND2D1BWP30P140LVT U14013 ( .A1(n9524), .A2(n9523), .ZN(N7064) );
  AOI22D1BWP30P140LVT U14014 ( .A1(i_data_bus[587]), .A2(n10469), .B1(
        i_data_bus[555]), .B2(n10472), .ZN(n9526) );
  AOI22D1BWP30P140LVT U14015 ( .A1(i_data_bus[523]), .A2(n10471), .B1(
        i_data_bus[619]), .B2(n10470), .ZN(n9525) );
  ND2D1BWP30P140LVT U14016 ( .A1(n9526), .A2(n9525), .ZN(N10816) );
  AOI22D1BWP30P140LVT U14017 ( .A1(i_data_bus[543]), .A2(n10533), .B1(
        i_data_bus[575]), .B2(n10535), .ZN(n9528) );
  AOI22D1BWP30P140LVT U14018 ( .A1(i_data_bus[607]), .A2(n10536), .B1(
        i_data_bus[639]), .B2(n10534), .ZN(n9527) );
  ND2D1BWP30P140LVT U14019 ( .A1(n9528), .A2(n9527), .ZN(N7088) );
  AOI22D1BWP30P140LVT U14020 ( .A1(i_data_bus[543]), .A2(n10471), .B1(
        i_data_bus[575]), .B2(n10472), .ZN(n9530) );
  AOI22D1BWP30P140LVT U14021 ( .A1(i_data_bus[607]), .A2(n10469), .B1(
        i_data_bus[639]), .B2(n10470), .ZN(n9529) );
  ND2D1BWP30P140LVT U14022 ( .A1(n9530), .A2(n9529), .ZN(N10836) );
  AOI22D1BWP30P140LVT U14023 ( .A1(i_data_bus[106]), .A2(n10549), .B1(
        i_data_bus[42]), .B2(n10550), .ZN(n9532) );
  AOI22D1BWP30P140LVT U14024 ( .A1(i_data_bus[74]), .A2(n10551), .B1(
        i_data_bus[10]), .B2(n10552), .ZN(n9531) );
  ND2D1BWP30P140LVT U14025 ( .A1(n9532), .A2(n9531), .ZN(N6203) );
  AOI22D1BWP30P140LVT U14026 ( .A1(i_data_bus[76]), .A2(n10551), .B1(
        i_data_bus[108]), .B2(n10549), .ZN(n9534) );
  AOI22D1BWP30P140LVT U14027 ( .A1(i_data_bus[44]), .A2(n10550), .B1(
        i_data_bus[12]), .B2(n10552), .ZN(n9533) );
  ND2D1BWP30P140LVT U14028 ( .A1(n9534), .A2(n9533), .ZN(N6205) );
  AOI22D1BWP30P140LVT U14029 ( .A1(i_data_bus[37]), .A2(n10550), .B1(
        i_data_bus[101]), .B2(n10549), .ZN(n9536) );
  AOI22D1BWP30P140LVT U14030 ( .A1(i_data_bus[69]), .A2(n10551), .B1(
        i_data_bus[5]), .B2(n10552), .ZN(n9535) );
  ND2D1BWP30P140LVT U14031 ( .A1(n9536), .A2(n9535), .ZN(N6198) );
  AOI22D1BWP30P140LVT U14032 ( .A1(i_data_bus[118]), .A2(n10549), .B1(
        i_data_bus[54]), .B2(n10550), .ZN(n9538) );
  AOI22D1BWP30P140LVT U14033 ( .A1(i_data_bus[86]), .A2(n10551), .B1(
        i_data_bus[22]), .B2(n10552), .ZN(n9537) );
  ND2D1BWP30P140LVT U14034 ( .A1(n9538), .A2(n9537), .ZN(N6215) );
  AOI22D1BWP30P140LVT U14035 ( .A1(i_data_bus[124]), .A2(n10549), .B1(
        i_data_bus[92]), .B2(n10551), .ZN(n9540) );
  AOI22D1BWP30P140LVT U14036 ( .A1(i_data_bus[60]), .A2(n10550), .B1(
        i_data_bus[28]), .B2(n10552), .ZN(n9539) );
  ND2D1BWP30P140LVT U14037 ( .A1(n9540), .A2(n9539), .ZN(N6221) );
  AOI22D1BWP30P140LVT U14038 ( .A1(i_data_bus[90]), .A2(n10551), .B1(
        i_data_bus[58]), .B2(n10550), .ZN(n9542) );
  AOI22D1BWP30P140LVT U14039 ( .A1(i_data_bus[122]), .A2(n10549), .B1(
        i_data_bus[26]), .B2(n10552), .ZN(n9541) );
  ND2D1BWP30P140LVT U14040 ( .A1(n9542), .A2(n9541), .ZN(N6219) );
  AOI22D1BWP30P140LVT U14041 ( .A1(i_data_bus[48]), .A2(n10550), .B1(
        i_data_bus[112]), .B2(n10549), .ZN(n9544) );
  AOI22D1BWP30P140LVT U14042 ( .A1(i_data_bus[80]), .A2(n10551), .B1(
        i_data_bus[16]), .B2(n10552), .ZN(n9543) );
  ND2D1BWP30P140LVT U14043 ( .A1(n9544), .A2(n9543), .ZN(N6209) );
  AOI22D1BWP30P140LVT U14044 ( .A1(i_data_bus[114]), .A2(n10549), .B1(
        i_data_bus[50]), .B2(n10550), .ZN(n9546) );
  AOI22D1BWP30P140LVT U14045 ( .A1(i_data_bus[82]), .A2(n10551), .B1(
        i_data_bus[18]), .B2(n10552), .ZN(n9545) );
  ND2D1BWP30P140LVT U14046 ( .A1(n9546), .A2(n9545), .ZN(N6211) );
  AOI22D1BWP30P140LVT U14047 ( .A1(i_data_bus[51]), .A2(n10550), .B1(
        i_data_bus[115]), .B2(n10549), .ZN(n9548) );
  AOI22D1BWP30P140LVT U14048 ( .A1(i_data_bus[83]), .A2(n10551), .B1(
        i_data_bus[19]), .B2(n10552), .ZN(n9547) );
  ND2D1BWP30P140LVT U14049 ( .A1(n9548), .A2(n9547), .ZN(N6212) );
  AOI22D1BWP30P140LVT U14050 ( .A1(i_data_bus[35]), .A2(n10550), .B1(
        i_data_bus[99]), .B2(n10549), .ZN(n9550) );
  AOI22D1BWP30P140LVT U14051 ( .A1(i_data_bus[67]), .A2(n10551), .B1(
        i_data_bus[3]), .B2(n10552), .ZN(n9549) );
  ND2D1BWP30P140LVT U14052 ( .A1(n9550), .A2(n9549), .ZN(N6196) );
  AOI22D1BWP30P140LVT U14053 ( .A1(i_data_bus[104]), .A2(n10549), .B1(
        i_data_bus[72]), .B2(n10551), .ZN(n9552) );
  AOI22D1BWP30P140LVT U14054 ( .A1(i_data_bus[40]), .A2(n10550), .B1(
        i_data_bus[8]), .B2(n10552), .ZN(n9551) );
  ND2D1BWP30P140LVT U14055 ( .A1(n9552), .A2(n9551), .ZN(N6201) );
  AOI22D1BWP30P140LVT U14056 ( .A1(i_data_bus[920]), .A2(n10395), .B1(
        i_data_bus[1016]), .B2(n10393), .ZN(n9554) );
  AOI22D1BWP30P140LVT U14057 ( .A1(i_data_bus[952]), .A2(n10394), .B1(
        i_data_bus[984]), .B2(n10396), .ZN(n9553) );
  ND2D1BWP30P140LVT U14058 ( .A1(n9554), .A2(n9553), .ZN(N15225) );
  AOI22D1BWP30P140LVT U14059 ( .A1(i_data_bus[913]), .A2(n10395), .B1(
        i_data_bus[945]), .B2(n10394), .ZN(n9556) );
  AOI22D1BWP30P140LVT U14060 ( .A1(i_data_bus[1009]), .A2(n10393), .B1(
        i_data_bus[977]), .B2(n10396), .ZN(n9555) );
  ND2D1BWP30P140LVT U14061 ( .A1(n9556), .A2(n9555), .ZN(N15218) );
  AOI22D1BWP30P140LVT U14062 ( .A1(i_data_bus[992]), .A2(n10393), .B1(
        i_data_bus[928]), .B2(n10394), .ZN(n9558) );
  AOI22D1BWP30P140LVT U14063 ( .A1(i_data_bus[896]), .A2(n10395), .B1(
        i_data_bus[960]), .B2(n10396), .ZN(n9557) );
  ND2D1BWP30P140LVT U14064 ( .A1(n9558), .A2(n9557), .ZN(N15201) );
  AOI22D1BWP30P140LVT U14065 ( .A1(i_data_bus[910]), .A2(n10395), .B1(
        i_data_bus[942]), .B2(n10394), .ZN(n9560) );
  AOI22D1BWP30P140LVT U14066 ( .A1(i_data_bus[1006]), .A2(n10393), .B1(
        i_data_bus[974]), .B2(n10396), .ZN(n9559) );
  ND2D1BWP30P140LVT U14067 ( .A1(n9560), .A2(n9559), .ZN(N15215) );
  AOI22D1BWP30P140LVT U14068 ( .A1(i_data_bus[923]), .A2(n10395), .B1(
        i_data_bus[1019]), .B2(n10393), .ZN(n9562) );
  AOI22D1BWP30P140LVT U14069 ( .A1(i_data_bus[955]), .A2(n10394), .B1(
        i_data_bus[987]), .B2(n10396), .ZN(n9561) );
  ND2D1BWP30P140LVT U14070 ( .A1(n9562), .A2(n9561), .ZN(N15228) );
  AOI22D1BWP30P140LVT U14071 ( .A1(i_data_bus[934]), .A2(n10394), .B1(
        i_data_bus[902]), .B2(n10395), .ZN(n9564) );
  AOI22D1BWP30P140LVT U14072 ( .A1(i_data_bus[998]), .A2(n10393), .B1(
        i_data_bus[966]), .B2(n10396), .ZN(n9563) );
  ND2D1BWP30P140LVT U14073 ( .A1(n9564), .A2(n9563), .ZN(N15207) );
  AOI22D1BWP30P140LVT U14074 ( .A1(i_data_bus[958]), .A2(n10394), .B1(
        i_data_bus[1022]), .B2(n10393), .ZN(n9566) );
  AOI22D1BWP30P140LVT U14075 ( .A1(i_data_bus[926]), .A2(n10395), .B1(
        i_data_bus[990]), .B2(n10396), .ZN(n9565) );
  ND2D1BWP30P140LVT U14076 ( .A1(n9566), .A2(n9565), .ZN(N15231) );
  AOI22D1BWP30P140LVT U14077 ( .A1(i_data_bus[951]), .A2(n10394), .B1(
        i_data_bus[1015]), .B2(n10393), .ZN(n9568) );
  AOI22D1BWP30P140LVT U14078 ( .A1(i_data_bus[919]), .A2(n10395), .B1(
        i_data_bus[983]), .B2(n10396), .ZN(n9567) );
  ND2D1BWP30P140LVT U14079 ( .A1(n9568), .A2(n9567), .ZN(N15224) );
  AOI22D1BWP30P140LVT U14080 ( .A1(i_data_bus[932]), .A2(n10394), .B1(
        i_data_bus[996]), .B2(n10393), .ZN(n9570) );
  AOI22D1BWP30P140LVT U14081 ( .A1(i_data_bus[900]), .A2(n10395), .B1(
        i_data_bus[964]), .B2(n10396), .ZN(n9569) );
  ND2D1BWP30P140LVT U14082 ( .A1(n9570), .A2(n9569), .ZN(N15205) );
  AOI22D1BWP30P140LVT U14083 ( .A1(i_data_bus[908]), .A2(n10395), .B1(
        i_data_bus[940]), .B2(n10394), .ZN(n9572) );
  AOI22D1BWP30P140LVT U14084 ( .A1(i_data_bus[1004]), .A2(n10393), .B1(
        i_data_bus[972]), .B2(n10396), .ZN(n9571) );
  ND2D1BWP30P140LVT U14085 ( .A1(n9572), .A2(n9571), .ZN(N15213) );
  AOI22D1BWP30P140LVT U14086 ( .A1(i_data_bus[995]), .A2(n10393), .B1(
        i_data_bus[931]), .B2(n10394), .ZN(n9574) );
  AOI22D1BWP30P140LVT U14087 ( .A1(i_data_bus[899]), .A2(n10395), .B1(
        i_data_bus[963]), .B2(n10396), .ZN(n9573) );
  ND2D1BWP30P140LVT U14088 ( .A1(n9574), .A2(n9573), .ZN(N15204) );
  AOI22D1BWP30P140LVT U14089 ( .A1(i_data_bus[1014]), .A2(n10393), .B1(
        i_data_bus[918]), .B2(n10395), .ZN(n9576) );
  AOI22D1BWP30P140LVT U14090 ( .A1(i_data_bus[950]), .A2(n10394), .B1(
        i_data_bus[982]), .B2(n10396), .ZN(n9575) );
  ND2D1BWP30P140LVT U14091 ( .A1(n9576), .A2(n9575), .ZN(N15223) );
  AOI22D1BWP30P140LVT U14092 ( .A1(i_data_bus[601]), .A2(n10565), .B1(
        i_data_bus[569]), .B2(n10567), .ZN(n9578) );
  AOI22D1BWP30P140LVT U14093 ( .A1(i_data_bus[537]), .A2(n10566), .B1(
        i_data_bus[633]), .B2(n10568), .ZN(n9577) );
  ND2D1BWP30P140LVT U14094 ( .A1(n9578), .A2(n9577), .ZN(N5208) );
  AOI22D1BWP30P140LVT U14095 ( .A1(i_data_bus[607]), .A2(n10565), .B1(
        i_data_bus[575]), .B2(n10567), .ZN(n9580) );
  AOI22D1BWP30P140LVT U14096 ( .A1(i_data_bus[543]), .A2(n10566), .B1(
        i_data_bus[639]), .B2(n10568), .ZN(n9579) );
  ND2D1BWP30P140LVT U14097 ( .A1(n9580), .A2(n9579), .ZN(N5214) );
  AOI22D1BWP30P140LVT U14098 ( .A1(i_data_bus[584]), .A2(n10565), .B1(
        i_data_bus[520]), .B2(n10566), .ZN(n9582) );
  AOI22D1BWP30P140LVT U14099 ( .A1(i_data_bus[552]), .A2(n10567), .B1(
        i_data_bus[616]), .B2(n10568), .ZN(n9581) );
  ND2D1BWP30P140LVT U14100 ( .A1(n9582), .A2(n9581), .ZN(N5191) );
  AOI22D1BWP30P140LVT U14101 ( .A1(i_data_bus[553]), .A2(n10567), .B1(
        i_data_bus[585]), .B2(n10565), .ZN(n9584) );
  AOI22D1BWP30P140LVT U14102 ( .A1(i_data_bus[521]), .A2(n10566), .B1(
        i_data_bus[617]), .B2(n10568), .ZN(n9583) );
  ND2D1BWP30P140LVT U14103 ( .A1(n9584), .A2(n9583), .ZN(N5192) );
  AOI22D1BWP30P140LVT U14104 ( .A1(i_data_bus[572]), .A2(n10567), .B1(
        i_data_bus[540]), .B2(n10566), .ZN(n9586) );
  AOI22D1BWP30P140LVT U14105 ( .A1(i_data_bus[604]), .A2(n10565), .B1(
        i_data_bus[636]), .B2(n10568), .ZN(n9585) );
  ND2D1BWP30P140LVT U14106 ( .A1(n9586), .A2(n9585), .ZN(N5211) );
  AOI22D1BWP30P140LVT U14107 ( .A1(i_data_bus[602]), .A2(n10565), .B1(
        i_data_bus[538]), .B2(n10566), .ZN(n9588) );
  AOI22D1BWP30P140LVT U14108 ( .A1(i_data_bus[570]), .A2(n10567), .B1(
        i_data_bus[634]), .B2(n10568), .ZN(n9587) );
  ND2D1BWP30P140LVT U14109 ( .A1(n9588), .A2(n9587), .ZN(N5209) );
  AOI22D1BWP30P140LVT U14110 ( .A1(i_data_bus[593]), .A2(n10565), .B1(
        i_data_bus[529]), .B2(n10566), .ZN(n9590) );
  AOI22D1BWP30P140LVT U14111 ( .A1(i_data_bus[561]), .A2(n10567), .B1(
        i_data_bus[625]), .B2(n10568), .ZN(n9589) );
  ND2D1BWP30P140LVT U14112 ( .A1(n9590), .A2(n9589), .ZN(N5200) );
  AOI22D1BWP30P140LVT U14113 ( .A1(i_data_bus[600]), .A2(n10565), .B1(
        i_data_bus[536]), .B2(n10566), .ZN(n9592) );
  AOI22D1BWP30P140LVT U14114 ( .A1(i_data_bus[568]), .A2(n10567), .B1(
        i_data_bus[632]), .B2(n10568), .ZN(n9591) );
  ND2D1BWP30P140LVT U14115 ( .A1(n9592), .A2(n9591), .ZN(N5207) );
  AOI22D1BWP30P140LVT U14116 ( .A1(i_data_bus[558]), .A2(n10504), .B1(
        i_data_bus[590]), .B2(n10502), .ZN(n9594) );
  AOI22D1BWP30P140LVT U14117 ( .A1(i_data_bus[526]), .A2(n10503), .B1(
        i_data_bus[622]), .B2(n10501), .ZN(n9593) );
  ND2D1BWP30P140LVT U14118 ( .A1(n9594), .A2(n9593), .ZN(N8945) );
  AOI22D1BWP30P140LVT U14119 ( .A1(i_data_bus[548]), .A2(n10504), .B1(
        i_data_bus[580]), .B2(n10502), .ZN(n9596) );
  AOI22D1BWP30P140LVT U14120 ( .A1(i_data_bus[516]), .A2(n10503), .B1(
        i_data_bus[612]), .B2(n10501), .ZN(n9595) );
  ND2D1BWP30P140LVT U14121 ( .A1(n9596), .A2(n9595), .ZN(N8935) );
  AOI22D1BWP30P140LVT U14122 ( .A1(i_data_bus[559]), .A2(n10504), .B1(
        i_data_bus[591]), .B2(n10502), .ZN(n9598) );
  AOI22D1BWP30P140LVT U14123 ( .A1(i_data_bus[527]), .A2(n10503), .B1(
        i_data_bus[623]), .B2(n10501), .ZN(n9597) );
  ND2D1BWP30P140LVT U14124 ( .A1(n9598), .A2(n9597), .ZN(N8946) );
  AOI22D1BWP30P140LVT U14125 ( .A1(i_data_bus[607]), .A2(n10502), .B1(
        i_data_bus[543]), .B2(n10503), .ZN(n9600) );
  AOI22D1BWP30P140LVT U14126 ( .A1(i_data_bus[575]), .A2(n10504), .B1(
        i_data_bus[639]), .B2(n10501), .ZN(n9599) );
  ND2D1BWP30P140LVT U14127 ( .A1(n9600), .A2(n9599), .ZN(N8962) );
  AOI22D1BWP30P140LVT U14128 ( .A1(i_data_bus[593]), .A2(n10502), .B1(
        i_data_bus[529]), .B2(n10503), .ZN(n9602) );
  AOI22D1BWP30P140LVT U14129 ( .A1(i_data_bus[561]), .A2(n10504), .B1(
        i_data_bus[625]), .B2(n10501), .ZN(n9601) );
  ND2D1BWP30P140LVT U14130 ( .A1(n9602), .A2(n9601), .ZN(N8948) );
  AOI22D1BWP30P140LVT U14131 ( .A1(i_data_bus[577]), .A2(n10502), .B1(
        i_data_bus[545]), .B2(n10504), .ZN(n9604) );
  AOI22D1BWP30P140LVT U14132 ( .A1(i_data_bus[513]), .A2(n10503), .B1(
        i_data_bus[609]), .B2(n10501), .ZN(n9603) );
  ND2D1BWP30P140LVT U14133 ( .A1(n9604), .A2(n9603), .ZN(N8932) );
  AOI22D1BWP30P140LVT U14134 ( .A1(i_data_bus[587]), .A2(n10502), .B1(
        i_data_bus[555]), .B2(n10504), .ZN(n9606) );
  AOI22D1BWP30P140LVT U14135 ( .A1(i_data_bus[523]), .A2(n10503), .B1(
        i_data_bus[619]), .B2(n10501), .ZN(n9605) );
  ND2D1BWP30P140LVT U14136 ( .A1(n9606), .A2(n9605), .ZN(N8942) );
  AOI22D1BWP30P140LVT U14137 ( .A1(i_data_bus[549]), .A2(n10504), .B1(
        i_data_bus[581]), .B2(n10502), .ZN(n9608) );
  AOI22D1BWP30P140LVT U14138 ( .A1(i_data_bus[517]), .A2(n10503), .B1(
        i_data_bus[613]), .B2(n10501), .ZN(n9607) );
  ND2D1BWP30P140LVT U14139 ( .A1(n9608), .A2(n9607), .ZN(N8936) );
  AOI22D1BWP30P140LVT U14140 ( .A1(i_data_bus[551]), .A2(n10504), .B1(
        i_data_bus[583]), .B2(n10502), .ZN(n9610) );
  AOI22D1BWP30P140LVT U14141 ( .A1(i_data_bus[519]), .A2(n10503), .B1(
        i_data_bus[615]), .B2(n10501), .ZN(n9609) );
  ND2D1BWP30P140LVT U14142 ( .A1(n9610), .A2(n9609), .ZN(N8938) );
  AOI22D1BWP30P140LVT U14143 ( .A1(i_data_bus[595]), .A2(n10502), .B1(
        i_data_bus[563]), .B2(n10504), .ZN(n9612) );
  AOI22D1BWP30P140LVT U14144 ( .A1(i_data_bus[531]), .A2(n10503), .B1(
        i_data_bus[627]), .B2(n10501), .ZN(n9611) );
  ND2D1BWP30P140LVT U14145 ( .A1(n9612), .A2(n9611), .ZN(N8950) );
  AOI22D1BWP30P140LVT U14146 ( .A1(i_data_bus[1006]), .A2(n10457), .B1(
        i_data_bus[942]), .B2(n10460), .ZN(n9614) );
  AOI22D1BWP30P140LVT U14147 ( .A1(i_data_bus[910]), .A2(n10458), .B1(
        i_data_bus[974]), .B2(n10459), .ZN(n9613) );
  ND2D1BWP30P140LVT U14148 ( .A1(n9614), .A2(n9613), .ZN(N11467) );
  AOI22D1BWP30P140LVT U14149 ( .A1(i_data_bus[896]), .A2(n10458), .B1(
        i_data_bus[992]), .B2(n10457), .ZN(n9616) );
  AOI22D1BWP30P140LVT U14150 ( .A1(i_data_bus[928]), .A2(n10460), .B1(
        i_data_bus[960]), .B2(n10459), .ZN(n9615) );
  ND2D1BWP30P140LVT U14151 ( .A1(n9616), .A2(n9615), .ZN(N11453) );
  AOI22D1BWP30P140LVT U14152 ( .A1(i_data_bus[957]), .A2(n10460), .B1(
        i_data_bus[1021]), .B2(n10457), .ZN(n9618) );
  AOI22D1BWP30P140LVT U14153 ( .A1(i_data_bus[925]), .A2(n10458), .B1(
        i_data_bus[989]), .B2(n10459), .ZN(n9617) );
  ND2D1BWP30P140LVT U14154 ( .A1(n9618), .A2(n9617), .ZN(N11482) );
  AOI22D1BWP30P140LVT U14155 ( .A1(i_data_bus[899]), .A2(n10458), .B1(
        i_data_bus[931]), .B2(n10460), .ZN(n9620) );
  AOI22D1BWP30P140LVT U14156 ( .A1(i_data_bus[995]), .A2(n10457), .B1(
        i_data_bus[963]), .B2(n10459), .ZN(n9619) );
  ND2D1BWP30P140LVT U14157 ( .A1(n9620), .A2(n9619), .ZN(N11456) );
  AOI22D1BWP30P140LVT U14158 ( .A1(i_data_bus[993]), .A2(n10457), .B1(
        i_data_bus[897]), .B2(n10458), .ZN(n9622) );
  AOI22D1BWP30P140LVT U14159 ( .A1(i_data_bus[929]), .A2(n10460), .B1(
        i_data_bus[961]), .B2(n10459), .ZN(n9621) );
  ND2D1BWP30P140LVT U14160 ( .A1(n9622), .A2(n9621), .ZN(N11454) );
  AOI22D1BWP30P140LVT U14161 ( .A1(i_data_bus[1018]), .A2(n10457), .B1(
        i_data_bus[922]), .B2(n10458), .ZN(n9624) );
  AOI22D1BWP30P140LVT U14162 ( .A1(i_data_bus[954]), .A2(n10460), .B1(
        i_data_bus[986]), .B2(n10459), .ZN(n9623) );
  ND2D1BWP30P140LVT U14163 ( .A1(n9624), .A2(n9623), .ZN(N11479) );
  AOI22D1BWP30P140LVT U14164 ( .A1(i_data_bus[998]), .A2(n10457), .B1(
        i_data_bus[902]), .B2(n10458), .ZN(n9626) );
  AOI22D1BWP30P140LVT U14165 ( .A1(i_data_bus[934]), .A2(n10460), .B1(
        i_data_bus[966]), .B2(n10459), .ZN(n9625) );
  ND2D1BWP30P140LVT U14166 ( .A1(n9626), .A2(n9625), .ZN(N11459) );
  AOI22D1BWP30P140LVT U14167 ( .A1(i_data_bus[903]), .A2(n10458), .B1(
        i_data_bus[999]), .B2(n10457), .ZN(n9628) );
  AOI22D1BWP30P140LVT U14168 ( .A1(i_data_bus[935]), .A2(n10460), .B1(
        i_data_bus[967]), .B2(n10459), .ZN(n9627) );
  ND2D1BWP30P140LVT U14169 ( .A1(n9628), .A2(n9627), .ZN(N11460) );
  AOI22D1BWP30P140LVT U14170 ( .A1(i_data_bus[950]), .A2(n10460), .B1(
        i_data_bus[918]), .B2(n10458), .ZN(n9630) );
  AOI22D1BWP30P140LVT U14171 ( .A1(i_data_bus[1014]), .A2(n10457), .B1(
        i_data_bus[982]), .B2(n10459), .ZN(n9629) );
  ND2D1BWP30P140LVT U14172 ( .A1(n9630), .A2(n9629), .ZN(N11475) );
  AOI22D1BWP30P140LVT U14173 ( .A1(i_data_bus[601]), .A2(n10600), .B1(
        i_data_bus[537]), .B2(n10597), .ZN(n9632) );
  AOI22D1BWP30P140LVT U14174 ( .A1(i_data_bus[569]), .A2(n10598), .B1(
        i_data_bus[633]), .B2(n10599), .ZN(n9631) );
  ND2D1BWP30P140LVT U14175 ( .A1(n9632), .A2(n9631), .ZN(N3334) );
  AOI22D1BWP30P140LVT U14176 ( .A1(i_data_bus[559]), .A2(n10598), .B1(
        i_data_bus[527]), .B2(n10597), .ZN(n9634) );
  AOI22D1BWP30P140LVT U14177 ( .A1(i_data_bus[591]), .A2(n10600), .B1(
        i_data_bus[623]), .B2(n10599), .ZN(n9633) );
  ND2D1BWP30P140LVT U14178 ( .A1(n9634), .A2(n9633), .ZN(N3324) );
  AOI22D1BWP30P140LVT U14179 ( .A1(i_data_bus[61]), .A2(n10518), .B1(
        i_data_bus[125]), .B2(n10519), .ZN(n9636) );
  AOI22D1BWP30P140LVT U14180 ( .A1(i_data_bus[93]), .A2(n10517), .B1(
        i_data_bus[29]), .B2(n10520), .ZN(n9635) );
  ND2D1BWP30P140LVT U14181 ( .A1(n9636), .A2(n9635), .ZN(N8096) );
  AOI22D1BWP30P140LVT U14182 ( .A1(i_data_bus[592]), .A2(n10600), .B1(
        i_data_bus[528]), .B2(n10597), .ZN(n9638) );
  AOI22D1BWP30P140LVT U14183 ( .A1(i_data_bus[560]), .A2(n10598), .B1(
        i_data_bus[624]), .B2(n10599), .ZN(n9637) );
  ND2D1BWP30P140LVT U14184 ( .A1(n9638), .A2(n9637), .ZN(N3325) );
  AOI22D1BWP30P140LVT U14185 ( .A1(i_data_bus[533]), .A2(n10597), .B1(
        i_data_bus[565]), .B2(n10598), .ZN(n9640) );
  AOI22D1BWP30P140LVT U14186 ( .A1(i_data_bus[597]), .A2(n10600), .B1(
        i_data_bus[629]), .B2(n10599), .ZN(n9639) );
  ND2D1BWP30P140LVT U14187 ( .A1(n9640), .A2(n9639), .ZN(N3330) );
  AOI22D1BWP30P140LVT U14188 ( .A1(i_data_bus[523]), .A2(n10597), .B1(
        i_data_bus[555]), .B2(n10598), .ZN(n9642) );
  AOI22D1BWP30P140LVT U14189 ( .A1(i_data_bus[587]), .A2(n10600), .B1(
        i_data_bus[619]), .B2(n10599), .ZN(n9641) );
  ND2D1BWP30P140LVT U14190 ( .A1(n9642), .A2(n9641), .ZN(N3320) );
  AOI22D1BWP30P140LVT U14191 ( .A1(i_data_bus[607]), .A2(n10600), .B1(
        i_data_bus[543]), .B2(n10597), .ZN(n9644) );
  AOI22D1BWP30P140LVT U14192 ( .A1(i_data_bus[575]), .A2(n10598), .B1(
        i_data_bus[639]), .B2(n10599), .ZN(n9643) );
  ND2D1BWP30P140LVT U14193 ( .A1(n9644), .A2(n9643), .ZN(N3340) );
  AOI22D1BWP30P140LVT U14194 ( .A1(i_data_bus[549]), .A2(n10598), .B1(
        i_data_bus[581]), .B2(n10600), .ZN(n9646) );
  AOI22D1BWP30P140LVT U14195 ( .A1(i_data_bus[517]), .A2(n10597), .B1(
        i_data_bus[613]), .B2(n10599), .ZN(n9645) );
  ND2D1BWP30P140LVT U14196 ( .A1(n9646), .A2(n9645), .ZN(N3314) );
  AOI22D1BWP30P140LVT U14197 ( .A1(i_data_bus[123]), .A2(n10519), .B1(
        i_data_bus[91]), .B2(n10517), .ZN(n9648) );
  AOI22D1BWP30P140LVT U14198 ( .A1(i_data_bus[59]), .A2(n10518), .B1(
        i_data_bus[27]), .B2(n10520), .ZN(n9647) );
  ND2D1BWP30P140LVT U14199 ( .A1(n9648), .A2(n9647), .ZN(N8094) );
  AOI22D1BWP30P140LVT U14200 ( .A1(i_data_bus[88]), .A2(n10517), .B1(
        i_data_bus[56]), .B2(n10518), .ZN(n9650) );
  AOI22D1BWP30P140LVT U14201 ( .A1(i_data_bus[120]), .A2(n10519), .B1(
        i_data_bus[24]), .B2(n10520), .ZN(n9649) );
  ND2D1BWP30P140LVT U14202 ( .A1(n9650), .A2(n9649), .ZN(N8091) );
  AOI22D1BWP30P140LVT U14203 ( .A1(i_data_bus[106]), .A2(n10519), .B1(
        i_data_bus[42]), .B2(n10518), .ZN(n9652) );
  AOI22D1BWP30P140LVT U14204 ( .A1(i_data_bus[74]), .A2(n10517), .B1(
        i_data_bus[10]), .B2(n10520), .ZN(n9651) );
  ND2D1BWP30P140LVT U14205 ( .A1(n9652), .A2(n9651), .ZN(N8077) );
  AOI22D1BWP30P140LVT U14206 ( .A1(i_data_bus[118]), .A2(n10519), .B1(
        i_data_bus[54]), .B2(n10518), .ZN(n9654) );
  AOI22D1BWP30P140LVT U14207 ( .A1(i_data_bus[86]), .A2(n10517), .B1(
        i_data_bus[22]), .B2(n10520), .ZN(n9653) );
  ND2D1BWP30P140LVT U14208 ( .A1(n9654), .A2(n9653), .ZN(N8089) );
  AOI22D1BWP30P140LVT U14209 ( .A1(i_data_bus[53]), .A2(n10518), .B1(
        i_data_bus[85]), .B2(n10517), .ZN(n9656) );
  AOI22D1BWP30P140LVT U14210 ( .A1(i_data_bus[117]), .A2(n10519), .B1(
        i_data_bus[21]), .B2(n10520), .ZN(n9655) );
  ND2D1BWP30P140LVT U14211 ( .A1(n9656), .A2(n9655), .ZN(N8088) );
  AOI22D1BWP30P140LVT U14212 ( .A1(i_data_bus[51]), .A2(n10518), .B1(
        i_data_bus[115]), .B2(n10519), .ZN(n9658) );
  AOI22D1BWP30P140LVT U14213 ( .A1(i_data_bus[83]), .A2(n10517), .B1(
        i_data_bus[19]), .B2(n10520), .ZN(n9657) );
  ND2D1BWP30P140LVT U14214 ( .A1(n9658), .A2(n9657), .ZN(N8086) );
  AOI22D1BWP30P140LVT U14215 ( .A1(i_data_bus[109]), .A2(n10519), .B1(
        i_data_bus[45]), .B2(n10518), .ZN(n9660) );
  AOI22D1BWP30P140LVT U14216 ( .A1(i_data_bus[77]), .A2(n10517), .B1(
        i_data_bus[13]), .B2(n10520), .ZN(n9659) );
  ND2D1BWP30P140LVT U14217 ( .A1(n9660), .A2(n9659), .ZN(N8080) );
  AOI22D1BWP30P140LVT U14218 ( .A1(i_data_bus[33]), .A2(n10518), .B1(
        i_data_bus[97]), .B2(n10519), .ZN(n9662) );
  AOI22D1BWP30P140LVT U14219 ( .A1(i_data_bus[65]), .A2(n10517), .B1(
        i_data_bus[1]), .B2(n10520), .ZN(n9661) );
  ND2D1BWP30P140LVT U14220 ( .A1(n9662), .A2(n9661), .ZN(N8068) );
  AOI22D1BWP30P140LVT U14221 ( .A1(i_data_bus[32]), .A2(n10518), .B1(
        i_data_bus[64]), .B2(n10517), .ZN(n9664) );
  AOI22D1BWP30P140LVT U14222 ( .A1(i_data_bus[96]), .A2(n10519), .B1(
        i_data_bus[0]), .B2(n10520), .ZN(n9663) );
  ND2D1BWP30P140LVT U14223 ( .A1(n9664), .A2(n9663), .ZN(N8067) );
  AOI22D1BWP30P140LVT U14224 ( .A1(i_data_bus[69]), .A2(n10517), .B1(
        i_data_bus[101]), .B2(n10519), .ZN(n9666) );
  AOI22D1BWP30P140LVT U14225 ( .A1(i_data_bus[37]), .A2(n10518), .B1(
        i_data_bus[5]), .B2(n10520), .ZN(n9665) );
  ND2D1BWP30P140LVT U14226 ( .A1(n9666), .A2(n9665), .ZN(N8072) );
  AOI22D1BWP30P140LVT U14227 ( .A1(i_data_bus[39]), .A2(n10518), .B1(
        i_data_bus[71]), .B2(n10517), .ZN(n9668) );
  AOI22D1BWP30P140LVT U14228 ( .A1(i_data_bus[103]), .A2(n10519), .B1(
        i_data_bus[7]), .B2(n10520), .ZN(n9667) );
  ND2D1BWP30P140LVT U14229 ( .A1(n9668), .A2(n9667), .ZN(N8074) );
  AOI22D1BWP30P140LVT U14230 ( .A1(i_data_bus[89]), .A2(n10517), .B1(
        i_data_bus[57]), .B2(n10518), .ZN(n9670) );
  AOI22D1BWP30P140LVT U14231 ( .A1(i_data_bus[121]), .A2(n10519), .B1(
        i_data_bus[25]), .B2(n10520), .ZN(n9669) );
  ND2D1BWP30P140LVT U14232 ( .A1(n9670), .A2(n9669), .ZN(N8092) );
  AOI22D1BWP30P140LVT U14233 ( .A1(i_data_bus[67]), .A2(n10517), .B1(
        i_data_bus[99]), .B2(n10519), .ZN(n9672) );
  AOI22D1BWP30P140LVT U14234 ( .A1(i_data_bus[35]), .A2(n10518), .B1(
        i_data_bus[3]), .B2(n10520), .ZN(n9671) );
  ND2D1BWP30P140LVT U14235 ( .A1(n9672), .A2(n9671), .ZN(N8070) );
  AOI22D1BWP30P140LVT U14236 ( .A1(i_data_bus[592]), .A2(n10437), .B1(
        i_data_bus[528]), .B2(n10438), .ZN(n9674) );
  AOI22D1BWP30P140LVT U14237 ( .A1(i_data_bus[560]), .A2(n10439), .B1(
        i_data_bus[624]), .B2(n10440), .ZN(n9673) );
  ND2D1BWP30P140LVT U14238 ( .A1(n9674), .A2(n9673), .ZN(N12695) );
  AOI22D1BWP30P140LVT U14239 ( .A1(i_data_bus[543]), .A2(n10438), .B1(
        i_data_bus[575]), .B2(n10439), .ZN(n9676) );
  AOI22D1BWP30P140LVT U14240 ( .A1(i_data_bus[607]), .A2(n10437), .B1(
        i_data_bus[639]), .B2(n10440), .ZN(n9675) );
  ND2D1BWP30P140LVT U14241 ( .A1(n9676), .A2(n9675), .ZN(N12710) );
  AOI22D1BWP30P140LVT U14242 ( .A1(i_data_bus[570]), .A2(n10439), .B1(
        i_data_bus[538]), .B2(n10438), .ZN(n9678) );
  AOI22D1BWP30P140LVT U14243 ( .A1(i_data_bus[602]), .A2(n10437), .B1(
        i_data_bus[634]), .B2(n10440), .ZN(n9677) );
  ND2D1BWP30P140LVT U14244 ( .A1(n9678), .A2(n9677), .ZN(N12705) );
  AOI22D1BWP30P140LVT U14245 ( .A1(i_data_bus[564]), .A2(n10439), .B1(
        i_data_bus[532]), .B2(n10438), .ZN(n9680) );
  AOI22D1BWP30P140LVT U14246 ( .A1(i_data_bus[596]), .A2(n10437), .B1(
        i_data_bus[628]), .B2(n10440), .ZN(n9679) );
  ND2D1BWP30P140LVT U14247 ( .A1(n9680), .A2(n9679), .ZN(N12699) );
  AOI22D1BWP30P140LVT U14248 ( .A1(i_data_bus[282]), .A2(n10543), .B1(
        i_data_bus[346]), .B2(n10544), .ZN(n9682) );
  AOI22D1BWP30P140LVT U14249 ( .A1(i_data_bus[314]), .A2(n10541), .B1(
        i_data_bus[378]), .B2(n10542), .ZN(n9681) );
  ND2D1BWP30P140LVT U14250 ( .A1(n9682), .A2(n9681), .ZN(N6651) );
  AOI22D1BWP30P140LVT U14251 ( .A1(i_data_bus[271]), .A2(n10543), .B1(
        i_data_bus[335]), .B2(n10544), .ZN(n9684) );
  AOI22D1BWP30P140LVT U14252 ( .A1(i_data_bus[303]), .A2(n10541), .B1(
        i_data_bus[367]), .B2(n10542), .ZN(n9683) );
  ND2D1BWP30P140LVT U14253 ( .A1(n9684), .A2(n9683), .ZN(N6640) );
  AOI22D1BWP30P140LVT U14254 ( .A1(i_data_bus[265]), .A2(n10543), .B1(
        i_data_bus[329]), .B2(n10544), .ZN(n9686) );
  AOI22D1BWP30P140LVT U14255 ( .A1(i_data_bus[297]), .A2(n10541), .B1(
        i_data_bus[361]), .B2(n10542), .ZN(n9685) );
  ND2D1BWP30P140LVT U14256 ( .A1(n9686), .A2(n9685), .ZN(N6634) );
  AOI22D1BWP30P140LVT U14257 ( .A1(i_data_bus[281]), .A2(n10543), .B1(
        i_data_bus[345]), .B2(n10544), .ZN(n9688) );
  AOI22D1BWP30P140LVT U14258 ( .A1(i_data_bus[313]), .A2(n10541), .B1(
        i_data_bus[377]), .B2(n10542), .ZN(n9687) );
  ND2D1BWP30P140LVT U14259 ( .A1(n9688), .A2(n9687), .ZN(N6650) );
  AOI22D1BWP30P140LVT U14260 ( .A1(i_data_bus[328]), .A2(n10544), .B1(
        i_data_bus[264]), .B2(n10543), .ZN(n9690) );
  AOI22D1BWP30P140LVT U14261 ( .A1(i_data_bus[296]), .A2(n10541), .B1(
        i_data_bus[360]), .B2(n10542), .ZN(n9689) );
  ND2D1BWP30P140LVT U14262 ( .A1(n9690), .A2(n9689), .ZN(N6633) );
  AOI22D1BWP30P140LVT U14263 ( .A1(i_data_bus[310]), .A2(n10541), .B1(
        i_data_bus[342]), .B2(n10544), .ZN(n9692) );
  AOI22D1BWP30P140LVT U14264 ( .A1(i_data_bus[278]), .A2(n10543), .B1(
        i_data_bus[374]), .B2(n10542), .ZN(n9691) );
  ND2D1BWP30P140LVT U14265 ( .A1(n9692), .A2(n9691), .ZN(N6647) );
  AOI22D1BWP30P140LVT U14266 ( .A1(i_data_bus[309]), .A2(n10541), .B1(
        i_data_bus[277]), .B2(n10543), .ZN(n9694) );
  AOI22D1BWP30P140LVT U14267 ( .A1(i_data_bus[341]), .A2(n10544), .B1(
        i_data_bus[373]), .B2(n10542), .ZN(n9693) );
  ND2D1BWP30P140LVT U14268 ( .A1(n9694), .A2(n9693), .ZN(N6646) );
  AOI22D1BWP30P140LVT U14269 ( .A1(i_data_bus[349]), .A2(n10544), .B1(
        i_data_bus[285]), .B2(n10543), .ZN(n9696) );
  AOI22D1BWP30P140LVT U14270 ( .A1(i_data_bus[317]), .A2(n10541), .B1(
        i_data_bus[381]), .B2(n10542), .ZN(n9695) );
  ND2D1BWP30P140LVT U14271 ( .A1(n9696), .A2(n9695), .ZN(N6654) );
  AOI22D1BWP30P140LVT U14272 ( .A1(i_data_bus[299]), .A2(n10541), .B1(
        i_data_bus[331]), .B2(n10544), .ZN(n9698) );
  AOI22D1BWP30P140LVT U14273 ( .A1(i_data_bus[267]), .A2(n10543), .B1(
        i_data_bus[363]), .B2(n10542), .ZN(n9697) );
  ND2D1BWP30P140LVT U14274 ( .A1(n9698), .A2(n9697), .ZN(N6636) );
  AOI22D1BWP30P140LVT U14275 ( .A1(i_data_bus[347]), .A2(n10544), .B1(
        i_data_bus[283]), .B2(n10543), .ZN(n9700) );
  AOI22D1BWP30P140LVT U14276 ( .A1(i_data_bus[315]), .A2(n10541), .B1(
        i_data_bus[379]), .B2(n10542), .ZN(n9699) );
  ND2D1BWP30P140LVT U14277 ( .A1(n9700), .A2(n9699), .ZN(N6652) );
  AOI22D1BWP30P140LVT U14278 ( .A1(i_data_bus[351]), .A2(n10478), .B1(
        i_data_bus[319]), .B2(n10477), .ZN(n9702) );
  AOI22D1BWP30P140LVT U14279 ( .A1(i_data_bus[287]), .A2(n10480), .B1(
        i_data_bus[383]), .B2(n10479), .ZN(n9701) );
  ND2D1BWP30P140LVT U14280 ( .A1(n9702), .A2(n9701), .ZN(N10404) );
  AOI22D1BWP30P140LVT U14281 ( .A1(i_data_bus[311]), .A2(n10477), .B1(
        i_data_bus[343]), .B2(n10478), .ZN(n9704) );
  AOI22D1BWP30P140LVT U14282 ( .A1(i_data_bus[279]), .A2(n10480), .B1(
        i_data_bus[375]), .B2(n10479), .ZN(n9703) );
  ND2D1BWP30P140LVT U14283 ( .A1(n9704), .A2(n9703), .ZN(N10396) );
  AOI22D1BWP30P140LVT U14284 ( .A1(i_data_bus[328]), .A2(n10478), .B1(
        i_data_bus[264]), .B2(n10480), .ZN(n9706) );
  AOI22D1BWP30P140LVT U14285 ( .A1(i_data_bus[296]), .A2(n10477), .B1(
        i_data_bus[360]), .B2(n10479), .ZN(n9705) );
  ND2D1BWP30P140LVT U14286 ( .A1(n9706), .A2(n9705), .ZN(N10381) );
  AOI22D1BWP30P140LVT U14287 ( .A1(i_data_bus[293]), .A2(n10477), .B1(
        i_data_bus[261]), .B2(n10480), .ZN(n9708) );
  AOI22D1BWP30P140LVT U14288 ( .A1(i_data_bus[325]), .A2(n10478), .B1(
        i_data_bus[357]), .B2(n10479), .ZN(n9707) );
  ND2D1BWP30P140LVT U14289 ( .A1(n9708), .A2(n9707), .ZN(N10378) );
  AOI22D1BWP30P140LVT U14290 ( .A1(i_data_bus[265]), .A2(n10480), .B1(
        i_data_bus[329]), .B2(n10478), .ZN(n9710) );
  AOI22D1BWP30P140LVT U14291 ( .A1(i_data_bus[297]), .A2(n10477), .B1(
        i_data_bus[361]), .B2(n10479), .ZN(n9709) );
  ND2D1BWP30P140LVT U14292 ( .A1(n9710), .A2(n9709), .ZN(N10382) );
  AOI22D1BWP30P140LVT U14293 ( .A1(i_data_bus[349]), .A2(n10478), .B1(
        i_data_bus[285]), .B2(n10480), .ZN(n9712) );
  AOI22D1BWP30P140LVT U14294 ( .A1(i_data_bus[317]), .A2(n10477), .B1(
        i_data_bus[381]), .B2(n10479), .ZN(n9711) );
  ND2D1BWP30P140LVT U14295 ( .A1(n9712), .A2(n9711), .ZN(N10402) );
  AOI22D1BWP30P140LVT U14296 ( .A1(i_data_bus[271]), .A2(n10480), .B1(
        i_data_bus[335]), .B2(n10478), .ZN(n9714) );
  AOI22D1BWP30P140LVT U14297 ( .A1(i_data_bus[303]), .A2(n10477), .B1(
        i_data_bus[367]), .B2(n10479), .ZN(n9713) );
  ND2D1BWP30P140LVT U14298 ( .A1(n9714), .A2(n9713), .ZN(N10388) );
  AOI22D1BWP30P140LVT U14299 ( .A1(i_data_bus[258]), .A2(n10480), .B1(
        i_data_bus[290]), .B2(n10477), .ZN(n9716) );
  AOI22D1BWP30P140LVT U14300 ( .A1(i_data_bus[322]), .A2(n10478), .B1(
        i_data_bus[354]), .B2(n10479), .ZN(n9715) );
  ND2D1BWP30P140LVT U14301 ( .A1(n9716), .A2(n9715), .ZN(N10375) );
  AOI22D1BWP30P140LVT U14302 ( .A1(i_data_bus[321]), .A2(n10478), .B1(
        i_data_bus[289]), .B2(n10477), .ZN(n9718) );
  AOI22D1BWP30P140LVT U14303 ( .A1(i_data_bus[257]), .A2(n10480), .B1(
        i_data_bus[353]), .B2(n10479), .ZN(n9717) );
  ND2D1BWP30P140LVT U14304 ( .A1(n9718), .A2(n9717), .ZN(N10374) );
  AOI22D1BWP30P140LVT U14305 ( .A1(i_data_bus[275]), .A2(n10415), .B1(
        i_data_bus[339]), .B2(n10413), .ZN(n9720) );
  AOI22D1BWP30P140LVT U14306 ( .A1(i_data_bus[307]), .A2(n10414), .B1(
        i_data_bus[371]), .B2(n10416), .ZN(n9719) );
  ND2D1BWP30P140LVT U14307 ( .A1(n9720), .A2(n9719), .ZN(N14140) );
  AOI22D1BWP30P140LVT U14308 ( .A1(i_data_bus[309]), .A2(n10414), .B1(
        i_data_bus[277]), .B2(n10415), .ZN(n9722) );
  AOI22D1BWP30P140LVT U14309 ( .A1(i_data_bus[341]), .A2(n10413), .B1(
        i_data_bus[373]), .B2(n10416), .ZN(n9721) );
  ND2D1BWP30P140LVT U14310 ( .A1(n9722), .A2(n9721), .ZN(N14142) );
  AOI22D1BWP30P140LVT U14311 ( .A1(i_data_bus[347]), .A2(n10413), .B1(
        i_data_bus[283]), .B2(n10415), .ZN(n9724) );
  AOI22D1BWP30P140LVT U14312 ( .A1(i_data_bus[315]), .A2(n10414), .B1(
        i_data_bus[379]), .B2(n10416), .ZN(n9723) );
  ND2D1BWP30P140LVT U14313 ( .A1(n9724), .A2(n9723), .ZN(N14148) );
  AOI22D1BWP30P140LVT U14314 ( .A1(i_data_bus[327]), .A2(n10413), .B1(
        i_data_bus[263]), .B2(n10415), .ZN(n9726) );
  AOI22D1BWP30P140LVT U14315 ( .A1(i_data_bus[295]), .A2(n10414), .B1(
        i_data_bus[359]), .B2(n10416), .ZN(n9725) );
  ND2D1BWP30P140LVT U14316 ( .A1(n9726), .A2(n9725), .ZN(N14128) );
  AOI22D1BWP30P140LVT U14317 ( .A1(i_data_bus[287]), .A2(n10415), .B1(
        i_data_bus[319]), .B2(n10414), .ZN(n9728) );
  AOI22D1BWP30P140LVT U14318 ( .A1(i_data_bus[351]), .A2(n10413), .B1(
        i_data_bus[383]), .B2(n10416), .ZN(n9727) );
  ND2D1BWP30P140LVT U14319 ( .A1(n9728), .A2(n9727), .ZN(N14152) );
  AOI22D1BWP30P140LVT U14320 ( .A1(i_data_bus[279]), .A2(n10415), .B1(
        i_data_bus[343]), .B2(n10413), .ZN(n9730) );
  AOI22D1BWP30P140LVT U14321 ( .A1(i_data_bus[311]), .A2(n10414), .B1(
        i_data_bus[375]), .B2(n10416), .ZN(n9729) );
  ND2D1BWP30P140LVT U14322 ( .A1(n9730), .A2(n9729), .ZN(N14144) );
  AOI22D1BWP30P140LVT U14323 ( .A1(i_data_bus[265]), .A2(n10415), .B1(
        i_data_bus[297]), .B2(n10414), .ZN(n9732) );
  AOI22D1BWP30P140LVT U14324 ( .A1(i_data_bus[329]), .A2(n10413), .B1(
        i_data_bus[361]), .B2(n10416), .ZN(n9731) );
  ND2D1BWP30P140LVT U14325 ( .A1(n9732), .A2(n9731), .ZN(N14130) );
  AOI22D1BWP30P140LVT U14326 ( .A1(i_data_bus[330]), .A2(n10413), .B1(
        i_data_bus[298]), .B2(n10414), .ZN(n9734) );
  AOI22D1BWP30P140LVT U14327 ( .A1(i_data_bus[266]), .A2(n10415), .B1(
        i_data_bus[362]), .B2(n10416), .ZN(n9733) );
  ND2D1BWP30P140LVT U14328 ( .A1(n9734), .A2(n9733), .ZN(N14131) );
  AOI22D1BWP30P140LVT U14329 ( .A1(i_data_bus[310]), .A2(n10414), .B1(
        i_data_bus[278]), .B2(n10415), .ZN(n9736) );
  AOI22D1BWP30P140LVT U14330 ( .A1(i_data_bus[342]), .A2(n10413), .B1(
        i_data_bus[374]), .B2(n10416), .ZN(n9735) );
  ND2D1BWP30P140LVT U14331 ( .A1(n9736), .A2(n9735), .ZN(N14143) );
  AOI22D1BWP30P140LVT U14332 ( .A1(i_data_bus[313]), .A2(n10414), .B1(
        i_data_bus[345]), .B2(n10413), .ZN(n9738) );
  AOI22D1BWP30P140LVT U14333 ( .A1(i_data_bus[281]), .A2(n10415), .B1(
        i_data_bus[377]), .B2(n10416), .ZN(n9737) );
  ND2D1BWP30P140LVT U14334 ( .A1(n9738), .A2(n9737), .ZN(N14146) );
  AOI22D1BWP30P140LVT U14335 ( .A1(i_data_bus[273]), .A2(n10415), .B1(
        i_data_bus[337]), .B2(n10413), .ZN(n9740) );
  AOI22D1BWP30P140LVT U14336 ( .A1(i_data_bus[305]), .A2(n10414), .B1(
        i_data_bus[369]), .B2(n10416), .ZN(n9739) );
  ND2D1BWP30P140LVT U14337 ( .A1(n9740), .A2(n9739), .ZN(N14138) );
  NR4D1BWP30P140LVT U14338 ( .A1(i_cmd[192]), .A2(n9746), .A3(n9741), .A4(
        n9742), .ZN(n10623) );
  INR4D1BWP30P140LVT U14339 ( .A1(i_cmd[200]), .B1(i_cmd[216]), .B2(n9743), 
        .B3(n9748), .ZN(n10622) );
  AOI22D1BWP30P140LVT U14340 ( .A1(n10623), .A2(i_data_bus[853]), .B1(n10622), 
        .B2(i_data_bus[821]), .ZN(n9751) );
  NR4D1BWP30P140LVT U14341 ( .A1(i_cmd[208]), .A2(n9746), .A3(n9745), .A4(
        n9744), .ZN(n10621) );
  AOI22D1BWP30P140LVT U14342 ( .A1(n10621), .A2(i_data_bus[789]), .B1(n9749), 
        .B2(i_data_bus[885]), .ZN(n9750) );
  ND2D1BWP30P140LVT U14343 ( .A1(n9751), .A2(n9750), .ZN(N1884) );
  AOI22D1BWP30P140LVT U14344 ( .A1(n10623), .A2(i_data_bus[847]), .B1(n10622), 
        .B2(i_data_bus[815]), .ZN(n9753) );
  AOI22D1BWP30P140LVT U14345 ( .A1(n10621), .A2(i_data_bus[783]), .B1(n9749), 
        .B2(i_data_bus[879]), .ZN(n9752) );
  ND2D1BWP30P140LVT U14346 ( .A1(n9753), .A2(n9752), .ZN(N1878) );
  AOI22D1BWP30P140LVT U14347 ( .A1(n10623), .A2(i_data_bus[835]), .B1(n10622), 
        .B2(i_data_bus[803]), .ZN(n9755) );
  AOI22D1BWP30P140LVT U14348 ( .A1(n10621), .A2(i_data_bus[771]), .B1(n9749), 
        .B2(i_data_bus[867]), .ZN(n9754) );
  ND2D1BWP30P140LVT U14349 ( .A1(n9755), .A2(n9754), .ZN(N1866) );
  AOI22D1BWP30P140LVT U14350 ( .A1(n10623), .A2(i_data_bus[851]), .B1(n10622), 
        .B2(i_data_bus[819]), .ZN(n9757) );
  AOI22D1BWP30P140LVT U14351 ( .A1(n10621), .A2(i_data_bus[787]), .B1(n9749), 
        .B2(i_data_bus[883]), .ZN(n9756) );
  ND2D1BWP30P140LVT U14352 ( .A1(n9757), .A2(n9756), .ZN(N1882) );
  NR4D1BWP30P140LVT U14353 ( .A1(i_cmd[112]), .A2(n9762), .A3(n9758), .A4(
        n9759), .ZN(n10634) );
  INR4D1BWP30P140LVT U14354 ( .A1(i_cmd[104]), .B1(i_cmd[120]), .B2(n9760), 
        .B3(n9765), .ZN(n10633) );
  AOI22D1BWP30P140LVT U14355 ( .A1(n10634), .A2(i_data_bus[393]), .B1(n10633), 
        .B2(i_data_bus[425]), .ZN(n9768) );
  NR4D1BWP30P140LVT U14356 ( .A1(i_cmd[96]), .A2(n9763), .A3(n9762), .A4(n9761), .ZN(n10632) );
  AOI22D1BWP30P140LVT U14357 ( .A1(n10632), .A2(i_data_bus[457]), .B1(n9766), 
        .B2(i_data_bus[489]), .ZN(n9767) );
  ND2D1BWP30P140LVT U14358 ( .A1(n9768), .A2(n9767), .ZN(N1212) );
  AOI22D1BWP30P140LVT U14359 ( .A1(n10634), .A2(i_data_bus[391]), .B1(n10633), 
        .B2(i_data_bus[423]), .ZN(n9770) );
  AOI22D1BWP30P140LVT U14360 ( .A1(n10632), .A2(i_data_bus[455]), .B1(n9766), 
        .B2(i_data_bus[487]), .ZN(n9769) );
  ND2D1BWP30P140LVT U14361 ( .A1(n9770), .A2(n9769), .ZN(N1210) );
  AOI22D1BWP30P140LVT U14362 ( .A1(n10634), .A2(i_data_bus[394]), .B1(n10633), 
        .B2(i_data_bus[426]), .ZN(n9772) );
  AOI22D1BWP30P140LVT U14363 ( .A1(n10632), .A2(i_data_bus[458]), .B1(n9766), 
        .B2(i_data_bus[490]), .ZN(n9771) );
  ND2D1BWP30P140LVT U14364 ( .A1(n9772), .A2(n9771), .ZN(N1213) );
  AOI22D1BWP30P140LVT U14365 ( .A1(n10634), .A2(i_data_bus[403]), .B1(n10633), 
        .B2(i_data_bus[435]), .ZN(n9774) );
  AOI22D1BWP30P140LVT U14366 ( .A1(n10632), .A2(i_data_bus[467]), .B1(n9766), 
        .B2(i_data_bus[499]), .ZN(n9773) );
  ND2D1BWP30P140LVT U14367 ( .A1(n9774), .A2(n9773), .ZN(N1222) );
  AOI22D1BWP30P140LVT U14368 ( .A1(n10634), .A2(i_data_bus[396]), .B1(n10633), 
        .B2(i_data_bus[428]), .ZN(n9776) );
  AOI22D1BWP30P140LVT U14369 ( .A1(n10632), .A2(i_data_bus[460]), .B1(n9766), 
        .B2(i_data_bus[492]), .ZN(n9775) );
  ND2D1BWP30P140LVT U14370 ( .A1(n9776), .A2(n9775), .ZN(N1215) );
  AOI22D1BWP30P140LVT U14371 ( .A1(n10634), .A2(i_data_bus[387]), .B1(n10633), 
        .B2(i_data_bus[419]), .ZN(n9778) );
  AOI22D1BWP30P140LVT U14372 ( .A1(n10632), .A2(i_data_bus[451]), .B1(n9766), 
        .B2(i_data_bus[483]), .ZN(n9777) );
  ND2D1BWP30P140LVT U14373 ( .A1(n9778), .A2(n9777), .ZN(N1206) );
  AOI22D1BWP30P140LVT U14374 ( .A1(i_data_bus[768]), .A2(n10621), .B1(
        i_data_bus[864]), .B2(n9749), .ZN(n9780) );
  AOI22D1BWP30P140LVT U14375 ( .A1(i_data_bus[832]), .A2(n10623), .B1(
        i_data_bus[800]), .B2(n10622), .ZN(n9779) );
  ND2D1BWP30P140LVT U14376 ( .A1(n9780), .A2(n9779), .ZN(N1863) );
  AOI22D1BWP30P140LVT U14377 ( .A1(n10633), .A2(i_data_bus[442]), .B1(n10632), 
        .B2(i_data_bus[474]), .ZN(n9782) );
  AOI22D1BWP30P140LVT U14378 ( .A1(n10634), .A2(i_data_bus[410]), .B1(n9766), 
        .B2(i_data_bus[506]), .ZN(n9781) );
  ND2D1BWP30P140LVT U14379 ( .A1(n9782), .A2(n9781), .ZN(N1229) );
  AOI22D1BWP30P140LVT U14380 ( .A1(n10633), .A2(i_data_bus[445]), .B1(n10632), 
        .B2(i_data_bus[477]), .ZN(n9784) );
  AOI22D1BWP30P140LVT U14381 ( .A1(n10634), .A2(i_data_bus[413]), .B1(n9766), 
        .B2(i_data_bus[509]), .ZN(n9783) );
  ND2D1BWP30P140LVT U14382 ( .A1(n9784), .A2(n9783), .ZN(N1232) );
  AOI22D1BWP30P140LVT U14383 ( .A1(n10633), .A2(i_data_bus[438]), .B1(n10632), 
        .B2(i_data_bus[470]), .ZN(n9786) );
  AOI22D1BWP30P140LVT U14384 ( .A1(n10634), .A2(i_data_bus[406]), .B1(n9766), 
        .B2(i_data_bus[502]), .ZN(n9785) );
  ND2D1BWP30P140LVT U14385 ( .A1(n9786), .A2(n9785), .ZN(N1225) );
  AOI22D1BWP30P140LVT U14386 ( .A1(n10633), .A2(i_data_bus[421]), .B1(n10632), 
        .B2(i_data_bus[453]), .ZN(n9788) );
  AOI22D1BWP30P140LVT U14387 ( .A1(n10634), .A2(i_data_bus[389]), .B1(n9766), 
        .B2(i_data_bus[485]), .ZN(n9787) );
  ND2D1BWP30P140LVT U14388 ( .A1(n9788), .A2(n9787), .ZN(N1208) );
  AOI22D1BWP30P140LVT U14389 ( .A1(n10633), .A2(i_data_bus[424]), .B1(n10632), 
        .B2(i_data_bus[456]), .ZN(n9790) );
  AOI22D1BWP30P140LVT U14390 ( .A1(n10634), .A2(i_data_bus[392]), .B1(n9766), 
        .B2(i_data_bus[488]), .ZN(n9789) );
  ND2D1BWP30P140LVT U14391 ( .A1(n9790), .A2(n9789), .ZN(N1211) );
  AOI22D1BWP30P140LVT U14392 ( .A1(n10634), .A2(i_data_bus[400]), .B1(n10632), 
        .B2(i_data_bus[464]), .ZN(n9792) );
  AOI22D1BWP30P140LVT U14393 ( .A1(n10633), .A2(i_data_bus[432]), .B1(n9766), 
        .B2(i_data_bus[496]), .ZN(n9791) );
  ND2D1BWP30P140LVT U14394 ( .A1(n9792), .A2(n9791), .ZN(N1219) );
  AOI22D1BWP30P140LVT U14395 ( .A1(n10634), .A2(i_data_bus[399]), .B1(n10632), 
        .B2(i_data_bus[463]), .ZN(n9794) );
  AOI22D1BWP30P140LVT U14396 ( .A1(n10633), .A2(i_data_bus[431]), .B1(n9766), 
        .B2(i_data_bus[495]), .ZN(n9793) );
  ND2D1BWP30P140LVT U14397 ( .A1(n9794), .A2(n9793), .ZN(N1218) );
  AOI22D1BWP30P140LVT U14398 ( .A1(n10634), .A2(i_data_bus[402]), .B1(n10632), 
        .B2(i_data_bus[466]), .ZN(n9796) );
  AOI22D1BWP30P140LVT U14399 ( .A1(n10633), .A2(i_data_bus[434]), .B1(n9766), 
        .B2(i_data_bus[498]), .ZN(n9795) );
  ND2D1BWP30P140LVT U14400 ( .A1(n9796), .A2(n9795), .ZN(N1221) );
  AOI22D1BWP30P140LVT U14401 ( .A1(n10634), .A2(i_data_bus[386]), .B1(n10632), 
        .B2(i_data_bus[450]), .ZN(n9798) );
  AOI22D1BWP30P140LVT U14402 ( .A1(n10633), .A2(i_data_bus[418]), .B1(n9766), 
        .B2(i_data_bus[482]), .ZN(n9797) );
  ND2D1BWP30P140LVT U14403 ( .A1(n9798), .A2(n9797), .ZN(N1205) );
  AOI22D1BWP30P140LVT U14404 ( .A1(n10634), .A2(i_data_bus[411]), .B1(n10632), 
        .B2(i_data_bus[475]), .ZN(n9800) );
  AOI22D1BWP30P140LVT U14405 ( .A1(n10633), .A2(i_data_bus[443]), .B1(n9766), 
        .B2(i_data_bus[507]), .ZN(n9799) );
  ND2D1BWP30P140LVT U14406 ( .A1(n9800), .A2(n9799), .ZN(N1230) );
  AOI22D1BWP30P140LVT U14407 ( .A1(n10621), .A2(i_data_bus[793]), .B1(n9749), 
        .B2(i_data_bus[889]), .ZN(n9802) );
  AOI22D1BWP30P140LVT U14408 ( .A1(n10623), .A2(i_data_bus[857]), .B1(n10622), 
        .B2(i_data_bus[825]), .ZN(n9801) );
  ND2D1BWP30P140LVT U14409 ( .A1(n9802), .A2(n9801), .ZN(N1888) );
  AOI22D1BWP30P140LVT U14410 ( .A1(n10621), .A2(i_data_bus[781]), .B1(n9749), 
        .B2(i_data_bus[877]), .ZN(n9804) );
  AOI22D1BWP30P140LVT U14411 ( .A1(n10623), .A2(i_data_bus[845]), .B1(n10622), 
        .B2(i_data_bus[813]), .ZN(n9803) );
  ND2D1BWP30P140LVT U14412 ( .A1(n9804), .A2(n9803), .ZN(N1876) );
  AOI22D1BWP30P140LVT U14413 ( .A1(i_data_bus[448]), .A2(n10632), .B1(
        i_data_bus[480]), .B2(n9766), .ZN(n9806) );
  AOI22D1BWP30P140LVT U14414 ( .A1(i_data_bus[384]), .A2(n10634), .B1(
        i_data_bus[416]), .B2(n10633), .ZN(n9805) );
  ND2D1BWP30P140LVT U14415 ( .A1(n9806), .A2(n9805), .ZN(N1203) );
  NR4D1BWP30P140LVT U14416 ( .A1(i_cmd[64]), .A2(n9811), .A3(n9807), .A4(n9809), .ZN(n10636) );
  NR4D1BWP30P140LVT U14417 ( .A1(i_cmd[80]), .A2(n9810), .A3(n9809), .A4(n9808), .ZN(n10635) );
  AOI22D1BWP30P140LVT U14418 ( .A1(i_data_bus[320]), .A2(n10636), .B1(
        i_data_bus[256]), .B2(n10635), .ZN(n9816) );
  INR4D1BWP30P140LVT U14419 ( .A1(i_cmd[88]), .B1(i_cmd[72]), .B2(n9812), .B3(
        n9814), .ZN(n10638) );
  INR4D1BWP30P140LVT U14420 ( .A1(i_cmd[72]), .B1(i_cmd[88]), .B2(n9814), .B3(
        n9813), .ZN(n10637) );
  AOI22D1BWP30P140LVT U14421 ( .A1(i_data_bus[352]), .A2(n10638), .B1(
        i_data_bus[288]), .B2(n10637), .ZN(n9815) );
  ND2D1BWP30P140LVT U14422 ( .A1(n9816), .A2(n9815), .ZN(N983) );
  AOI22D1BWP30P140LVT U14423 ( .A1(n10632), .A2(i_data_bus[449]), .B1(n9766), 
        .B2(i_data_bus[481]), .ZN(n9818) );
  AOI22D1BWP30P140LVT U14424 ( .A1(n10634), .A2(i_data_bus[385]), .B1(n10633), 
        .B2(i_data_bus[417]), .ZN(n9817) );
  ND2D1BWP30P140LVT U14425 ( .A1(n9818), .A2(n9817), .ZN(N1204) );
  AOI22D1BWP30P140LVT U14426 ( .A1(n10632), .A2(i_data_bus[462]), .B1(n9766), 
        .B2(i_data_bus[494]), .ZN(n9820) );
  AOI22D1BWP30P140LVT U14427 ( .A1(n10634), .A2(i_data_bus[398]), .B1(n10633), 
        .B2(i_data_bus[430]), .ZN(n9819) );
  ND2D1BWP30P140LVT U14428 ( .A1(n9820), .A2(n9819), .ZN(N1217) );
  AOI22D1BWP30P140LVT U14429 ( .A1(n10632), .A2(i_data_bus[465]), .B1(n9766), 
        .B2(i_data_bus[497]), .ZN(n9822) );
  AOI22D1BWP30P140LVT U14430 ( .A1(n10634), .A2(i_data_bus[401]), .B1(n10633), 
        .B2(i_data_bus[433]), .ZN(n9821) );
  ND2D1BWP30P140LVT U14431 ( .A1(n9822), .A2(n9821), .ZN(N1220) );
  AOI22D1BWP30P140LVT U14432 ( .A1(n10632), .A2(i_data_bus[478]), .B1(n9766), 
        .B2(i_data_bus[510]), .ZN(n9824) );
  AOI22D1BWP30P140LVT U14433 ( .A1(n10634), .A2(i_data_bus[414]), .B1(n10633), 
        .B2(i_data_bus[446]), .ZN(n9823) );
  ND2D1BWP30P140LVT U14434 ( .A1(n9824), .A2(n9823), .ZN(N1233) );
  AOI22D1BWP30P140LVT U14435 ( .A1(n10632), .A2(i_data_bus[459]), .B1(n9766), 
        .B2(i_data_bus[491]), .ZN(n9826) );
  AOI22D1BWP30P140LVT U14436 ( .A1(n10634), .A2(i_data_bus[395]), .B1(n10633), 
        .B2(i_data_bus[427]), .ZN(n9825) );
  ND2D1BWP30P140LVT U14437 ( .A1(n9826), .A2(n9825), .ZN(N1214) );
  AOI22D1BWP30P140LVT U14438 ( .A1(n10632), .A2(i_data_bus[461]), .B1(n9766), 
        .B2(i_data_bus[493]), .ZN(n9828) );
  AOI22D1BWP30P140LVT U14439 ( .A1(n10634), .A2(i_data_bus[397]), .B1(n10633), 
        .B2(i_data_bus[429]), .ZN(n9827) );
  ND2D1BWP30P140LVT U14440 ( .A1(n9828), .A2(n9827), .ZN(N1216) );
  AOI22D1BWP30P140LVT U14441 ( .A1(n10632), .A2(i_data_bus[469]), .B1(n9766), 
        .B2(i_data_bus[501]), .ZN(n9830) );
  AOI22D1BWP30P140LVT U14442 ( .A1(n10634), .A2(i_data_bus[405]), .B1(n10633), 
        .B2(i_data_bus[437]), .ZN(n9829) );
  ND2D1BWP30P140LVT U14443 ( .A1(n9830), .A2(n9829), .ZN(N1224) );
  AOI22D1BWP30P140LVT U14444 ( .A1(n10632), .A2(i_data_bus[468]), .B1(n9766), 
        .B2(i_data_bus[500]), .ZN(n9832) );
  AOI22D1BWP30P140LVT U14445 ( .A1(n10634), .A2(i_data_bus[404]), .B1(n10633), 
        .B2(i_data_bus[436]), .ZN(n9831) );
  ND2D1BWP30P140LVT U14446 ( .A1(n9832), .A2(n9831), .ZN(N1223) );
  INR4D1BWP30P140LVT U14447 ( .A1(i_cmd[136]), .B1(i_cmd[152]), .B2(n9836), 
        .B3(n9833), .ZN(n10629) );
  NR4D1BWP30P140LVT U14448 ( .A1(i_cmd[128]), .A2(n9835), .A3(n9838), .A4(
        n9834), .ZN(n10628) );
  AOI22D1BWP30P140LVT U14449 ( .A1(i_data_bus[544]), .A2(n10629), .B1(
        i_data_bus[576]), .B2(n10628), .ZN(n9842) );
  INR4D1BWP30P140LVT U14450 ( .A1(i_cmd[152]), .B1(i_cmd[136]), .B2(n9837), 
        .B3(n9836), .ZN(n10631) );
  NR4D1BWP30P140LVT U14451 ( .A1(i_cmd[144]), .A2(n9840), .A3(n9839), .A4(
        n9838), .ZN(n10630) );
  AOI22D1BWP30P140LVT U14452 ( .A1(i_data_bus[608]), .A2(n10631), .B1(
        i_data_bus[512]), .B2(n10630), .ZN(n9841) );
  ND2D1BWP30P140LVT U14453 ( .A1(n9842), .A2(n9841), .ZN(N1423) );
  INR4D1BWP30P140LVT U14454 ( .A1(i_cmd[160]), .B1(i_cmd[176]), .B2(n9849), 
        .B3(n9843), .ZN(n10625) );
  NR4D1BWP30P140LVT U14455 ( .A1(i_cmd[168]), .A2(n9848), .A3(n9845), .A4(
        n9844), .ZN(n10624) );
  AOI22D1BWP30P140LVT U14456 ( .A1(i_data_bus[640]), .A2(n10625), .B1(
        i_data_bus[736]), .B2(n10624), .ZN(n9852) );
  NR4D1BWP30P140LVT U14457 ( .A1(i_cmd[184]), .A2(n9848), .A3(n9847), .A4(
        n9846), .ZN(n10627) );
  INR4D1BWP30P140LVT U14458 ( .A1(i_cmd[176]), .B1(i_cmd[160]), .B2(n9850), 
        .B3(n9849), .ZN(n10626) );
  AOI22D1BWP30P140LVT U14459 ( .A1(i_data_bus[672]), .A2(n10627), .B1(
        i_data_bus[704]), .B2(n10626), .ZN(n9851) );
  ND2D1BWP30P140LVT U14460 ( .A1(n9852), .A2(n9851), .ZN(N1643) );
  INR4D1BWP30P140LVT U14461 ( .A1(i_cmd[40]), .B1(i_cmd[56]), .B2(n9859), .B3(
        n9853), .ZN(n10640) );
  NR4D1BWP30P140LVT U14462 ( .A1(i_cmd[32]), .A2(n9855), .A3(n9858), .A4(n9854), .ZN(n10639) );
  AOI22D1BWP30P140LVT U14463 ( .A1(i_data_bus[160]), .A2(n10640), .B1(
        i_data_bus[192]), .B2(n10639), .ZN(n9862) );
  NR4D1BWP30P140LVT U14464 ( .A1(i_cmd[48]), .A2(n9858), .A3(n9857), .A4(n9856), .ZN(n10642) );
  INR4D1BWP30P140LVT U14465 ( .A1(i_cmd[56]), .B1(i_cmd[40]), .B2(n9860), .B3(
        n9859), .ZN(n10641) );
  AOI22D1BWP30P140LVT U14466 ( .A1(i_data_bus[128]), .A2(n10642), .B1(
        i_data_bus[224]), .B2(n10641), .ZN(n9861) );
  ND2D1BWP30P140LVT U14467 ( .A1(n9862), .A2(n9861), .ZN(N763) );
  AOI22D1BWP30P140LVT U14468 ( .A1(n10622), .A2(i_data_bus[808]), .B1(n10621), 
        .B2(i_data_bus[776]), .ZN(n9864) );
  AOI22D1BWP30P140LVT U14469 ( .A1(n10623), .A2(i_data_bus[840]), .B1(n9749), 
        .B2(i_data_bus[872]), .ZN(n9863) );
  ND2D1BWP30P140LVT U14470 ( .A1(n9864), .A2(n9863), .ZN(N1871) );
  AOI22D1BWP30P140LVT U14471 ( .A1(n10622), .A2(i_data_bus[830]), .B1(n10621), 
        .B2(i_data_bus[798]), .ZN(n9866) );
  AOI22D1BWP30P140LVT U14472 ( .A1(n10623), .A2(i_data_bus[862]), .B1(n9749), 
        .B2(i_data_bus[894]), .ZN(n9865) );
  ND2D1BWP30P140LVT U14473 ( .A1(n9866), .A2(n9865), .ZN(N1893) );
  AOI22D1BWP30P140LVT U14474 ( .A1(n10622), .A2(i_data_bus[831]), .B1(n10621), 
        .B2(i_data_bus[799]), .ZN(n9868) );
  AOI22D1BWP30P140LVT U14475 ( .A1(n10623), .A2(i_data_bus[863]), .B1(n9749), 
        .B2(i_data_bus[895]), .ZN(n9867) );
  ND2D1BWP30P140LVT U14476 ( .A1(n9868), .A2(n9867), .ZN(N1894) );
  AOI22D1BWP30P140LVT U14477 ( .A1(n10622), .A2(i_data_bus[824]), .B1(n10621), 
        .B2(i_data_bus[792]), .ZN(n9870) );
  AOI22D1BWP30P140LVT U14478 ( .A1(n10623), .A2(i_data_bus[856]), .B1(n9749), 
        .B2(i_data_bus[888]), .ZN(n9869) );
  ND2D1BWP30P140LVT U14479 ( .A1(n9870), .A2(n9869), .ZN(N1887) );
  AOI22D1BWP30P140LVT U14480 ( .A1(n10622), .A2(i_data_bus[802]), .B1(n10621), 
        .B2(i_data_bus[770]), .ZN(n9872) );
  AOI22D1BWP30P140LVT U14481 ( .A1(n10623), .A2(i_data_bus[834]), .B1(n9749), 
        .B2(i_data_bus[866]), .ZN(n9871) );
  ND2D1BWP30P140LVT U14482 ( .A1(n9872), .A2(n9871), .ZN(N1865) );
  AOI22D1BWP30P140LVT U14483 ( .A1(n10622), .A2(i_data_bus[823]), .B1(n10621), 
        .B2(i_data_bus[791]), .ZN(n9874) );
  AOI22D1BWP30P140LVT U14484 ( .A1(n10623), .A2(i_data_bus[855]), .B1(n9749), 
        .B2(i_data_bus[887]), .ZN(n9873) );
  ND2D1BWP30P140LVT U14485 ( .A1(n9874), .A2(n9873), .ZN(N1886) );
  AOI22D1BWP30P140LVT U14486 ( .A1(n10622), .A2(i_data_bus[804]), .B1(n10621), 
        .B2(i_data_bus[772]), .ZN(n9876) );
  AOI22D1BWP30P140LVT U14487 ( .A1(n10623), .A2(i_data_bus[836]), .B1(n9749), 
        .B2(i_data_bus[868]), .ZN(n9875) );
  ND2D1BWP30P140LVT U14488 ( .A1(n9876), .A2(n9875), .ZN(N1867) );
  AOI22D1BWP30P140LVT U14489 ( .A1(n10622), .A2(i_data_bus[817]), .B1(n10621), 
        .B2(i_data_bus[785]), .ZN(n9878) );
  AOI22D1BWP30P140LVT U14490 ( .A1(n10623), .A2(i_data_bus[849]), .B1(n9749), 
        .B2(i_data_bus[881]), .ZN(n9877) );
  ND2D1BWP30P140LVT U14491 ( .A1(n9878), .A2(n9877), .ZN(N1880) );
  AOI22D1BWP30P140LVT U14492 ( .A1(n10622), .A2(i_data_bus[818]), .B1(n10621), 
        .B2(i_data_bus[786]), .ZN(n9880) );
  AOI22D1BWP30P140LVT U14493 ( .A1(n10623), .A2(i_data_bus[850]), .B1(n9749), 
        .B2(i_data_bus[882]), .ZN(n9879) );
  ND2D1BWP30P140LVT U14494 ( .A1(n9880), .A2(n9879), .ZN(N1881) );
  AOI22D1BWP30P140LVT U14495 ( .A1(n10623), .A2(i_data_bus[859]), .B1(n10621), 
        .B2(i_data_bus[795]), .ZN(n9882) );
  AOI22D1BWP30P140LVT U14496 ( .A1(n10622), .A2(i_data_bus[827]), .B1(n9749), 
        .B2(i_data_bus[891]), .ZN(n9881) );
  ND2D1BWP30P140LVT U14497 ( .A1(n9882), .A2(n9881), .ZN(N1890) );
  AOI22D1BWP30P140LVT U14498 ( .A1(n10623), .A2(i_data_bus[861]), .B1(n10621), 
        .B2(i_data_bus[797]), .ZN(n9884) );
  AOI22D1BWP30P140LVT U14499 ( .A1(n10622), .A2(i_data_bus[829]), .B1(n9749), 
        .B2(i_data_bus[893]), .ZN(n9883) );
  ND2D1BWP30P140LVT U14500 ( .A1(n9884), .A2(n9883), .ZN(N1892) );
  AOI22D1BWP30P140LVT U14501 ( .A1(n10623), .A2(i_data_bus[838]), .B1(n10621), 
        .B2(i_data_bus[774]), .ZN(n9886) );
  AOI22D1BWP30P140LVT U14502 ( .A1(n10622), .A2(i_data_bus[806]), .B1(n9749), 
        .B2(i_data_bus[870]), .ZN(n9885) );
  ND2D1BWP30P140LVT U14503 ( .A1(n9886), .A2(n9885), .ZN(N1869) );
  AOI22D1BWP30P140LVT U14504 ( .A1(n10623), .A2(i_data_bus[852]), .B1(n10621), 
        .B2(i_data_bus[788]), .ZN(n9888) );
  AOI22D1BWP30P140LVT U14505 ( .A1(n10622), .A2(i_data_bus[820]), .B1(n9749), 
        .B2(i_data_bus[884]), .ZN(n9887) );
  ND2D1BWP30P140LVT U14506 ( .A1(n9888), .A2(n9887), .ZN(N1883) );
  AOI22D1BWP30P140LVT U14507 ( .A1(n10623), .A2(i_data_bus[833]), .B1(n10621), 
        .B2(i_data_bus[769]), .ZN(n9890) );
  AOI22D1BWP30P140LVT U14508 ( .A1(n10622), .A2(i_data_bus[801]), .B1(n9749), 
        .B2(i_data_bus[865]), .ZN(n9889) );
  ND2D1BWP30P140LVT U14509 ( .A1(n9890), .A2(n9889), .ZN(N1864) );
  AOI22D1BWP30P140LVT U14510 ( .A1(n10623), .A2(i_data_bus[854]), .B1(n10621), 
        .B2(i_data_bus[790]), .ZN(n9892) );
  AOI22D1BWP30P140LVT U14511 ( .A1(n10622), .A2(i_data_bus[822]), .B1(n9749), 
        .B2(i_data_bus[886]), .ZN(n9891) );
  ND2D1BWP30P140LVT U14512 ( .A1(n9892), .A2(n9891), .ZN(N1885) );
  AOI22D1BWP30P140LVT U14513 ( .A1(n10623), .A2(i_data_bus[846]), .B1(n10621), 
        .B2(i_data_bus[782]), .ZN(n9894) );
  AOI22D1BWP30P140LVT U14514 ( .A1(n10622), .A2(i_data_bus[814]), .B1(n9749), 
        .B2(i_data_bus[878]), .ZN(n9893) );
  ND2D1BWP30P140LVT U14515 ( .A1(n9894), .A2(n9893), .ZN(N1877) );
  AOI22D1BWP30P140LVT U14516 ( .A1(n10623), .A2(i_data_bus[839]), .B1(n10621), 
        .B2(i_data_bus[775]), .ZN(n9896) );
  AOI22D1BWP30P140LVT U14517 ( .A1(n10622), .A2(i_data_bus[807]), .B1(n9749), 
        .B2(i_data_bus[871]), .ZN(n9895) );
  ND2D1BWP30P140LVT U14518 ( .A1(n9896), .A2(n9895), .ZN(N1870) );
  AOI22D1BWP30P140LVT U14519 ( .A1(n10623), .A2(i_data_bus[837]), .B1(n10621), 
        .B2(i_data_bus[773]), .ZN(n9898) );
  AOI22D1BWP30P140LVT U14520 ( .A1(n10622), .A2(i_data_bus[805]), .B1(n9749), 
        .B2(i_data_bus[869]), .ZN(n9897) );
  ND2D1BWP30P140LVT U14521 ( .A1(n9898), .A2(n9897), .ZN(N1868) );
  AOI22D1BWP30P140LVT U14522 ( .A1(n10636), .A2(i_data_bus[323]), .B1(n10635), 
        .B2(i_data_bus[259]), .ZN(n9900) );
  AOI22D1BWP30P140LVT U14523 ( .A1(n10638), .A2(i_data_bus[355]), .B1(n10637), 
        .B2(i_data_bus[291]), .ZN(n9899) );
  ND2D1BWP30P140LVT U14524 ( .A1(n9900), .A2(n9899), .ZN(N986) );
  AOI22D1BWP30P140LVT U14525 ( .A1(n10636), .A2(i_data_bus[340]), .B1(n10635), 
        .B2(i_data_bus[276]), .ZN(n9902) );
  AOI22D1BWP30P140LVT U14526 ( .A1(n10638), .A2(i_data_bus[372]), .B1(n10637), 
        .B2(i_data_bus[308]), .ZN(n9901) );
  ND2D1BWP30P140LVT U14527 ( .A1(n9902), .A2(n9901), .ZN(N1003) );
  AOI22D1BWP30P140LVT U14528 ( .A1(n10629), .A2(i_data_bus[553]), .B1(n10628), 
        .B2(i_data_bus[585]), .ZN(n9904) );
  AOI22D1BWP30P140LVT U14529 ( .A1(n10631), .A2(i_data_bus[617]), .B1(n10630), 
        .B2(i_data_bus[521]), .ZN(n9903) );
  ND2D1BWP30P140LVT U14530 ( .A1(n9904), .A2(n9903), .ZN(N1432) );
  AOI22D1BWP30P140LVT U14531 ( .A1(n10629), .A2(i_data_bus[548]), .B1(n10628), 
        .B2(i_data_bus[580]), .ZN(n9906) );
  AOI22D1BWP30P140LVT U14532 ( .A1(n10631), .A2(i_data_bus[612]), .B1(n10630), 
        .B2(i_data_bus[516]), .ZN(n9905) );
  ND2D1BWP30P140LVT U14533 ( .A1(n9906), .A2(n9905), .ZN(N1427) );
  AOI22D1BWP30P140LVT U14534 ( .A1(n10629), .A2(i_data_bus[563]), .B1(n10628), 
        .B2(i_data_bus[595]), .ZN(n9908) );
  AOI22D1BWP30P140LVT U14535 ( .A1(n10631), .A2(i_data_bus[627]), .B1(n10630), 
        .B2(i_data_bus[531]), .ZN(n9907) );
  ND2D1BWP30P140LVT U14536 ( .A1(n9908), .A2(n9907), .ZN(N1442) );
  AOI22D1BWP30P140LVT U14537 ( .A1(n10629), .A2(i_data_bus[574]), .B1(n10628), 
        .B2(i_data_bus[606]), .ZN(n9910) );
  AOI22D1BWP30P140LVT U14538 ( .A1(n10631), .A2(i_data_bus[638]), .B1(n10630), 
        .B2(i_data_bus[542]), .ZN(n9909) );
  ND2D1BWP30P140LVT U14539 ( .A1(n9910), .A2(n9909), .ZN(N1453) );
  AOI22D1BWP30P140LVT U14540 ( .A1(n10629), .A2(i_data_bus[551]), .B1(n10628), 
        .B2(i_data_bus[583]), .ZN(n9912) );
  AOI22D1BWP30P140LVT U14541 ( .A1(n10631), .A2(i_data_bus[615]), .B1(n10630), 
        .B2(i_data_bus[519]), .ZN(n9911) );
  ND2D1BWP30P140LVT U14542 ( .A1(n9912), .A2(n9911), .ZN(N1430) );
  AOI22D1BWP30P140LVT U14543 ( .A1(n10630), .A2(i_data_bus[539]), .B1(n10628), 
        .B2(i_data_bus[603]), .ZN(n9914) );
  AOI22D1BWP30P140LVT U14544 ( .A1(n10631), .A2(i_data_bus[635]), .B1(n10629), 
        .B2(i_data_bus[571]), .ZN(n9913) );
  ND2D1BWP30P140LVT U14545 ( .A1(n9914), .A2(n9913), .ZN(N1450) );
  AOI22D1BWP30P140LVT U14546 ( .A1(n10630), .A2(i_data_bus[518]), .B1(n10628), 
        .B2(i_data_bus[582]), .ZN(n9916) );
  AOI22D1BWP30P140LVT U14547 ( .A1(n10631), .A2(i_data_bus[614]), .B1(n10629), 
        .B2(i_data_bus[550]), .ZN(n9915) );
  ND2D1BWP30P140LVT U14548 ( .A1(n9916), .A2(n9915), .ZN(N1429) );
  AOI22D1BWP30P140LVT U14549 ( .A1(n10631), .A2(i_data_bus[613]), .B1(n10628), 
        .B2(i_data_bus[581]), .ZN(n9918) );
  AOI22D1BWP30P140LVT U14550 ( .A1(n10630), .A2(i_data_bus[517]), .B1(n10629), 
        .B2(i_data_bus[549]), .ZN(n9917) );
  ND2D1BWP30P140LVT U14551 ( .A1(n9918), .A2(n9917), .ZN(N1428) );
  AOI22D1BWP30P140LVT U14552 ( .A1(n10631), .A2(i_data_bus[622]), .B1(n10628), 
        .B2(i_data_bus[590]), .ZN(n9920) );
  AOI22D1BWP30P140LVT U14553 ( .A1(n10630), .A2(i_data_bus[526]), .B1(n10629), 
        .B2(i_data_bus[558]), .ZN(n9919) );
  ND2D1BWP30P140LVT U14554 ( .A1(n9920), .A2(n9919), .ZN(N1437) );
  AOI22D1BWP30P140LVT U14555 ( .A1(n10630), .A2(i_data_bus[520]), .B1(n10628), 
        .B2(i_data_bus[584]), .ZN(n9922) );
  AOI22D1BWP30P140LVT U14556 ( .A1(n10631), .A2(i_data_bus[616]), .B1(n10629), 
        .B2(i_data_bus[552]), .ZN(n9921) );
  ND2D1BWP30P140LVT U14557 ( .A1(n9922), .A2(n9921), .ZN(N1431) );
  AOI22D1BWP30P140LVT U14558 ( .A1(n10630), .A2(i_data_bus[525]), .B1(n10628), 
        .B2(i_data_bus[589]), .ZN(n9924) );
  AOI22D1BWP30P140LVT U14559 ( .A1(n10631), .A2(i_data_bus[621]), .B1(n10629), 
        .B2(i_data_bus[557]), .ZN(n9923) );
  ND2D1BWP30P140LVT U14560 ( .A1(n9924), .A2(n9923), .ZN(N1436) );
  AOI22D1BWP30P140LVT U14561 ( .A1(n10630), .A2(i_data_bus[528]), .B1(n10628), 
        .B2(i_data_bus[592]), .ZN(n9926) );
  AOI22D1BWP30P140LVT U14562 ( .A1(n10631), .A2(i_data_bus[624]), .B1(n10629), 
        .B2(i_data_bus[560]), .ZN(n9925) );
  ND2D1BWP30P140LVT U14563 ( .A1(n9926), .A2(n9925), .ZN(N1439) );
  AOI22D1BWP30P140LVT U14564 ( .A1(n10631), .A2(i_data_bus[620]), .B1(n10628), 
        .B2(i_data_bus[588]), .ZN(n9928) );
  AOI22D1BWP30P140LVT U14565 ( .A1(n10630), .A2(i_data_bus[524]), .B1(n10629), 
        .B2(i_data_bus[556]), .ZN(n9927) );
  ND2D1BWP30P140LVT U14566 ( .A1(n9928), .A2(n9927), .ZN(N1435) );
  AOI22D1BWP30P140LVT U14567 ( .A1(n10630), .A2(i_data_bus[534]), .B1(n10628), 
        .B2(i_data_bus[598]), .ZN(n9930) );
  AOI22D1BWP30P140LVT U14568 ( .A1(n10631), .A2(i_data_bus[630]), .B1(n10629), 
        .B2(i_data_bus[566]), .ZN(n9929) );
  ND2D1BWP30P140LVT U14569 ( .A1(n9930), .A2(n9929), .ZN(N1445) );
  AOI22D1BWP30P140LVT U14570 ( .A1(n10634), .A2(i_data_bus[407]), .B1(n9766), 
        .B2(i_data_bus[503]), .ZN(n9932) );
  AOI22D1BWP30P140LVT U14571 ( .A1(n10633), .A2(i_data_bus[439]), .B1(n10632), 
        .B2(i_data_bus[471]), .ZN(n9931) );
  ND2D1BWP30P140LVT U14572 ( .A1(n9932), .A2(n9931), .ZN(N1226) );
  AOI22D1BWP30P140LVT U14573 ( .A1(n10633), .A2(i_data_bus[441]), .B1(n9766), 
        .B2(i_data_bus[505]), .ZN(n9934) );
  AOI22D1BWP30P140LVT U14574 ( .A1(n10634), .A2(i_data_bus[409]), .B1(n10632), 
        .B2(i_data_bus[473]), .ZN(n9933) );
  ND2D1BWP30P140LVT U14575 ( .A1(n9934), .A2(n9933), .ZN(N1228) );
  AOI22D1BWP30P140LVT U14576 ( .A1(n10633), .A2(i_data_bus[447]), .B1(n9766), 
        .B2(i_data_bus[511]), .ZN(n9936) );
  AOI22D1BWP30P140LVT U14577 ( .A1(n10634), .A2(i_data_bus[415]), .B1(n10632), 
        .B2(i_data_bus[479]), .ZN(n9935) );
  ND2D1BWP30P140LVT U14578 ( .A1(n9936), .A2(n9935), .ZN(N1234) );
  AOI22D1BWP30P140LVT U14579 ( .A1(n10633), .A2(i_data_bus[420]), .B1(n9766), 
        .B2(i_data_bus[484]), .ZN(n9938) );
  AOI22D1BWP30P140LVT U14580 ( .A1(n10634), .A2(i_data_bus[388]), .B1(n10632), 
        .B2(i_data_bus[452]), .ZN(n9937) );
  ND2D1BWP30P140LVT U14581 ( .A1(n9938), .A2(n9937), .ZN(N1207) );
  AOI22D1BWP30P140LVT U14582 ( .A1(n10633), .A2(i_data_bus[440]), .B1(n9766), 
        .B2(i_data_bus[504]), .ZN(n9940) );
  AOI22D1BWP30P140LVT U14583 ( .A1(n10634), .A2(i_data_bus[408]), .B1(n10632), 
        .B2(i_data_bus[472]), .ZN(n9939) );
  ND2D1BWP30P140LVT U14584 ( .A1(n9940), .A2(n9939), .ZN(N1227) );
  AOI22D1BWP30P140LVT U14585 ( .A1(n10634), .A2(i_data_bus[390]), .B1(n9766), 
        .B2(i_data_bus[486]), .ZN(n9942) );
  AOI22D1BWP30P140LVT U14586 ( .A1(n10633), .A2(i_data_bus[422]), .B1(n10632), 
        .B2(i_data_bus[454]), .ZN(n9941) );
  ND2D1BWP30P140LVT U14587 ( .A1(n9942), .A2(n9941), .ZN(N1209) );
  AOI22D1BWP30P140LVT U14588 ( .A1(n10634), .A2(i_data_bus[412]), .B1(n9766), 
        .B2(i_data_bus[508]), .ZN(n9944) );
  AOI22D1BWP30P140LVT U14589 ( .A1(n10633), .A2(i_data_bus[444]), .B1(n10632), 
        .B2(i_data_bus[476]), .ZN(n9943) );
  ND2D1BWP30P140LVT U14590 ( .A1(n9944), .A2(n9943), .ZN(N1231) );
  AOI22D1BWP30P140LVT U14591 ( .A1(n10625), .A2(i_data_bus[654]), .B1(n10624), 
        .B2(i_data_bus[750]), .ZN(n9946) );
  AOI22D1BWP30P140LVT U14592 ( .A1(n10627), .A2(i_data_bus[686]), .B1(n10626), 
        .B2(i_data_bus[718]), .ZN(n9945) );
  ND2D1BWP30P140LVT U14593 ( .A1(n9946), .A2(n9945), .ZN(N1657) );
  AOI22D1BWP30P140LVT U14594 ( .A1(n10625), .A2(i_data_bus[649]), .B1(n10624), 
        .B2(i_data_bus[745]), .ZN(n9948) );
  AOI22D1BWP30P140LVT U14595 ( .A1(n10627), .A2(i_data_bus[681]), .B1(n10626), 
        .B2(i_data_bus[713]), .ZN(n9947) );
  ND2D1BWP30P140LVT U14596 ( .A1(n9948), .A2(n9947), .ZN(N1652) );
  AOI22D1BWP30P140LVT U14597 ( .A1(n10625), .A2(i_data_bus[664]), .B1(n10624), 
        .B2(i_data_bus[760]), .ZN(n9950) );
  AOI22D1BWP30P140LVT U14598 ( .A1(n10627), .A2(i_data_bus[696]), .B1(n10626), 
        .B2(i_data_bus[728]), .ZN(n9949) );
  ND2D1BWP30P140LVT U14599 ( .A1(n9950), .A2(n9949), .ZN(N1667) );
  AOI22D1BWP30P140LVT U14600 ( .A1(n10625), .A2(i_data_bus[671]), .B1(n10624), 
        .B2(i_data_bus[767]), .ZN(n9952) );
  AOI22D1BWP30P140LVT U14601 ( .A1(n10627), .A2(i_data_bus[703]), .B1(n10626), 
        .B2(i_data_bus[735]), .ZN(n9951) );
  ND2D1BWP30P140LVT U14602 ( .A1(n9952), .A2(n9951), .ZN(N1674) );
  AOI22D1BWP30P140LVT U14603 ( .A1(n10625), .A2(i_data_bus[647]), .B1(n10624), 
        .B2(i_data_bus[743]), .ZN(n9954) );
  AOI22D1BWP30P140LVT U14604 ( .A1(n10627), .A2(i_data_bus[679]), .B1(n10626), 
        .B2(i_data_bus[711]), .ZN(n9953) );
  ND2D1BWP30P140LVT U14605 ( .A1(n9954), .A2(n9953), .ZN(N1650) );
  AOI22D1BWP30P140LVT U14606 ( .A1(n10625), .A2(i_data_bus[655]), .B1(n10624), 
        .B2(i_data_bus[751]), .ZN(n9956) );
  AOI22D1BWP30P140LVT U14607 ( .A1(n10627), .A2(i_data_bus[687]), .B1(n10626), 
        .B2(i_data_bus[719]), .ZN(n9955) );
  ND2D1BWP30P140LVT U14608 ( .A1(n9956), .A2(n9955), .ZN(N1658) );
  AOI22D1BWP30P140LVT U14609 ( .A1(n10625), .A2(i_data_bus[645]), .B1(n10624), 
        .B2(i_data_bus[741]), .ZN(n9958) );
  AOI22D1BWP30P140LVT U14610 ( .A1(n10627), .A2(i_data_bus[677]), .B1(n10626), 
        .B2(i_data_bus[709]), .ZN(n9957) );
  ND2D1BWP30P140LVT U14611 ( .A1(n9958), .A2(n9957), .ZN(N1648) );
  AOI22D1BWP30P140LVT U14612 ( .A1(n10625), .A2(i_data_bus[652]), .B1(n10624), 
        .B2(i_data_bus[748]), .ZN(n9960) );
  AOI22D1BWP30P140LVT U14613 ( .A1(n10627), .A2(i_data_bus[684]), .B1(n10626), 
        .B2(i_data_bus[716]), .ZN(n9959) );
  ND2D1BWP30P140LVT U14614 ( .A1(n9960), .A2(n9959), .ZN(N1655) );
  AOI22D1BWP30P140LVT U14615 ( .A1(n10626), .A2(i_data_bus[727]), .B1(n10624), 
        .B2(i_data_bus[759]), .ZN(n9962) );
  AOI22D1BWP30P140LVT U14616 ( .A1(n10627), .A2(i_data_bus[695]), .B1(n10625), 
        .B2(i_data_bus[663]), .ZN(n9961) );
  ND2D1BWP30P140LVT U14617 ( .A1(n9962), .A2(n9961), .ZN(N1666) );
  AOI22D1BWP30P140LVT U14618 ( .A1(n10627), .A2(i_data_bus[701]), .B1(n10624), 
        .B2(i_data_bus[765]), .ZN(n9964) );
  AOI22D1BWP30P140LVT U14619 ( .A1(n10626), .A2(i_data_bus[733]), .B1(n10625), 
        .B2(i_data_bus[669]), .ZN(n9963) );
  ND2D1BWP30P140LVT U14620 ( .A1(n9964), .A2(n9963), .ZN(N1672) );
  AOI22D1BWP30P140LVT U14621 ( .A1(n10626), .A2(i_data_bus[730]), .B1(n10624), 
        .B2(i_data_bus[762]), .ZN(n9966) );
  AOI22D1BWP30P140LVT U14622 ( .A1(n10627), .A2(i_data_bus[698]), .B1(n10625), 
        .B2(i_data_bus[666]), .ZN(n9965) );
  ND2D1BWP30P140LVT U14623 ( .A1(n9966), .A2(n9965), .ZN(N1669) );
  AOI22D1BWP30P140LVT U14624 ( .A1(n10626), .A2(i_data_bus[724]), .B1(n10624), 
        .B2(i_data_bus[756]), .ZN(n9968) );
  AOI22D1BWP30P140LVT U14625 ( .A1(n10627), .A2(i_data_bus[692]), .B1(n10625), 
        .B2(i_data_bus[660]), .ZN(n9967) );
  ND2D1BWP30P140LVT U14626 ( .A1(n9968), .A2(n9967), .ZN(N1663) );
  AOI22D1BWP30P140LVT U14627 ( .A1(n10626), .A2(i_data_bus[705]), .B1(n10624), 
        .B2(i_data_bus[737]), .ZN(n9970) );
  AOI22D1BWP30P140LVT U14628 ( .A1(n10627), .A2(i_data_bus[673]), .B1(n10625), 
        .B2(i_data_bus[641]), .ZN(n9969) );
  ND2D1BWP30P140LVT U14629 ( .A1(n9970), .A2(n9969), .ZN(N1644) );
  AOI22D1BWP30P140LVT U14630 ( .A1(n10627), .A2(i_data_bus[678]), .B1(n10624), 
        .B2(i_data_bus[742]), .ZN(n9972) );
  AOI22D1BWP30P140LVT U14631 ( .A1(n10626), .A2(i_data_bus[710]), .B1(n10625), 
        .B2(i_data_bus[646]), .ZN(n9971) );
  ND2D1BWP30P140LVT U14632 ( .A1(n9972), .A2(n9971), .ZN(N1649) );
  AOI22D1BWP30P140LVT U14633 ( .A1(n10627), .A2(i_data_bus[675]), .B1(n10624), 
        .B2(i_data_bus[739]), .ZN(n9974) );
  AOI22D1BWP30P140LVT U14634 ( .A1(n10626), .A2(i_data_bus[707]), .B1(n10625), 
        .B2(i_data_bus[643]), .ZN(n9973) );
  ND2D1BWP30P140LVT U14635 ( .A1(n9974), .A2(n9973), .ZN(N1646) );
  AOI22D1BWP30P140LVT U14636 ( .A1(n10627), .A2(i_data_bus[683]), .B1(n10624), 
        .B2(i_data_bus[747]), .ZN(n9976) );
  AOI22D1BWP30P140LVT U14637 ( .A1(n10626), .A2(i_data_bus[715]), .B1(n10625), 
        .B2(i_data_bus[651]), .ZN(n9975) );
  ND2D1BWP30P140LVT U14638 ( .A1(n9976), .A2(n9975), .ZN(N1654) );
  AOI22D1BWP30P140LVT U14639 ( .A1(n10627), .A2(i_data_bus[690]), .B1(n10624), 
        .B2(i_data_bus[754]), .ZN(n9978) );
  AOI22D1BWP30P140LVT U14640 ( .A1(n10626), .A2(i_data_bus[722]), .B1(n10625), 
        .B2(i_data_bus[658]), .ZN(n9977) );
  ND2D1BWP30P140LVT U14641 ( .A1(n9978), .A2(n9977), .ZN(N1661) );
  AOI22D1BWP30P140LVT U14642 ( .A1(n10627), .A2(i_data_bus[674]), .B1(n10624), 
        .B2(i_data_bus[738]), .ZN(n9980) );
  AOI22D1BWP30P140LVT U14643 ( .A1(n10626), .A2(i_data_bus[706]), .B1(n10625), 
        .B2(i_data_bus[642]), .ZN(n9979) );
  ND2D1BWP30P140LVT U14644 ( .A1(n9980), .A2(n9979), .ZN(N1645) );
  AOI22D1BWP30P140LVT U14645 ( .A1(n10640), .A2(i_data_bus[181]), .B1(n10639), 
        .B2(i_data_bus[213]), .ZN(n9982) );
  AOI22D1BWP30P140LVT U14646 ( .A1(n10642), .A2(i_data_bus[149]), .B1(n10641), 
        .B2(i_data_bus[245]), .ZN(n9981) );
  ND2D1BWP30P140LVT U14647 ( .A1(n9982), .A2(n9981), .ZN(N784) );
  AOI22D1BWP30P140LVT U14648 ( .A1(n10640), .A2(i_data_bus[164]), .B1(n10639), 
        .B2(i_data_bus[196]), .ZN(n9984) );
  AOI22D1BWP30P140LVT U14649 ( .A1(n10642), .A2(i_data_bus[132]), .B1(n10641), 
        .B2(i_data_bus[228]), .ZN(n9983) );
  ND2D1BWP30P140LVT U14650 ( .A1(n9984), .A2(n9983), .ZN(N767) );
  AOI22D1BWP30P140LVT U14651 ( .A1(n10640), .A2(i_data_bus[188]), .B1(n10639), 
        .B2(i_data_bus[220]), .ZN(n9986) );
  AOI22D1BWP30P140LVT U14652 ( .A1(n10642), .A2(i_data_bus[156]), .B1(n10641), 
        .B2(i_data_bus[252]), .ZN(n9985) );
  ND2D1BWP30P140LVT U14653 ( .A1(n9986), .A2(n9985), .ZN(N791) );
  AOI22D1BWP30P140LVT U14654 ( .A1(n10641), .A2(i_data_bus[251]), .B1(n10639), 
        .B2(i_data_bus[219]), .ZN(n9988) );
  AOI22D1BWP30P140LVT U14655 ( .A1(n10642), .A2(i_data_bus[155]), .B1(n10640), 
        .B2(i_data_bus[187]), .ZN(n9987) );
  ND2D1BWP30P140LVT U14656 ( .A1(n9988), .A2(n9987), .ZN(N790) );
  AOI22D1BWP30P140LVT U14657 ( .A1(n10641), .A2(i_data_bus[250]), .B1(n10639), 
        .B2(i_data_bus[218]), .ZN(n9990) );
  AOI22D1BWP30P140LVT U14658 ( .A1(n10642), .A2(i_data_bus[154]), .B1(n10640), 
        .B2(i_data_bus[186]), .ZN(n9989) );
  ND2D1BWP30P140LVT U14659 ( .A1(n9990), .A2(n9989), .ZN(N789) );
  AOI22D1BWP30P140LVT U14660 ( .A1(n10641), .A2(i_data_bus[229]), .B1(n10639), 
        .B2(i_data_bus[197]), .ZN(n9992) );
  AOI22D1BWP30P140LVT U14661 ( .A1(n10642), .A2(i_data_bus[133]), .B1(n10640), 
        .B2(i_data_bus[165]), .ZN(n9991) );
  ND2D1BWP30P140LVT U14662 ( .A1(n9992), .A2(n9991), .ZN(N768) );
  AOI22D1BWP30P140LVT U14663 ( .A1(n10641), .A2(i_data_bus[243]), .B1(n10639), 
        .B2(i_data_bus[211]), .ZN(n9994) );
  AOI22D1BWP30P140LVT U14664 ( .A1(n10642), .A2(i_data_bus[147]), .B1(n10640), 
        .B2(i_data_bus[179]), .ZN(n9993) );
  ND2D1BWP30P140LVT U14665 ( .A1(n9994), .A2(n9993), .ZN(N782) );
  AOI22D1BWP30P140LVT U14666 ( .A1(n10641), .A2(i_data_bus[244]), .B1(n10639), 
        .B2(i_data_bus[212]), .ZN(n9996) );
  AOI22D1BWP30P140LVT U14667 ( .A1(n10642), .A2(i_data_bus[148]), .B1(n10640), 
        .B2(i_data_bus[180]), .ZN(n9995) );
  ND2D1BWP30P140LVT U14668 ( .A1(n9996), .A2(n9995), .ZN(N783) );
  AOI22D1BWP30P140LVT U14669 ( .A1(n10641), .A2(i_data_bus[247]), .B1(n10639), 
        .B2(i_data_bus[215]), .ZN(n9998) );
  AOI22D1BWP30P140LVT U14670 ( .A1(n10642), .A2(i_data_bus[151]), .B1(n10640), 
        .B2(i_data_bus[183]), .ZN(n9997) );
  ND2D1BWP30P140LVT U14671 ( .A1(n9998), .A2(n9997), .ZN(N786) );
  AOI22D1BWP30P140LVT U14672 ( .A1(n10642), .A2(i_data_bus[142]), .B1(n10639), 
        .B2(i_data_bus[206]), .ZN(n10000) );
  AOI22D1BWP30P140LVT U14673 ( .A1(n10641), .A2(i_data_bus[238]), .B1(n10640), 
        .B2(i_data_bus[174]), .ZN(n9999) );
  ND2D1BWP30P140LVT U14674 ( .A1(n10000), .A2(n9999), .ZN(N777) );
  AOI22D1BWP30P140LVT U14675 ( .A1(n10642), .A2(i_data_bus[153]), .B1(n10639), 
        .B2(i_data_bus[217]), .ZN(n10002) );
  AOI22D1BWP30P140LVT U14676 ( .A1(n10641), .A2(i_data_bus[249]), .B1(n10640), 
        .B2(i_data_bus[185]), .ZN(n10001) );
  ND2D1BWP30P140LVT U14677 ( .A1(n10002), .A2(n10001), .ZN(N788) );
  AOI22D1BWP30P140LVT U14678 ( .A1(n10642), .A2(i_data_bus[135]), .B1(n10639), 
        .B2(i_data_bus[199]), .ZN(n10004) );
  AOI22D1BWP30P140LVT U14679 ( .A1(n10641), .A2(i_data_bus[231]), .B1(n10640), 
        .B2(i_data_bus[167]), .ZN(n10003) );
  ND2D1BWP30P140LVT U14680 ( .A1(n10004), .A2(n10003), .ZN(N770) );
  AOI22D1BWP30P140LVT U14681 ( .A1(n10642), .A2(i_data_bus[131]), .B1(n10639), 
        .B2(i_data_bus[195]), .ZN(n10006) );
  AOI22D1BWP30P140LVT U14682 ( .A1(n10641), .A2(i_data_bus[227]), .B1(n10640), 
        .B2(i_data_bus[163]), .ZN(n10005) );
  ND2D1BWP30P140LVT U14683 ( .A1(n10006), .A2(n10005), .ZN(N766) );
  AOI22D1BWP30P140LVT U14684 ( .A1(n10641), .A2(i_data_bus[225]), .B1(n10639), 
        .B2(i_data_bus[193]), .ZN(n10008) );
  AOI22D1BWP30P140LVT U14685 ( .A1(n10642), .A2(i_data_bus[129]), .B1(n10640), 
        .B2(i_data_bus[161]), .ZN(n10007) );
  ND2D1BWP30P140LVT U14686 ( .A1(n10008), .A2(n10007), .ZN(N764) );
  AOI22D1BWP30P140LVT U14687 ( .A1(n10642), .A2(i_data_bus[138]), .B1(n10639), 
        .B2(i_data_bus[202]), .ZN(n10010) );
  AOI22D1BWP30P140LVT U14688 ( .A1(n10641), .A2(i_data_bus[234]), .B1(n10640), 
        .B2(i_data_bus[170]), .ZN(n10009) );
  ND2D1BWP30P140LVT U14689 ( .A1(n10010), .A2(n10009), .ZN(N773) );
  AOI22D1BWP30P140LVT U14690 ( .A1(n10641), .A2(i_data_bus[242]), .B1(n10639), 
        .B2(i_data_bus[210]), .ZN(n10012) );
  AOI22D1BWP30P140LVT U14691 ( .A1(n10642), .A2(i_data_bus[146]), .B1(n10640), 
        .B2(i_data_bus[178]), .ZN(n10011) );
  ND2D1BWP30P140LVT U14692 ( .A1(n10012), .A2(n10011), .ZN(N781) );
  NR4D1BWP30P140LVT U14693 ( .A1(i_cmd[16]), .A2(n10016), .A3(n10013), .A4(
        n10015), .ZN(n10644) );
  NR4D1BWP30P140LVT U14694 ( .A1(i_cmd[0]), .A2(n10017), .A3(n10015), .A4(
        n10014), .ZN(n10643) );
  AOI22D1BWP30P140LVT U14695 ( .A1(i_data_bus[0]), .A2(n10644), .B1(
        i_data_bus[64]), .B2(n10643), .ZN(n10022) );
  INR4D1BWP30P140LVT U14696 ( .A1(i_cmd[8]), .B1(i_cmd[24]), .B2(n10018), .B3(
        n10020), .ZN(n10646) );
  INR4D1BWP30P140LVT U14697 ( .A1(i_cmd[24]), .B1(i_cmd[8]), .B2(n10020), .B3(
        n10019), .ZN(n10645) );
  AOI22D1BWP30P140LVT U14698 ( .A1(i_data_bus[32]), .A2(n10646), .B1(
        i_data_bus[96]), .B2(n10645), .ZN(n10021) );
  ND2D1BWP30P140LVT U14699 ( .A1(n10022), .A2(n10021), .ZN(N543) );
  INR4D1BWP30P140LVT U14700 ( .A1(i_cmd[232]), .B1(i_cmd[248]), .B2(n10029), 
        .B3(n10023), .ZN(n10618) );
  NR4D1BWP30P140LVT U14701 ( .A1(i_cmd[224]), .A2(n10025), .A3(n10026), .A4(
        n10024), .ZN(n10617) );
  AOI22D1BWP30P140LVT U14702 ( .A1(i_data_bus[928]), .A2(n10618), .B1(
        i_data_bus[960]), .B2(n10617), .ZN(n10032) );
  NR4D1BWP30P140LVT U14703 ( .A1(i_cmd[240]), .A2(n10028), .A3(n10027), .A4(
        n10026), .ZN(n10620) );
  INR4D1BWP30P140LVT U14704 ( .A1(i_cmd[248]), .B1(i_cmd[232]), .B2(n10030), 
        .B3(n10029), .ZN(n10619) );
  AOI22D1BWP30P140LVT U14705 ( .A1(i_data_bus[896]), .A2(n10620), .B1(
        i_data_bus[992]), .B2(n10619), .ZN(n10031) );
  ND2D1BWP30P140LVT U14706 ( .A1(n10032), .A2(n10031), .ZN(N2083) );
  AOI22D1BWP30P140LVT U14707 ( .A1(n10637), .A2(i_data_bus[293]), .B1(n10635), 
        .B2(i_data_bus[261]), .ZN(n10034) );
  AOI22D1BWP30P140LVT U14708 ( .A1(n10638), .A2(i_data_bus[357]), .B1(n10636), 
        .B2(i_data_bus[325]), .ZN(n10033) );
  ND2D1BWP30P140LVT U14709 ( .A1(n10034), .A2(n10033), .ZN(N988) );
  AOI22D1BWP30P140LVT U14710 ( .A1(n10637), .A2(i_data_bus[304]), .B1(n10635), 
        .B2(i_data_bus[272]), .ZN(n10036) );
  AOI22D1BWP30P140LVT U14711 ( .A1(n10638), .A2(i_data_bus[368]), .B1(n10636), 
        .B2(i_data_bus[336]), .ZN(n10035) );
  ND2D1BWP30P140LVT U14712 ( .A1(n10036), .A2(n10035), .ZN(N999) );
  AOI22D1BWP30P140LVT U14713 ( .A1(n10637), .A2(i_data_bus[318]), .B1(n10635), 
        .B2(i_data_bus[286]), .ZN(n10038) );
  AOI22D1BWP30P140LVT U14714 ( .A1(n10638), .A2(i_data_bus[382]), .B1(n10636), 
        .B2(i_data_bus[350]), .ZN(n10037) );
  ND2D1BWP30P140LVT U14715 ( .A1(n10038), .A2(n10037), .ZN(N1013) );
  AOI22D1BWP30P140LVT U14716 ( .A1(n10637), .A2(i_data_bus[306]), .B1(n10635), 
        .B2(i_data_bus[274]), .ZN(n10040) );
  AOI22D1BWP30P140LVT U14717 ( .A1(n10638), .A2(i_data_bus[370]), .B1(n10636), 
        .B2(i_data_bus[338]), .ZN(n10039) );
  ND2D1BWP30P140LVT U14718 ( .A1(n10040), .A2(n10039), .ZN(N1001) );
  AOI22D1BWP30P140LVT U14719 ( .A1(n10638), .A2(i_data_bus[373]), .B1(n10635), 
        .B2(i_data_bus[277]), .ZN(n10042) );
  AOI22D1BWP30P140LVT U14720 ( .A1(n10637), .A2(i_data_bus[309]), .B1(n10636), 
        .B2(i_data_bus[341]), .ZN(n10041) );
  ND2D1BWP30P140LVT U14721 ( .A1(n10042), .A2(n10041), .ZN(N1004) );
  AOI22D1BWP30P140LVT U14722 ( .A1(n10638), .A2(i_data_bus[359]), .B1(n10635), 
        .B2(i_data_bus[263]), .ZN(n10044) );
  AOI22D1BWP30P140LVT U14723 ( .A1(n10637), .A2(i_data_bus[295]), .B1(n10636), 
        .B2(i_data_bus[327]), .ZN(n10043) );
  ND2D1BWP30P140LVT U14724 ( .A1(n10044), .A2(n10043), .ZN(N990) );
  AOI22D1BWP30P140LVT U14725 ( .A1(n10638), .A2(i_data_bus[379]), .B1(n10635), 
        .B2(i_data_bus[283]), .ZN(n10046) );
  AOI22D1BWP30P140LVT U14726 ( .A1(n10637), .A2(i_data_bus[315]), .B1(n10636), 
        .B2(i_data_bus[347]), .ZN(n10045) );
  ND2D1BWP30P140LVT U14727 ( .A1(n10046), .A2(n10045), .ZN(N1010) );
  AOI22D1BWP30P140LVT U14728 ( .A1(n10638), .A2(i_data_bus[381]), .B1(n10635), 
        .B2(i_data_bus[285]), .ZN(n10048) );
  AOI22D1BWP30P140LVT U14729 ( .A1(n10637), .A2(i_data_bus[317]), .B1(n10636), 
        .B2(i_data_bus[349]), .ZN(n10047) );
  ND2D1BWP30P140LVT U14730 ( .A1(n10048), .A2(n10047), .ZN(N1012) );
  AOI22D1BWP30P140LVT U14731 ( .A1(n10638), .A2(i_data_bus[356]), .B1(n10635), 
        .B2(i_data_bus[260]), .ZN(n10050) );
  AOI22D1BWP30P140LVT U14732 ( .A1(n10637), .A2(i_data_bus[292]), .B1(n10636), 
        .B2(i_data_bus[324]), .ZN(n10049) );
  ND2D1BWP30P140LVT U14733 ( .A1(n10050), .A2(n10049), .ZN(N987) );
  AOI22D1BWP30P140LVT U14734 ( .A1(n10637), .A2(i_data_bus[301]), .B1(n10635), 
        .B2(i_data_bus[269]), .ZN(n10052) );
  AOI22D1BWP30P140LVT U14735 ( .A1(n10638), .A2(i_data_bus[365]), .B1(n10636), 
        .B2(i_data_bus[333]), .ZN(n10051) );
  ND2D1BWP30P140LVT U14736 ( .A1(n10052), .A2(n10051), .ZN(N996) );
  AOI22D1BWP30P140LVT U14737 ( .A1(n10638), .A2(i_data_bus[360]), .B1(n10635), 
        .B2(i_data_bus[264]), .ZN(n10054) );
  AOI22D1BWP30P140LVT U14738 ( .A1(n10637), .A2(i_data_bus[296]), .B1(n10636), 
        .B2(i_data_bus[328]), .ZN(n10053) );
  ND2D1BWP30P140LVT U14739 ( .A1(n10054), .A2(n10053), .ZN(N991) );
  AOI22D1BWP30P140LVT U14740 ( .A1(n10644), .A2(i_data_bus[16]), .B1(n10643), 
        .B2(i_data_bus[80]), .ZN(n10056) );
  AOI22D1BWP30P140LVT U14741 ( .A1(n10646), .A2(i_data_bus[48]), .B1(n10645), 
        .B2(i_data_bus[112]), .ZN(n10055) );
  ND2D1BWP30P140LVT U14742 ( .A1(n10056), .A2(n10055), .ZN(N559) );
  AOI22D1BWP30P140LVT U14743 ( .A1(n10644), .A2(i_data_bus[27]), .B1(n10643), 
        .B2(i_data_bus[91]), .ZN(n10058) );
  AOI22D1BWP30P140LVT U14744 ( .A1(n10646), .A2(i_data_bus[59]), .B1(n10645), 
        .B2(i_data_bus[123]), .ZN(n10057) );
  ND2D1BWP30P140LVT U14745 ( .A1(n10058), .A2(n10057), .ZN(N570) );
  AOI22D1BWP30P140LVT U14746 ( .A1(n10644), .A2(i_data_bus[1]), .B1(n10643), 
        .B2(i_data_bus[65]), .ZN(n10060) );
  AOI22D1BWP30P140LVT U14747 ( .A1(n10646), .A2(i_data_bus[33]), .B1(n10645), 
        .B2(i_data_bus[97]), .ZN(n10059) );
  ND2D1BWP30P140LVT U14748 ( .A1(n10060), .A2(n10059), .ZN(N544) );
  AOI22D1BWP30P140LVT U14749 ( .A1(n10644), .A2(i_data_bus[20]), .B1(n10643), 
        .B2(i_data_bus[84]), .ZN(n10062) );
  AOI22D1BWP30P140LVT U14750 ( .A1(n10646), .A2(i_data_bus[52]), .B1(n10645), 
        .B2(i_data_bus[116]), .ZN(n10061) );
  ND2D1BWP30P140LVT U14751 ( .A1(n10062), .A2(n10061), .ZN(N563) );
  AOI22D1BWP30P140LVT U14752 ( .A1(n10644), .A2(i_data_bus[28]), .B1(n10643), 
        .B2(i_data_bus[92]), .ZN(n10064) );
  AOI22D1BWP30P140LVT U14753 ( .A1(n10646), .A2(i_data_bus[60]), .B1(n10645), 
        .B2(i_data_bus[124]), .ZN(n10063) );
  ND2D1BWP30P140LVT U14754 ( .A1(n10064), .A2(n10063), .ZN(N571) );
  AOI22D1BWP30P140LVT U14755 ( .A1(n10618), .A2(i_data_bus[942]), .B1(n10617), 
        .B2(i_data_bus[974]), .ZN(n10066) );
  AOI22D1BWP30P140LVT U14756 ( .A1(n10620), .A2(i_data_bus[910]), .B1(n10619), 
        .B2(i_data_bus[1006]), .ZN(n10065) );
  ND2D1BWP30P140LVT U14757 ( .A1(n10066), .A2(n10065), .ZN(N2097) );
  AOI22D1BWP30P140LVT U14758 ( .A1(n10618), .A2(i_data_bus[931]), .B1(n10617), 
        .B2(i_data_bus[963]), .ZN(n10068) );
  AOI22D1BWP30P140LVT U14759 ( .A1(n10620), .A2(i_data_bus[899]), .B1(n10619), 
        .B2(i_data_bus[995]), .ZN(n10067) );
  ND2D1BWP30P140LVT U14760 ( .A1(n10068), .A2(n10067), .ZN(N2086) );
  AOI22D1BWP30P140LVT U14761 ( .A1(n10618), .A2(i_data_bus[945]), .B1(n10617), 
        .B2(i_data_bus[977]), .ZN(n10070) );
  AOI22D1BWP30P140LVT U14762 ( .A1(n10620), .A2(i_data_bus[913]), .B1(n10619), 
        .B2(i_data_bus[1009]), .ZN(n10069) );
  ND2D1BWP30P140LVT U14763 ( .A1(n10070), .A2(n10069), .ZN(N2100) );
  AOI22D1BWP30P140LVT U14764 ( .A1(n10618), .A2(i_data_bus[959]), .B1(n10617), 
        .B2(i_data_bus[991]), .ZN(n10072) );
  AOI22D1BWP30P140LVT U14765 ( .A1(n10620), .A2(i_data_bus[927]), .B1(n10619), 
        .B2(i_data_bus[1023]), .ZN(n10071) );
  ND2D1BWP30P140LVT U14766 ( .A1(n10072), .A2(n10071), .ZN(N2114) );
  AOI22D1BWP30P140LVT U14767 ( .A1(n10618), .A2(i_data_bus[944]), .B1(n10617), 
        .B2(i_data_bus[976]), .ZN(n10074) );
  AOI22D1BWP30P140LVT U14768 ( .A1(n10620), .A2(i_data_bus[912]), .B1(n10619), 
        .B2(i_data_bus[1008]), .ZN(n10073) );
  ND2D1BWP30P140LVT U14769 ( .A1(n10074), .A2(n10073), .ZN(N2099) );
  AOI22D1BWP30P140LVT U14770 ( .A1(n10646), .A2(i_data_bus[36]), .B1(n10643), 
        .B2(i_data_bus[68]), .ZN(n10076) );
  AOI22D1BWP30P140LVT U14771 ( .A1(n10645), .A2(i_data_bus[100]), .B1(n10644), 
        .B2(i_data_bus[4]), .ZN(n10075) );
  ND2D1BWP30P140LVT U14772 ( .A1(n10076), .A2(n10075), .ZN(N547) );
  AOI22D1BWP30P140LVT U14773 ( .A1(n10645), .A2(i_data_bus[113]), .B1(n10643), 
        .B2(i_data_bus[81]), .ZN(n10078) );
  AOI22D1BWP30P140LVT U14774 ( .A1(n10646), .A2(i_data_bus[49]), .B1(n10644), 
        .B2(i_data_bus[17]), .ZN(n10077) );
  ND2D1BWP30P140LVT U14775 ( .A1(n10078), .A2(n10077), .ZN(N560) );
  AOI22D1BWP30P140LVT U14776 ( .A1(n10646), .A2(i_data_bus[56]), .B1(n10643), 
        .B2(i_data_bus[88]), .ZN(n10080) );
  AOI22D1BWP30P140LVT U14777 ( .A1(n10645), .A2(i_data_bus[120]), .B1(n10644), 
        .B2(i_data_bus[24]), .ZN(n10079) );
  ND2D1BWP30P140LVT U14778 ( .A1(n10080), .A2(n10079), .ZN(N567) );
  AOI22D1BWP30P140LVT U14779 ( .A1(n10645), .A2(i_data_bus[104]), .B1(n10643), 
        .B2(i_data_bus[72]), .ZN(n10082) );
  AOI22D1BWP30P140LVT U14780 ( .A1(n10646), .A2(i_data_bus[40]), .B1(n10644), 
        .B2(i_data_bus[8]), .ZN(n10081) );
  ND2D1BWP30P140LVT U14781 ( .A1(n10082), .A2(n10081), .ZN(N551) );
  AOI22D1BWP30P140LVT U14782 ( .A1(n10646), .A2(i_data_bus[46]), .B1(n10643), 
        .B2(i_data_bus[78]), .ZN(n10084) );
  AOI22D1BWP30P140LVT U14783 ( .A1(n10645), .A2(i_data_bus[110]), .B1(n10644), 
        .B2(i_data_bus[14]), .ZN(n10083) );
  ND2D1BWP30P140LVT U14784 ( .A1(n10084), .A2(n10083), .ZN(N557) );
  AOI22D1BWP30P140LVT U14785 ( .A1(n10645), .A2(i_data_bus[102]), .B1(n10643), 
        .B2(i_data_bus[70]), .ZN(n10086) );
  AOI22D1BWP30P140LVT U14786 ( .A1(n10646), .A2(i_data_bus[38]), .B1(n10644), 
        .B2(i_data_bus[6]), .ZN(n10085) );
  ND2D1BWP30P140LVT U14787 ( .A1(n10086), .A2(n10085), .ZN(N549) );
  AOI22D1BWP30P140LVT U14788 ( .A1(n10646), .A2(i_data_bus[53]), .B1(n10643), 
        .B2(i_data_bus[85]), .ZN(n10088) );
  AOI22D1BWP30P140LVT U14789 ( .A1(n10645), .A2(i_data_bus[117]), .B1(n10644), 
        .B2(i_data_bus[21]), .ZN(n10087) );
  ND2D1BWP30P140LVT U14790 ( .A1(n10088), .A2(n10087), .ZN(N564) );
  AOI22D1BWP30P140LVT U14791 ( .A1(n10646), .A2(i_data_bus[55]), .B1(n10643), 
        .B2(i_data_bus[87]), .ZN(n10090) );
  AOI22D1BWP30P140LVT U14792 ( .A1(n10645), .A2(i_data_bus[119]), .B1(n10644), 
        .B2(i_data_bus[23]), .ZN(n10089) );
  ND2D1BWP30P140LVT U14793 ( .A1(n10090), .A2(n10089), .ZN(N566) );
  AOI22D1BWP30P140LVT U14794 ( .A1(n10646), .A2(i_data_bus[47]), .B1(n10643), 
        .B2(i_data_bus[79]), .ZN(n10092) );
  AOI22D1BWP30P140LVT U14795 ( .A1(n10645), .A2(i_data_bus[111]), .B1(n10644), 
        .B2(i_data_bus[15]), .ZN(n10091) );
  ND2D1BWP30P140LVT U14796 ( .A1(n10092), .A2(n10091), .ZN(N558) );
  AOI22D1BWP30P140LVT U14797 ( .A1(n10620), .A2(i_data_bus[900]), .B1(n10617), 
        .B2(i_data_bus[964]), .ZN(n10094) );
  AOI22D1BWP30P140LVT U14798 ( .A1(n10619), .A2(i_data_bus[996]), .B1(n10618), 
        .B2(i_data_bus[932]), .ZN(n10093) );
  ND2D1BWP30P140LVT U14799 ( .A1(n10094), .A2(n10093), .ZN(N2087) );
  AOI22D1BWP30P140LVT U14800 ( .A1(n10619), .A2(i_data_bus[1022]), .B1(n10617), 
        .B2(i_data_bus[990]), .ZN(n10096) );
  AOI22D1BWP30P140LVT U14801 ( .A1(n10620), .A2(i_data_bus[926]), .B1(n10618), 
        .B2(i_data_bus[958]), .ZN(n10095) );
  ND2D1BWP30P140LVT U14802 ( .A1(n10096), .A2(n10095), .ZN(N2113) );
  AOI22D1BWP30P140LVT U14803 ( .A1(n10619), .A2(i_data_bus[1016]), .B1(n10617), 
        .B2(i_data_bus[984]), .ZN(n10098) );
  AOI22D1BWP30P140LVT U14804 ( .A1(n10620), .A2(i_data_bus[920]), .B1(n10618), 
        .B2(i_data_bus[952]), .ZN(n10097) );
  ND2D1BWP30P140LVT U14805 ( .A1(n10098), .A2(n10097), .ZN(N2107) );
  AOI22D1BWP30P140LVT U14806 ( .A1(n10620), .A2(i_data_bus[907]), .B1(n10617), 
        .B2(i_data_bus[971]), .ZN(n10100) );
  AOI22D1BWP30P140LVT U14807 ( .A1(n10619), .A2(i_data_bus[1003]), .B1(n10618), 
        .B2(i_data_bus[939]), .ZN(n10099) );
  ND2D1BWP30P140LVT U14808 ( .A1(n10100), .A2(n10099), .ZN(N2094) );
  AOI22D1BWP30P140LVT U14809 ( .A1(n10619), .A2(i_data_bus[1019]), .B1(n10617), 
        .B2(i_data_bus[987]), .ZN(n10102) );
  AOI22D1BWP30P140LVT U14810 ( .A1(n10620), .A2(i_data_bus[923]), .B1(n10618), 
        .B2(i_data_bus[955]), .ZN(n10101) );
  ND2D1BWP30P140LVT U14811 ( .A1(n10102), .A2(n10101), .ZN(N2110) );
  AOI22D1BWP30P140LVT U14812 ( .A1(n10619), .A2(i_data_bus[999]), .B1(n10617), 
        .B2(i_data_bus[967]), .ZN(n10104) );
  AOI22D1BWP30P140LVT U14813 ( .A1(n10620), .A2(i_data_bus[903]), .B1(n10618), 
        .B2(i_data_bus[935]), .ZN(n10103) );
  ND2D1BWP30P140LVT U14814 ( .A1(n10104), .A2(n10103), .ZN(N2090) );
  AOI22D1BWP30P140LVT U14815 ( .A1(n10620), .A2(i_data_bus[918]), .B1(n10617), 
        .B2(i_data_bus[982]), .ZN(n10106) );
  AOI22D1BWP30P140LVT U14816 ( .A1(n10619), .A2(i_data_bus[1014]), .B1(n10618), 
        .B2(i_data_bus[950]), .ZN(n10105) );
  ND2D1BWP30P140LVT U14817 ( .A1(n10106), .A2(n10105), .ZN(N2105) );
  AOI22D1BWP30P140LVT U14818 ( .A1(n10620), .A2(i_data_bus[902]), .B1(n10617), 
        .B2(i_data_bus[966]), .ZN(n10108) );
  AOI22D1BWP30P140LVT U14819 ( .A1(n10619), .A2(i_data_bus[998]), .B1(n10618), 
        .B2(i_data_bus[934]), .ZN(n10107) );
  ND2D1BWP30P140LVT U14820 ( .A1(n10108), .A2(n10107), .ZN(N2089) );
  AOI22D1BWP30P140LVT U14821 ( .A1(n10620), .A2(i_data_bus[897]), .B1(n10617), 
        .B2(i_data_bus[961]), .ZN(n10110) );
  AOI22D1BWP30P140LVT U14822 ( .A1(n10619), .A2(i_data_bus[993]), .B1(n10618), 
        .B2(i_data_bus[929]), .ZN(n10109) );
  ND2D1BWP30P140LVT U14823 ( .A1(n10110), .A2(n10109), .ZN(N2084) );
  AOI22D1BWP30P140LVT U14824 ( .A1(n10619), .A2(i_data_bus[1015]), .B1(n10617), 
        .B2(i_data_bus[983]), .ZN(n10112) );
  AOI22D1BWP30P140LVT U14825 ( .A1(n10620), .A2(i_data_bus[919]), .B1(n10618), 
        .B2(i_data_bus[951]), .ZN(n10111) );
  ND2D1BWP30P140LVT U14826 ( .A1(n10112), .A2(n10111), .ZN(N2106) );
  AOI22D1BWP30P140LVT U14827 ( .A1(n10620), .A2(i_data_bus[915]), .B1(n10617), 
        .B2(i_data_bus[979]), .ZN(n10114) );
  AOI22D1BWP30P140LVT U14828 ( .A1(n10619), .A2(i_data_bus[1011]), .B1(n10618), 
        .B2(i_data_bus[947]), .ZN(n10113) );
  ND2D1BWP30P140LVT U14829 ( .A1(n10114), .A2(n10113), .ZN(N2102) );
  AOI22D1BWP30P140LVT U14830 ( .A1(n10619), .A2(i_data_bus[1004]), .B1(n10617), 
        .B2(i_data_bus[972]), .ZN(n10116) );
  AOI22D1BWP30P140LVT U14831 ( .A1(n10620), .A2(i_data_bus[908]), .B1(n10618), 
        .B2(i_data_bus[940]), .ZN(n10115) );
  ND2D1BWP30P140LVT U14832 ( .A1(n10116), .A2(n10115), .ZN(N2095) );
  AOI22D1BWP30P140LVT U14833 ( .A1(n10620), .A2(i_data_bus[911]), .B1(n10617), 
        .B2(i_data_bus[975]), .ZN(n10118) );
  AOI22D1BWP30P140LVT U14834 ( .A1(n10619), .A2(i_data_bus[1007]), .B1(n10618), 
        .B2(i_data_bus[943]), .ZN(n10117) );
  ND2D1BWP30P140LVT U14835 ( .A1(n10118), .A2(n10117), .ZN(N2098) );
  AOI22D1BWP30P140LVT U14836 ( .A1(n10622), .A2(i_data_bus[809]), .B1(n9749), 
        .B2(i_data_bus[873]), .ZN(n10120) );
  AOI22D1BWP30P140LVT U14837 ( .A1(n10623), .A2(i_data_bus[841]), .B1(n10621), 
        .B2(i_data_bus[777]), .ZN(n10119) );
  ND2D1BWP30P140LVT U14838 ( .A1(n10120), .A2(n10119), .ZN(N1872) );
  AOI22D1BWP30P140LVT U14839 ( .A1(n10622), .A2(i_data_bus[828]), .B1(n9749), 
        .B2(i_data_bus[892]), .ZN(n10122) );
  AOI22D1BWP30P140LVT U14840 ( .A1(n10623), .A2(i_data_bus[860]), .B1(n10621), 
        .B2(i_data_bus[796]), .ZN(n10121) );
  ND2D1BWP30P140LVT U14841 ( .A1(n10122), .A2(n10121), .ZN(N1891) );
  AOI22D1BWP30P140LVT U14842 ( .A1(n10623), .A2(i_data_bus[844]), .B1(n9749), 
        .B2(i_data_bus[876]), .ZN(n10124) );
  AOI22D1BWP30P140LVT U14843 ( .A1(n10622), .A2(i_data_bus[812]), .B1(n10621), 
        .B2(i_data_bus[780]), .ZN(n10123) );
  ND2D1BWP30P140LVT U14844 ( .A1(n10124), .A2(n10123), .ZN(N1875) );
  AOI22D1BWP30P140LVT U14845 ( .A1(n10622), .A2(i_data_bus[826]), .B1(n9749), 
        .B2(i_data_bus[890]), .ZN(n10126) );
  AOI22D1BWP30P140LVT U14846 ( .A1(n10623), .A2(i_data_bus[858]), .B1(n10621), 
        .B2(i_data_bus[794]), .ZN(n10125) );
  ND2D1BWP30P140LVT U14847 ( .A1(n10126), .A2(n10125), .ZN(N1889) );
  AOI22D1BWP30P140LVT U14848 ( .A1(n10622), .A2(i_data_bus[810]), .B1(n9749), 
        .B2(i_data_bus[874]), .ZN(n10128) );
  AOI22D1BWP30P140LVT U14849 ( .A1(n10623), .A2(i_data_bus[842]), .B1(n10621), 
        .B2(i_data_bus[778]), .ZN(n10127) );
  ND2D1BWP30P140LVT U14850 ( .A1(n10128), .A2(n10127), .ZN(N1873) );
  AOI22D1BWP30P140LVT U14851 ( .A1(n10622), .A2(i_data_bus[816]), .B1(n9749), 
        .B2(i_data_bus[880]), .ZN(n10130) );
  AOI22D1BWP30P140LVT U14852 ( .A1(n10623), .A2(i_data_bus[848]), .B1(n10621), 
        .B2(i_data_bus[784]), .ZN(n10129) );
  ND2D1BWP30P140LVT U14853 ( .A1(n10130), .A2(n10129), .ZN(N1879) );
  AOI22D1BWP30P140LVT U14854 ( .A1(n10622), .A2(i_data_bus[811]), .B1(n9749), 
        .B2(i_data_bus[875]), .ZN(n10132) );
  AOI22D1BWP30P140LVT U14855 ( .A1(n10623), .A2(i_data_bus[843]), .B1(n10621), 
        .B2(i_data_bus[779]), .ZN(n10131) );
  ND2D1BWP30P140LVT U14856 ( .A1(n10132), .A2(n10131), .ZN(N1874) );
  AOI22D1BWP30P140LVT U14857 ( .A1(n10637), .A2(i_data_bus[316]), .B1(n10636), 
        .B2(i_data_bus[348]), .ZN(n10134) );
  AOI22D1BWP30P140LVT U14858 ( .A1(n10638), .A2(i_data_bus[380]), .B1(n10635), 
        .B2(i_data_bus[284]), .ZN(n10133) );
  ND2D1BWP30P140LVT U14859 ( .A1(n10134), .A2(n10133), .ZN(N1011) );
  AOI22D1BWP30P140LVT U14860 ( .A1(n10638), .A2(i_data_bus[361]), .B1(n10637), 
        .B2(i_data_bus[297]), .ZN(n10136) );
  AOI22D1BWP30P140LVT U14861 ( .A1(n10636), .A2(i_data_bus[329]), .B1(n10635), 
        .B2(i_data_bus[265]), .ZN(n10135) );
  ND2D1BWP30P140LVT U14862 ( .A1(n10136), .A2(n10135), .ZN(N992) );
  AOI22D1BWP30P140LVT U14863 ( .A1(n10638), .A2(i_data_bus[362]), .B1(n10637), 
        .B2(i_data_bus[298]), .ZN(n10138) );
  AOI22D1BWP30P140LVT U14864 ( .A1(n10636), .A2(i_data_bus[330]), .B1(n10635), 
        .B2(i_data_bus[266]), .ZN(n10137) );
  ND2D1BWP30P140LVT U14865 ( .A1(n10138), .A2(n10137), .ZN(N993) );
  AOI22D1BWP30P140LVT U14866 ( .A1(n10637), .A2(i_data_bus[299]), .B1(n10636), 
        .B2(i_data_bus[331]), .ZN(n10140) );
  AOI22D1BWP30P140LVT U14867 ( .A1(n10638), .A2(i_data_bus[363]), .B1(n10635), 
        .B2(i_data_bus[267]), .ZN(n10139) );
  ND2D1BWP30P140LVT U14868 ( .A1(n10140), .A2(n10139), .ZN(N994) );
  AOI22D1BWP30P140LVT U14869 ( .A1(n10637), .A2(i_data_bus[300]), .B1(n10636), 
        .B2(i_data_bus[332]), .ZN(n10142) );
  AOI22D1BWP30P140LVT U14870 ( .A1(n10638), .A2(i_data_bus[364]), .B1(n10635), 
        .B2(i_data_bus[268]), .ZN(n10141) );
  ND2D1BWP30P140LVT U14871 ( .A1(n10142), .A2(n10141), .ZN(N995) );
  AOI22D1BWP30P140LVT U14872 ( .A1(n10637), .A2(i_data_bus[302]), .B1(n10636), 
        .B2(i_data_bus[334]), .ZN(n10144) );
  AOI22D1BWP30P140LVT U14873 ( .A1(n10638), .A2(i_data_bus[366]), .B1(n10635), 
        .B2(i_data_bus[270]), .ZN(n10143) );
  ND2D1BWP30P140LVT U14874 ( .A1(n10144), .A2(n10143), .ZN(N997) );
  AOI22D1BWP30P140LVT U14875 ( .A1(n10638), .A2(i_data_bus[374]), .B1(n10636), 
        .B2(i_data_bus[342]), .ZN(n10146) );
  AOI22D1BWP30P140LVT U14876 ( .A1(n10637), .A2(i_data_bus[310]), .B1(n10635), 
        .B2(i_data_bus[278]), .ZN(n10145) );
  ND2D1BWP30P140LVT U14877 ( .A1(n10146), .A2(n10145), .ZN(N1005) );
  AOI22D1BWP30P140LVT U14878 ( .A1(n10638), .A2(i_data_bus[367]), .B1(n10636), 
        .B2(i_data_bus[335]), .ZN(n10148) );
  AOI22D1BWP30P140LVT U14879 ( .A1(n10637), .A2(i_data_bus[303]), .B1(n10635), 
        .B2(i_data_bus[271]), .ZN(n10147) );
  ND2D1BWP30P140LVT U14880 ( .A1(n10148), .A2(n10147), .ZN(N998) );
  AOI22D1BWP30P140LVT U14881 ( .A1(n10637), .A2(i_data_bus[312]), .B1(n10636), 
        .B2(i_data_bus[344]), .ZN(n10150) );
  AOI22D1BWP30P140LVT U14882 ( .A1(n10638), .A2(i_data_bus[376]), .B1(n10635), 
        .B2(i_data_bus[280]), .ZN(n10149) );
  ND2D1BWP30P140LVT U14883 ( .A1(n10150), .A2(n10149), .ZN(N1007) );
  AOI22D1BWP30P140LVT U14884 ( .A1(n10638), .A2(i_data_bus[369]), .B1(n10636), 
        .B2(i_data_bus[337]), .ZN(n10152) );
  AOI22D1BWP30P140LVT U14885 ( .A1(n10637), .A2(i_data_bus[305]), .B1(n10635), 
        .B2(i_data_bus[273]), .ZN(n10151) );
  ND2D1BWP30P140LVT U14886 ( .A1(n10152), .A2(n10151), .ZN(N1000) );
  AOI22D1BWP30P140LVT U14887 ( .A1(n10638), .A2(i_data_bus[371]), .B1(n10636), 
        .B2(i_data_bus[339]), .ZN(n10154) );
  AOI22D1BWP30P140LVT U14888 ( .A1(n10637), .A2(i_data_bus[307]), .B1(n10635), 
        .B2(i_data_bus[275]), .ZN(n10153) );
  ND2D1BWP30P140LVT U14889 ( .A1(n10154), .A2(n10153), .ZN(N1002) );
  AOI22D1BWP30P140LVT U14890 ( .A1(n10638), .A2(i_data_bus[383]), .B1(n10637), 
        .B2(i_data_bus[319]), .ZN(n10156) );
  AOI22D1BWP30P140LVT U14891 ( .A1(n10636), .A2(i_data_bus[351]), .B1(n10635), 
        .B2(i_data_bus[287]), .ZN(n10155) );
  ND2D1BWP30P140LVT U14892 ( .A1(n10156), .A2(n10155), .ZN(N1014) );
  AOI22D1BWP30P140LVT U14893 ( .A1(n10638), .A2(i_data_bus[375]), .B1(n10636), 
        .B2(i_data_bus[343]), .ZN(n10158) );
  AOI22D1BWP30P140LVT U14894 ( .A1(n10637), .A2(i_data_bus[311]), .B1(n10635), 
        .B2(i_data_bus[279]), .ZN(n10157) );
  ND2D1BWP30P140LVT U14895 ( .A1(n10158), .A2(n10157), .ZN(N1006) );
  AOI22D1BWP30P140LVT U14896 ( .A1(n10638), .A2(i_data_bus[378]), .B1(n10636), 
        .B2(i_data_bus[346]), .ZN(n10160) );
  AOI22D1BWP30P140LVT U14897 ( .A1(n10637), .A2(i_data_bus[314]), .B1(n10635), 
        .B2(i_data_bus[282]), .ZN(n10159) );
  ND2D1BWP30P140LVT U14898 ( .A1(n10160), .A2(n10159), .ZN(N1009) );
  AOI22D1BWP30P140LVT U14899 ( .A1(n10638), .A2(i_data_bus[377]), .B1(n10636), 
        .B2(i_data_bus[345]), .ZN(n10162) );
  AOI22D1BWP30P140LVT U14900 ( .A1(n10637), .A2(i_data_bus[313]), .B1(n10635), 
        .B2(i_data_bus[281]), .ZN(n10161) );
  ND2D1BWP30P140LVT U14901 ( .A1(n10162), .A2(n10161), .ZN(N1008) );
  AOI22D1BWP30P140LVT U14902 ( .A1(n10637), .A2(i_data_bus[294]), .B1(n10636), 
        .B2(i_data_bus[326]), .ZN(n10164) );
  AOI22D1BWP30P140LVT U14903 ( .A1(n10638), .A2(i_data_bus[358]), .B1(n10635), 
        .B2(i_data_bus[262]), .ZN(n10163) );
  ND2D1BWP30P140LVT U14904 ( .A1(n10164), .A2(n10163), .ZN(N989) );
  AOI22D1BWP30P140LVT U14905 ( .A1(n10638), .A2(i_data_bus[354]), .B1(n10636), 
        .B2(i_data_bus[322]), .ZN(n10166) );
  AOI22D1BWP30P140LVT U14906 ( .A1(n10637), .A2(i_data_bus[290]), .B1(n10635), 
        .B2(i_data_bus[258]), .ZN(n10165) );
  ND2D1BWP30P140LVT U14907 ( .A1(n10166), .A2(n10165), .ZN(N985) );
  AOI22D1BWP30P140LVT U14908 ( .A1(n10638), .A2(i_data_bus[353]), .B1(n10637), 
        .B2(i_data_bus[289]), .ZN(n10168) );
  AOI22D1BWP30P140LVT U14909 ( .A1(n10636), .A2(i_data_bus[321]), .B1(n10635), 
        .B2(i_data_bus[257]), .ZN(n10167) );
  ND2D1BWP30P140LVT U14910 ( .A1(n10168), .A2(n10167), .ZN(N984) );
  AOI22D1BWP30P140LVT U14911 ( .A1(n10631), .A2(i_data_bus[618]), .B1(n10630), 
        .B2(i_data_bus[522]), .ZN(n10170) );
  AOI22D1BWP30P140LVT U14912 ( .A1(n10629), .A2(i_data_bus[554]), .B1(n10628), 
        .B2(i_data_bus[586]), .ZN(n10169) );
  ND2D1BWP30P140LVT U14913 ( .A1(n10170), .A2(n10169), .ZN(N1433) );
  AOI22D1BWP30P140LVT U14914 ( .A1(n10631), .A2(i_data_bus[632]), .B1(n10629), 
        .B2(i_data_bus[568]), .ZN(n10172) );
  AOI22D1BWP30P140LVT U14915 ( .A1(n10630), .A2(i_data_bus[536]), .B1(n10628), 
        .B2(i_data_bus[600]), .ZN(n10171) );
  AOI22D1BWP30P140LVT U14916 ( .A1(n10631), .A2(i_data_bus[628]), .B1(n10630), 
        .B2(i_data_bus[532]), .ZN(n10174) );
  AOI22D1BWP30P140LVT U14917 ( .A1(n10629), .A2(i_data_bus[564]), .B1(n10628), 
        .B2(i_data_bus[596]), .ZN(n10173) );
  ND2D1BWP30P140LVT U14918 ( .A1(n10174), .A2(n10173), .ZN(N1443) );
  AOI22D1BWP30P140LVT U14919 ( .A1(n10630), .A2(i_data_bus[535]), .B1(n10629), 
        .B2(i_data_bus[567]), .ZN(n10176) );
  AOI22D1BWP30P140LVT U14920 ( .A1(n10631), .A2(i_data_bus[631]), .B1(n10628), 
        .B2(i_data_bus[599]), .ZN(n10175) );
  AOI22D1BWP30P140LVT U14921 ( .A1(n10630), .A2(i_data_bus[530]), .B1(n10629), 
        .B2(i_data_bus[562]), .ZN(n10178) );
  AOI22D1BWP30P140LVT U14922 ( .A1(n10631), .A2(i_data_bus[626]), .B1(n10628), 
        .B2(i_data_bus[594]), .ZN(n10177) );
  AOI22D1BWP30P140LVT U14923 ( .A1(n10630), .A2(i_data_bus[541]), .B1(n10629), 
        .B2(i_data_bus[573]), .ZN(n10180) );
  AOI22D1BWP30P140LVT U14924 ( .A1(n10631), .A2(i_data_bus[637]), .B1(n10628), 
        .B2(i_data_bus[605]), .ZN(n10179) );
  AOI22D1BWP30P140LVT U14925 ( .A1(n10631), .A2(i_data_bus[639]), .B1(n10629), 
        .B2(i_data_bus[575]), .ZN(n10182) );
  AOI22D1BWP30P140LVT U14926 ( .A1(n10630), .A2(i_data_bus[543]), .B1(n10628), 
        .B2(i_data_bus[607]), .ZN(n10181) );
  AOI22D1BWP30P140LVT U14927 ( .A1(n10631), .A2(i_data_bus[633]), .B1(n10630), 
        .B2(i_data_bus[537]), .ZN(n10184) );
  AOI22D1BWP30P140LVT U14928 ( .A1(n10629), .A2(i_data_bus[569]), .B1(n10628), 
        .B2(i_data_bus[601]), .ZN(n10183) );
  ND2D1BWP30P140LVT U14929 ( .A1(n10184), .A2(n10183), .ZN(N1448) );
  AOI22D1BWP30P140LVT U14930 ( .A1(n10631), .A2(i_data_bus[634]), .B1(n10630), 
        .B2(i_data_bus[538]), .ZN(n10186) );
  AOI22D1BWP30P140LVT U14931 ( .A1(n10629), .A2(i_data_bus[570]), .B1(n10628), 
        .B2(i_data_bus[602]), .ZN(n10185) );
  ND2D1BWP30P140LVT U14932 ( .A1(n10186), .A2(n10185), .ZN(N1449) );
  AOI22D1BWP30P140LVT U14933 ( .A1(n10631), .A2(i_data_bus[636]), .B1(n10630), 
        .B2(i_data_bus[540]), .ZN(n10188) );
  AOI22D1BWP30P140LVT U14934 ( .A1(n10629), .A2(i_data_bus[572]), .B1(n10628), 
        .B2(i_data_bus[604]), .ZN(n10187) );
  ND2D1BWP30P140LVT U14935 ( .A1(n10188), .A2(n10187), .ZN(N1451) );
  AOI22D1BWP30P140LVT U14936 ( .A1(n10631), .A2(i_data_bus[623]), .B1(n10630), 
        .B2(i_data_bus[527]), .ZN(n10190) );
  AOI22D1BWP30P140LVT U14937 ( .A1(n10629), .A2(i_data_bus[559]), .B1(n10628), 
        .B2(i_data_bus[591]), .ZN(n10189) );
  ND2D1BWP30P140LVT U14938 ( .A1(n10190), .A2(n10189), .ZN(N1438) );
  AOI22D1BWP30P140LVT U14939 ( .A1(n10630), .A2(i_data_bus[515]), .B1(n10629), 
        .B2(i_data_bus[547]), .ZN(n10192) );
  AOI22D1BWP30P140LVT U14940 ( .A1(n10631), .A2(i_data_bus[611]), .B1(n10628), 
        .B2(i_data_bus[579]), .ZN(n10191) );
  AOI22D1BWP30P140LVT U14941 ( .A1(n10630), .A2(i_data_bus[514]), .B1(n10629), 
        .B2(i_data_bus[546]), .ZN(n10194) );
  AOI22D1BWP30P140LVT U14942 ( .A1(n10631), .A2(i_data_bus[610]), .B1(n10628), 
        .B2(i_data_bus[578]), .ZN(n10193) );
  AOI22D1BWP30P140LVT U14943 ( .A1(n10631), .A2(i_data_bus[609]), .B1(n10629), 
        .B2(i_data_bus[545]), .ZN(n10196) );
  AOI22D1BWP30P140LVT U14944 ( .A1(n10630), .A2(i_data_bus[513]), .B1(n10628), 
        .B2(i_data_bus[577]), .ZN(n10195) );
  AOI22D1BWP30P140LVT U14945 ( .A1(n10631), .A2(i_data_bus[625]), .B1(n10630), 
        .B2(i_data_bus[529]), .ZN(n10198) );
  AOI22D1BWP30P140LVT U14946 ( .A1(n10629), .A2(i_data_bus[561]), .B1(n10628), 
        .B2(i_data_bus[593]), .ZN(n10197) );
  ND2D1BWP30P140LVT U14947 ( .A1(n10198), .A2(n10197), .ZN(N1440) );
  AOI22D1BWP30P140LVT U14948 ( .A1(n10631), .A2(i_data_bus[629]), .B1(n10629), 
        .B2(i_data_bus[565]), .ZN(n10200) );
  AOI22D1BWP30P140LVT U14949 ( .A1(n10630), .A2(i_data_bus[533]), .B1(n10628), 
        .B2(i_data_bus[597]), .ZN(n10199) );
  AOI22D1BWP30P140LVT U14950 ( .A1(n10631), .A2(i_data_bus[619]), .B1(n10629), 
        .B2(i_data_bus[555]), .ZN(n10202) );
  AOI22D1BWP30P140LVT U14951 ( .A1(n10630), .A2(i_data_bus[523]), .B1(n10628), 
        .B2(i_data_bus[587]), .ZN(n10201) );
  AOI22D1BWP30P140LVT U14952 ( .A1(n10627), .A2(i_data_bus[688]), .B1(n10625), 
        .B2(i_data_bus[656]), .ZN(n10204) );
  AOI22D1BWP30P140LVT U14953 ( .A1(n10626), .A2(i_data_bus[720]), .B1(n10624), 
        .B2(i_data_bus[752]), .ZN(n10203) );
  AOI22D1BWP30P140LVT U14954 ( .A1(n10627), .A2(i_data_bus[697]), .B1(n10626), 
        .B2(i_data_bus[729]), .ZN(n10206) );
  AOI22D1BWP30P140LVT U14955 ( .A1(n10625), .A2(i_data_bus[665]), .B1(n10624), 
        .B2(i_data_bus[761]), .ZN(n10205) );
  AOI22D1BWP30P140LVT U14956 ( .A1(n10626), .A2(i_data_bus[726]), .B1(n10625), 
        .B2(i_data_bus[662]), .ZN(n10208) );
  AOI22D1BWP30P140LVT U14957 ( .A1(n10627), .A2(i_data_bus[694]), .B1(n10624), 
        .B2(i_data_bus[758]), .ZN(n10207) );
  AOI22D1BWP30P140LVT U14958 ( .A1(n10627), .A2(i_data_bus[699]), .B1(n10626), 
        .B2(i_data_bus[731]), .ZN(n10210) );
  AOI22D1BWP30P140LVT U14959 ( .A1(n10625), .A2(i_data_bus[667]), .B1(n10624), 
        .B2(i_data_bus[763]), .ZN(n10209) );
  AOI22D1BWP30P140LVT U14960 ( .A1(n10627), .A2(i_data_bus[691]), .B1(n10626), 
        .B2(i_data_bus[723]), .ZN(n10212) );
  AOI22D1BWP30P140LVT U14961 ( .A1(n10625), .A2(i_data_bus[659]), .B1(n10624), 
        .B2(i_data_bus[755]), .ZN(n10211) );
  AOI22D1BWP30P140LVT U14962 ( .A1(n10627), .A2(i_data_bus[693]), .B1(n10625), 
        .B2(i_data_bus[661]), .ZN(n10214) );
  AOI22D1BWP30P140LVT U14963 ( .A1(n10626), .A2(i_data_bus[725]), .B1(n10624), 
        .B2(i_data_bus[757]), .ZN(n10213) );
  AOI22D1BWP30P140LVT U14964 ( .A1(n10627), .A2(i_data_bus[700]), .B1(n10625), 
        .B2(i_data_bus[668]), .ZN(n10216) );
  AOI22D1BWP30P140LVT U14965 ( .A1(n10626), .A2(i_data_bus[732]), .B1(n10624), 
        .B2(i_data_bus[764]), .ZN(n10215) );
  AOI22D1BWP30P140LVT U14966 ( .A1(n10627), .A2(i_data_bus[702]), .B1(n10625), 
        .B2(i_data_bus[670]), .ZN(n10218) );
  AOI22D1BWP30P140LVT U14967 ( .A1(n10626), .A2(i_data_bus[734]), .B1(n10624), 
        .B2(i_data_bus[766]), .ZN(n10217) );
  AOI22D1BWP30P140LVT U14968 ( .A1(n10627), .A2(i_data_bus[689]), .B1(n10626), 
        .B2(i_data_bus[721]), .ZN(n10220) );
  AOI22D1BWP30P140LVT U14969 ( .A1(n10625), .A2(i_data_bus[657]), .B1(n10624), 
        .B2(i_data_bus[753]), .ZN(n10219) );
  AOI22D1BWP30P140LVT U14970 ( .A1(n10627), .A2(i_data_bus[676]), .B1(n10625), 
        .B2(i_data_bus[644]), .ZN(n10222) );
  AOI22D1BWP30P140LVT U14971 ( .A1(n10626), .A2(i_data_bus[708]), .B1(n10624), 
        .B2(i_data_bus[740]), .ZN(n10221) );
  AOI22D1BWP30P140LVT U14972 ( .A1(n10627), .A2(i_data_bus[682]), .B1(n10626), 
        .B2(i_data_bus[714]), .ZN(n10224) );
  AOI22D1BWP30P140LVT U14973 ( .A1(n10625), .A2(i_data_bus[650]), .B1(n10624), 
        .B2(i_data_bus[746]), .ZN(n10223) );
  AOI22D1BWP30P140LVT U14974 ( .A1(n10627), .A2(i_data_bus[685]), .B1(n10626), 
        .B2(i_data_bus[717]), .ZN(n10226) );
  AOI22D1BWP30P140LVT U14975 ( .A1(n10625), .A2(i_data_bus[653]), .B1(n10624), 
        .B2(i_data_bus[749]), .ZN(n10225) );
  AOI22D1BWP30P140LVT U14976 ( .A1(n10627), .A2(i_data_bus[680]), .B1(n10626), 
        .B2(i_data_bus[712]), .ZN(n10228) );
  AOI22D1BWP30P140LVT U14977 ( .A1(n10625), .A2(i_data_bus[648]), .B1(n10624), 
        .B2(i_data_bus[744]), .ZN(n10227) );
  AOI22D1BWP30P140LVT U14978 ( .A1(n10642), .A2(i_data_bus[137]), .B1(n10640), 
        .B2(i_data_bus[169]), .ZN(n10230) );
  AOI22D1BWP30P140LVT U14979 ( .A1(n10641), .A2(i_data_bus[233]), .B1(n10639), 
        .B2(i_data_bus[201]), .ZN(n10229) );
  AOI22D1BWP30P140LVT U14980 ( .A1(n10642), .A2(i_data_bus[140]), .B1(n10640), 
        .B2(i_data_bus[172]), .ZN(n10232) );
  AOI22D1BWP30P140LVT U14981 ( .A1(n10641), .A2(i_data_bus[236]), .B1(n10639), 
        .B2(i_data_bus[204]), .ZN(n10231) );
  AOI22D1BWP30P140LVT U14982 ( .A1(n10642), .A2(i_data_bus[130]), .B1(n10641), 
        .B2(i_data_bus[226]), .ZN(n10234) );
  AOI22D1BWP30P140LVT U14983 ( .A1(n10640), .A2(i_data_bus[162]), .B1(n10639), 
        .B2(i_data_bus[194]), .ZN(n10233) );
  AOI22D1BWP30P140LVT U14984 ( .A1(n10642), .A2(i_data_bus[136]), .B1(n10641), 
        .B2(i_data_bus[232]), .ZN(n10236) );
  AOI22D1BWP30P140LVT U14985 ( .A1(n10640), .A2(i_data_bus[168]), .B1(n10639), 
        .B2(i_data_bus[200]), .ZN(n10235) );
  AOI22D1BWP30P140LVT U14986 ( .A1(n10642), .A2(i_data_bus[143]), .B1(n10641), 
        .B2(i_data_bus[239]), .ZN(n10238) );
  AOI22D1BWP30P140LVT U14987 ( .A1(n10640), .A2(i_data_bus[175]), .B1(n10639), 
        .B2(i_data_bus[207]), .ZN(n10237) );
  AOI22D1BWP30P140LVT U14988 ( .A1(n10642), .A2(i_data_bus[145]), .B1(n10641), 
        .B2(i_data_bus[241]), .ZN(n10240) );
  AOI22D1BWP30P140LVT U14989 ( .A1(n10640), .A2(i_data_bus[177]), .B1(n10639), 
        .B2(i_data_bus[209]), .ZN(n10239) );
  AOI22D1BWP30P140LVT U14990 ( .A1(n10642), .A2(i_data_bus[150]), .B1(n10641), 
        .B2(i_data_bus[246]), .ZN(n10242) );
  AOI22D1BWP30P140LVT U14991 ( .A1(n10640), .A2(i_data_bus[182]), .B1(n10639), 
        .B2(i_data_bus[214]), .ZN(n10241) );
  AOI22D1BWP30P140LVT U14992 ( .A1(n10642), .A2(i_data_bus[141]), .B1(n10641), 
        .B2(i_data_bus[237]), .ZN(n10244) );
  AOI22D1BWP30P140LVT U14993 ( .A1(n10640), .A2(i_data_bus[173]), .B1(n10639), 
        .B2(i_data_bus[205]), .ZN(n10243) );
  AOI22D1BWP30P140LVT U14994 ( .A1(n10642), .A2(i_data_bus[152]), .B1(n10640), 
        .B2(i_data_bus[184]), .ZN(n10246) );
  AOI22D1BWP30P140LVT U14995 ( .A1(n10641), .A2(i_data_bus[248]), .B1(n10639), 
        .B2(i_data_bus[216]), .ZN(n10245) );
  AOI22D1BWP30P140LVT U14996 ( .A1(n10642), .A2(i_data_bus[134]), .B1(n10640), 
        .B2(i_data_bus[166]), .ZN(n10248) );
  AOI22D1BWP30P140LVT U14997 ( .A1(n10641), .A2(i_data_bus[230]), .B1(n10639), 
        .B2(i_data_bus[198]), .ZN(n10247) );
  AOI22D1BWP30P140LVT U14998 ( .A1(n10642), .A2(i_data_bus[157]), .B1(n10640), 
        .B2(i_data_bus[189]), .ZN(n10250) );
  AOI22D1BWP30P140LVT U14999 ( .A1(n10641), .A2(i_data_bus[253]), .B1(n10639), 
        .B2(i_data_bus[221]), .ZN(n10249) );
  AOI22D1BWP30P140LVT U15000 ( .A1(n10642), .A2(i_data_bus[158]), .B1(n10641), 
        .B2(i_data_bus[254]), .ZN(n10252) );
  AOI22D1BWP30P140LVT U15001 ( .A1(n10640), .A2(i_data_bus[190]), .B1(n10639), 
        .B2(i_data_bus[222]), .ZN(n10251) );
  AOI22D1BWP30P140LVT U15002 ( .A1(n10642), .A2(i_data_bus[139]), .B1(n10640), 
        .B2(i_data_bus[171]), .ZN(n10254) );
  AOI22D1BWP30P140LVT U15003 ( .A1(n10641), .A2(i_data_bus[235]), .B1(n10639), 
        .B2(i_data_bus[203]), .ZN(n10253) );
  AOI22D1BWP30P140LVT U15004 ( .A1(n10641), .A2(i_data_bus[255]), .B1(n10640), 
        .B2(i_data_bus[191]), .ZN(n10256) );
  AOI22D1BWP30P140LVT U15005 ( .A1(n10642), .A2(i_data_bus[159]), .B1(n10639), 
        .B2(i_data_bus[223]), .ZN(n10255) );
  AOI22D1BWP30P140LVT U15006 ( .A1(n10641), .A2(i_data_bus[240]), .B1(n10640), 
        .B2(i_data_bus[176]), .ZN(n10258) );
  AOI22D1BWP30P140LVT U15007 ( .A1(n10642), .A2(i_data_bus[144]), .B1(n10639), 
        .B2(i_data_bus[208]), .ZN(n10257) );
  AOI22D1BWP30P140LVT U15008 ( .A1(n10646), .A2(i_data_bus[45]), .B1(n10644), 
        .B2(i_data_bus[13]), .ZN(n10260) );
  AOI22D1BWP30P140LVT U15009 ( .A1(n10645), .A2(i_data_bus[109]), .B1(n10643), 
        .B2(i_data_bus[77]), .ZN(n10259) );
  AOI22D1BWP30P140LVT U15010 ( .A1(n10645), .A2(i_data_bus[108]), .B1(n10644), 
        .B2(i_data_bus[12]), .ZN(n10262) );
  AOI22D1BWP30P140LVT U15011 ( .A1(n10646), .A2(i_data_bus[44]), .B1(n10643), 
        .B2(i_data_bus[76]), .ZN(n10261) );
  AOI22D1BWP30P140LVT U15012 ( .A1(n10645), .A2(i_data_bus[107]), .B1(n10644), 
        .B2(i_data_bus[11]), .ZN(n10264) );
  AOI22D1BWP30P140LVT U15013 ( .A1(n10646), .A2(i_data_bus[43]), .B1(n10643), 
        .B2(i_data_bus[75]), .ZN(n10263) );
  AOI22D1BWP30P140LVT U15014 ( .A1(n10646), .A2(i_data_bus[42]), .B1(n10645), 
        .B2(i_data_bus[106]), .ZN(n10266) );
  AOI22D1BWP30P140LVT U15015 ( .A1(n10644), .A2(i_data_bus[10]), .B1(n10643), 
        .B2(i_data_bus[74]), .ZN(n10265) );
  AOI22D1BWP30P140LVT U15016 ( .A1(n10646), .A2(i_data_bus[54]), .B1(n10644), 
        .B2(i_data_bus[22]), .ZN(n10268) );
  AOI22D1BWP30P140LVT U15017 ( .A1(n10645), .A2(i_data_bus[118]), .B1(n10643), 
        .B2(i_data_bus[86]), .ZN(n10267) );
  AOI22D1BWP30P140LVT U15018 ( .A1(n10645), .A2(i_data_bus[101]), .B1(n10644), 
        .B2(i_data_bus[5]), .ZN(n10270) );
  AOI22D1BWP30P140LVT U15019 ( .A1(n10646), .A2(i_data_bus[37]), .B1(n10643), 
        .B2(i_data_bus[69]), .ZN(n10269) );
  AOI22D1BWP30P140LVT U15020 ( .A1(n10646), .A2(i_data_bus[41]), .B1(n10644), 
        .B2(i_data_bus[9]), .ZN(n10272) );
  AOI22D1BWP30P140LVT U15021 ( .A1(n10645), .A2(i_data_bus[105]), .B1(n10643), 
        .B2(i_data_bus[73]), .ZN(n10271) );
  AOI22D1BWP30P140LVT U15022 ( .A1(n10645), .A2(i_data_bus[103]), .B1(n10644), 
        .B2(i_data_bus[7]), .ZN(n10274) );
  AOI22D1BWP30P140LVT U15023 ( .A1(n10646), .A2(i_data_bus[39]), .B1(n10643), 
        .B2(i_data_bus[71]), .ZN(n10273) );
  AOI22D1BWP30P140LVT U15024 ( .A1(n10645), .A2(i_data_bus[125]), .B1(n10644), 
        .B2(i_data_bus[29]), .ZN(n10276) );
  AOI22D1BWP30P140LVT U15025 ( .A1(n10646), .A2(i_data_bus[61]), .B1(n10643), 
        .B2(i_data_bus[93]), .ZN(n10275) );
  AOI22D1BWP30P140LVT U15026 ( .A1(n10646), .A2(i_data_bus[58]), .B1(n10644), 
        .B2(i_data_bus[26]), .ZN(n10278) );
  AOI22D1BWP30P140LVT U15027 ( .A1(n10645), .A2(i_data_bus[122]), .B1(n10643), 
        .B2(i_data_bus[90]), .ZN(n10277) );
  AOI22D1BWP30P140LVT U15028 ( .A1(n10646), .A2(i_data_bus[57]), .B1(n10644), 
        .B2(i_data_bus[25]), .ZN(n10280) );
  AOI22D1BWP30P140LVT U15029 ( .A1(n10645), .A2(i_data_bus[121]), .B1(n10643), 
        .B2(i_data_bus[89]), .ZN(n10279) );
  AOI22D1BWP30P140LVT U15030 ( .A1(n10646), .A2(i_data_bus[63]), .B1(n10644), 
        .B2(i_data_bus[31]), .ZN(n10282) );
  AOI22D1BWP30P140LVT U15031 ( .A1(n10645), .A2(i_data_bus[127]), .B1(n10643), 
        .B2(i_data_bus[95]), .ZN(n10281) );
  AOI22D1BWP30P140LVT U15032 ( .A1(n10645), .A2(i_data_bus[115]), .B1(n10644), 
        .B2(i_data_bus[19]), .ZN(n10284) );
  AOI22D1BWP30P140LVT U15033 ( .A1(n10646), .A2(i_data_bus[51]), .B1(n10643), 
        .B2(i_data_bus[83]), .ZN(n10283) );
  AOI22D1BWP30P140LVT U15034 ( .A1(n10645), .A2(i_data_bus[99]), .B1(n10644), 
        .B2(i_data_bus[3]), .ZN(n10286) );
  AOI22D1BWP30P140LVT U15035 ( .A1(n10646), .A2(i_data_bus[35]), .B1(n10643), 
        .B2(i_data_bus[67]), .ZN(n10285) );
  AOI22D1BWP30P140LVT U15036 ( .A1(n10646), .A2(i_data_bus[62]), .B1(n10644), 
        .B2(i_data_bus[30]), .ZN(n10288) );
  AOI22D1BWP30P140LVT U15037 ( .A1(n10645), .A2(i_data_bus[126]), .B1(n10643), 
        .B2(i_data_bus[94]), .ZN(n10287) );
  AOI22D1BWP30P140LVT U15038 ( .A1(n10646), .A2(i_data_bus[50]), .B1(n10644), 
        .B2(i_data_bus[18]), .ZN(n10290) );
  AOI22D1BWP30P140LVT U15039 ( .A1(n10645), .A2(i_data_bus[114]), .B1(n10643), 
        .B2(i_data_bus[82]), .ZN(n10289) );
  AOI22D1BWP30P140LVT U15040 ( .A1(n10646), .A2(i_data_bus[34]), .B1(n10644), 
        .B2(i_data_bus[2]), .ZN(n10292) );
  AOI22D1BWP30P140LVT U15041 ( .A1(n10645), .A2(i_data_bus[98]), .B1(n10643), 
        .B2(i_data_bus[66]), .ZN(n10291) );
  NR3D0P7BWP30P140LVT U15042 ( .A1(inner_first_stage_valid_reg[62]), .A2(
        inner_first_stage_valid_reg[63]), .A3(n10380), .ZN(n10302) );
  NR3D0P7BWP30P140LVT U15043 ( .A1(inner_first_stage_valid_reg[61]), .A2(
        inner_first_stage_valid_reg[57]), .A3(inner_first_stage_valid_reg[59]), 
        .ZN(n10294) );
  IND3D1BWP30P140LVT U15044 ( .A1(inner_first_stage_valid_reg[60]), .B1(n10302), .B2(n10294), .ZN(n10300) );
  INR3D2BWP30P140LVT U15045 ( .A1(inner_first_stage_valid_reg[58]), .B1(
        inner_first_stage_valid_reg[56]), .B2(n10300), .ZN(n11760) );
  INVD1BWP30P140LVT U15046 ( .I(inner_first_stage_valid_reg[62]), .ZN(n10296)
         );
  INVD1BWP30P140LVT U15047 ( .I(inner_first_stage_valid_reg[63]), .ZN(n10298)
         );
  INR4D0BWP30P140LVT U15048 ( .A1(n10295), .B1(inner_first_stage_valid_reg[58]), .B2(inner_first_stage_valid_reg[56]), .B3(n10293), .ZN(n10304) );
  INVD1BWP30P140LVT U15049 ( .I(inner_first_stage_valid_reg[59]), .ZN(n10303)
         );
  INR3D2BWP30P140LVT U15050 ( .A1(inner_first_stage_valid_reg[57]), .B1(
        inner_first_stage_valid_reg[61]), .B2(n10299), .ZN(n11759) );
  INR3D0BWP30P140LVT U15051 ( .A1(n10294), .B1(inner_first_stage_valid_reg[56]), .B2(inner_first_stage_valid_reg[58]), .ZN(n10301) );
  NR4D0BWP30P140LVT U15052 ( .A1(n11760), .A2(n11759), .A3(n11762), .A4(n11761), .ZN(n10306) );
  INR3D2BWP30P140LVT U15053 ( .A1(inner_first_stage_valid_reg[61]), .B1(
        inner_first_stage_valid_reg[57]), .B2(n10299), .ZN(n11756) );
  INR3D2BWP30P140LVT U15054 ( .A1(inner_first_stage_valid_reg[56]), .B1(
        inner_first_stage_valid_reg[58]), .B2(n10300), .ZN(n11758) );
  INR4D1BWP30P140LVT U15055 ( .A1(n10304), .B1(inner_first_stage_valid_reg[57]), .B2(inner_first_stage_valid_reg[61]), .B3(n10303), .ZN(n11755) );
  NR4D0BWP30P140LVT U15056 ( .A1(n11756), .A2(n11758), .A3(n11757), .A4(n11755), .ZN(n10305) );
  AOI22D1BWP30P140LVT U15057 ( .A1(n10620), .A2(i_data_bus[904]), .B1(n10619), 
        .B2(i_data_bus[1000]), .ZN(n10308) );
  AOI22D1BWP30P140LVT U15058 ( .A1(n10618), .A2(i_data_bus[936]), .B1(n10617), 
        .B2(i_data_bus[968]), .ZN(n10307) );
  AOI22D1BWP30P140LVT U15059 ( .A1(n10620), .A2(i_data_bus[901]), .B1(n10619), 
        .B2(i_data_bus[997]), .ZN(n10310) );
  AOI22D1BWP30P140LVT U15060 ( .A1(n10618), .A2(i_data_bus[933]), .B1(n10617), 
        .B2(i_data_bus[965]), .ZN(n10309) );
  AOI22D1BWP30P140LVT U15061 ( .A1(n10620), .A2(i_data_bus[909]), .B1(n10618), 
        .B2(i_data_bus[941]), .ZN(n10312) );
  AOI22D1BWP30P140LVT U15062 ( .A1(n10619), .A2(i_data_bus[1005]), .B1(n10617), 
        .B2(i_data_bus[973]), .ZN(n10311) );
  AOI22D1BWP30P140LVT U15063 ( .A1(n10619), .A2(i_data_bus[1002]), .B1(n10618), 
        .B2(i_data_bus[938]), .ZN(n10314) );
  AOI22D1BWP30P140LVT U15064 ( .A1(n10620), .A2(i_data_bus[906]), .B1(n10617), 
        .B2(i_data_bus[970]), .ZN(n10313) );
  AOI22D1BWP30P140LVT U15065 ( .A1(n10620), .A2(i_data_bus[916]), .B1(n10618), 
        .B2(i_data_bus[948]), .ZN(n10316) );
  AOI22D1BWP30P140LVT U15066 ( .A1(n10619), .A2(i_data_bus[1012]), .B1(n10617), 
        .B2(i_data_bus[980]), .ZN(n10315) );
  AOI22D1BWP30P140LVT U15067 ( .A1(n10620), .A2(i_data_bus[914]), .B1(n10619), 
        .B2(i_data_bus[1010]), .ZN(n10318) );
  AOI22D1BWP30P140LVT U15068 ( .A1(n10618), .A2(i_data_bus[946]), .B1(n10617), 
        .B2(i_data_bus[978]), .ZN(n10317) );
  AOI22D1BWP30P140LVT U15069 ( .A1(n10619), .A2(i_data_bus[1020]), .B1(n10618), 
        .B2(i_data_bus[956]), .ZN(n10320) );
  AOI22D1BWP30P140LVT U15070 ( .A1(n10620), .A2(i_data_bus[924]), .B1(n10617), 
        .B2(i_data_bus[988]), .ZN(n10319) );
  AOI22D1BWP30P140LVT U15071 ( .A1(n10619), .A2(i_data_bus[1021]), .B1(n10618), 
        .B2(i_data_bus[957]), .ZN(n10322) );
  AOI22D1BWP30P140LVT U15072 ( .A1(n10620), .A2(i_data_bus[925]), .B1(n10617), 
        .B2(i_data_bus[989]), .ZN(n10321) );
  AOI22D1BWP30P140LVT U15073 ( .A1(n10620), .A2(i_data_bus[922]), .B1(n10619), 
        .B2(i_data_bus[1018]), .ZN(n10324) );
  AOI22D1BWP30P140LVT U15074 ( .A1(n10618), .A2(i_data_bus[954]), .B1(n10617), 
        .B2(i_data_bus[986]), .ZN(n10323) );
  AOI22D1BWP30P140LVT U15075 ( .A1(n10619), .A2(i_data_bus[1017]), .B1(n10618), 
        .B2(i_data_bus[953]), .ZN(n10326) );
  AOI22D1BWP30P140LVT U15076 ( .A1(n10620), .A2(i_data_bus[921]), .B1(n10617), 
        .B2(i_data_bus[985]), .ZN(n10325) );
  AOI22D1BWP30P140LVT U15077 ( .A1(n10620), .A2(i_data_bus[905]), .B1(n10618), 
        .B2(i_data_bus[937]), .ZN(n10328) );
  AOI22D1BWP30P140LVT U15078 ( .A1(n10619), .A2(i_data_bus[1001]), .B1(n10617), 
        .B2(i_data_bus[969]), .ZN(n10327) );
  AOI22D1BWP30P140LVT U15079 ( .A1(n10619), .A2(i_data_bus[1013]), .B1(n10618), 
        .B2(i_data_bus[949]), .ZN(n10330) );
  AOI22D1BWP30P140LVT U15080 ( .A1(n10620), .A2(i_data_bus[917]), .B1(n10617), 
        .B2(i_data_bus[981]), .ZN(n10329) );
  AOI22D1BWP30P140LVT U15081 ( .A1(n10619), .A2(i_data_bus[994]), .B1(n10618), 
        .B2(i_data_bus[930]), .ZN(n10332) );
  AOI22D1BWP30P140LVT U15082 ( .A1(n10620), .A2(i_data_bus[898]), .B1(n10617), 
        .B2(i_data_bus[962]), .ZN(n10331) );
  NR3D0P7BWP30P140LVT U15083 ( .A1(inner_first_stage_valid_reg[8]), .A2(
        inner_first_stage_valid_reg[14]), .A3(inner_first_stage_valid_reg[15]), 
        .ZN(n10338) );
  NR2D1BWP30P140LVT U15084 ( .A1(inner_first_stage_valid_reg[9]), .A2(
        inner_first_stage_valid_reg[13]), .ZN(n10333) );
  INR3D2BWP30P140LVT U15085 ( .A1(inner_first_stage_valid_reg[11]), .B1(
        inner_first_stage_valid_reg[10]), .B2(n10337), .ZN(n10944) );
  NR2D1BWP30P140LVT U15086 ( .A1(inner_first_stage_valid_reg[8]), .A2(
        inner_first_stage_valid_reg[13]), .ZN(n10339) );
  NR3D0P7BWP30P140LVT U15087 ( .A1(inner_first_stage_valid_reg[10]), .A2(
        inner_first_stage_valid_reg[11]), .A3(inner_first_stage_valid_reg[9]), 
        .ZN(n10334) );
  ND3D1BWP30P140LVT U15088 ( .A1(n10339), .A2(n10335), .A3(n10334), .ZN(n10336) );
  INR3D2BWP30P140LVT U15089 ( .A1(inner_first_stage_valid_reg[15]), .B1(
        inner_first_stage_valid_reg[14]), .B2(n10336), .ZN(n10946) );
  INR3D2BWP30P140LVT U15090 ( .A1(inner_first_stage_valid_reg[14]), .B1(
        inner_first_stage_valid_reg[15]), .B2(n10336), .ZN(n10943) );
  INR3D2BWP30P140LVT U15091 ( .A1(inner_first_stage_valid_reg[10]), .B1(
        inner_first_stage_valid_reg[11]), .B2(n10337), .ZN(n10945) );
  NR4D0BWP30P140LVT U15092 ( .A1(n10944), .A2(n10946), .A3(n10943), .A4(n10945), .ZN(n10346) );
  NR4D0BWP30P140LVT U15093 ( .A1(inner_first_stage_valid_reg[10]), .A2(
        inner_first_stage_valid_reg[11]), .A3(inner_first_stage_valid_reg[9]), 
        .A4(inner_first_stage_valid_reg[13]), .ZN(n10341) );
  NR2D1BWP30P140LVT U15094 ( .A1(inner_first_stage_valid_reg[10]), .A2(
        inner_first_stage_valid_reg[11]), .ZN(n10342) );
  NR4D0BWP30P140LVT U15095 ( .A1(inner_first_stage_valid_reg[14]), .A2(
        inner_first_stage_valid_reg[12]), .A3(inner_first_stage_valid_reg[15]), 
        .A4(n10380), .ZN(n10340) );
  INVD1BWP30P140LVT U15096 ( .I(n10342), .ZN(n10344) );
  INR4D1BWP30P140LVT U15097 ( .A1(inner_first_stage_valid_reg[13]), .B1(n10344), .B2(inner_first_stage_valid_reg[9]), .B3(n10343), .ZN(n10941) );
  NR4D0BWP30P140LVT U15098 ( .A1(n10940), .A2(n10939), .A3(n10942), .A4(n10941), .ZN(n10345) );
  ND2D1BWP30P140LVT U15099 ( .A1(n10346), .A2(n10345), .ZN(N4102) );
  INVD1BWP30P140LVT U15100 ( .I(inner_first_stage_valid_reg[41]), .ZN(n10349)
         );
  INVD1BWP30P140LVT U15101 ( .I(inner_first_stage_valid_reg[45]), .ZN(n10355)
         );
  ND4D1BWP30P140LVT U15102 ( .A1(n10349), .A2(n10355), .A3(n10347), .A4(n10352), .ZN(n10357) );
  INR3D2BWP30P140LVT U15103 ( .A1(inner_first_stage_valid_reg[46]), .B1(
        inner_first_stage_valid_reg[47]), .B2(n10356), .ZN(n11488) );
  NR4D0BWP30P140LVT U15104 ( .A1(inner_first_stage_valid_reg[44]), .A2(
        inner_first_stage_valid_reg[47]), .A3(inner_first_stage_valid_reg[46]), 
        .A4(n10359), .ZN(n10348) );
  NR3D0P7BWP30P140LVT U15105 ( .A1(inner_first_stage_valid_reg[44]), .A2(
        inner_first_stage_valid_reg[47]), .A3(inner_first_stage_valid_reg[46]), 
        .ZN(n10351) );
  NR2D1BWP30P140LVT U15106 ( .A1(inner_first_stage_valid_reg[41]), .A2(
        inner_first_stage_valid_reg[45]), .ZN(n10350) );
  ND2D1BWP30P140LVT U15107 ( .A1(n10351), .A2(n10350), .ZN(n10358) );
  INR3D2BWP30P140LVT U15108 ( .A1(inner_first_stage_valid_reg[42]), .B1(
        inner_first_stage_valid_reg[43]), .B2(n10353), .ZN(n11489) );
  NR4D0BWP30P140LVT U15109 ( .A1(n11488), .A2(n11487), .A3(n11490), .A4(n11489), .ZN(n10362) );
  INR3D2BWP30P140LVT U15110 ( .A1(inner_first_stage_valid_reg[47]), .B1(
        inner_first_stage_valid_reg[46]), .B2(n10356), .ZN(n11484) );
  INR4D1BWP30P140LVT U15111 ( .A1(inner_first_stage_valid_reg[44]), .B1(
        inner_first_stage_valid_reg[46]), .B2(inner_first_stage_valid_reg[47]), 
        .B3(n10357), .ZN(n11485) );
  NR4D0BWP30P140LVT U15112 ( .A1(n11486), .A2(n11484), .A3(n11485), .A4(n5893), 
        .ZN(n10361) );
  INVD1BWP30P140LVT U15113 ( .I(inner_first_stage_valid_reg[16]), .ZN(n10364)
         );
  ND3D1BWP30P140LVT U15114 ( .A1(n11767), .A2(n10368), .A3(n5900), .ZN(n10369)
         );
  NR3D0P7BWP30P140LVT U15115 ( .A1(inner_first_stage_valid_reg[22]), .A2(
        inner_first_stage_valid_reg[23]), .A3(inner_first_stage_valid_reg[20]), 
        .ZN(n10365) );
  NR4D1BWP30P140LVT U15116 ( .A1(inner_first_stage_valid_reg[17]), .A2(
        inner_first_stage_valid_reg[21]), .A3(n10364), .A4(n10363), .ZN(n11080) );
  INR4D1BWP30P140LVT U15117 ( .A1(inner_first_stage_valid_reg[21]), .B1(
        inner_first_stage_valid_reg[16]), .B2(inner_first_stage_valid_reg[17]), 
        .B3(n10363), .ZN(n11079) );
  NR2D1BWP30P140LVT U15118 ( .A1(inner_first_stage_valid_reg[21]), .A2(
        inner_first_stage_valid_reg[17]), .ZN(n10366) );
  ND4D1BWP30P140LVT U15119 ( .A1(n5900), .A2(n10366), .A3(n10365), .A4(n10364), 
        .ZN(n10367) );
  NR4D0BWP30P140LVT U15120 ( .A1(n11080), .A2(n11079), .A3(n11082), .A4(n11081), .ZN(n10377) );
  INVD1BWP30P140LVT U15121 ( .I(inner_first_stage_valid_reg[17]), .ZN(n10373)
         );
  NR2D1BWP30P140LVT U15122 ( .A1(inner_first_stage_valid_reg[22]), .A2(
        inner_first_stage_valid_reg[23]), .ZN(n10370) );
  NR3D0P7BWP30P140LVT U15123 ( .A1(inner_first_stage_valid_reg[16]), .A2(
        inner_first_stage_valid_reg[21]), .A3(n10369), .ZN(n10374) );
  INVD1BWP30P140LVT U15124 ( .I(inner_first_stage_valid_reg[20]), .ZN(n10372)
         );
  ND3D1BWP30P140LVT U15125 ( .A1(n10374), .A2(n10373), .A3(n10372), .ZN(n10375) );
  INR3D2BWP30P140LVT U15126 ( .A1(inner_first_stage_valid_reg[22]), .B1(
        inner_first_stage_valid_reg[23]), .B2(n10375), .ZN(n11078) );
  INR3D2BWP30P140LVT U15127 ( .A1(inner_first_stage_valid_reg[23]), .B1(
        inner_first_stage_valid_reg[22]), .B2(n10375), .ZN(n11077) );
  NR4D0BWP30P140LVT U15128 ( .A1(n11076), .A2(n11075), .A3(n11078), .A4(n11077), .ZN(n10376) );
  INVD1BWP30P140LVT U15129 ( .I(inner_first_stage_valid_reg[27]), .ZN(n10379)
         );
  NR2D1BWP30P140LVT U15130 ( .A1(inner_first_stage_valid_reg[25]), .A2(
        inner_first_stage_valid_reg[29]), .ZN(n10378) );
  NR3D0P7BWP30P140LVT U15131 ( .A1(inner_first_stage_valid_reg[30]), .A2(
        inner_first_stage_valid_reg[31]), .A3(n10380), .ZN(n10388) );
  INVD1BWP30P140LVT U15132 ( .I(inner_first_stage_valid_reg[24]), .ZN(n10385)
         );
  IND4D1BWP30P140LVT U15133 ( .A1(inner_first_stage_valid_reg[28]), .B1(n10378), .B2(n10388), .B3(n10385), .ZN(n10389) );
  INVD1BWP30P140LVT U15134 ( .I(inner_first_stage_valid_reg[26]), .ZN(n10390)
         );
  NR2D1BWP30P140LVT U15135 ( .A1(inner_first_stage_valid_reg[30]), .A2(
        inner_first_stage_valid_reg[31]), .ZN(n10381) );
  IND3D1BWP30P140LVT U15136 ( .A1(n10382), .B1(n10381), .B2(n10383), .ZN(
        n10386) );
  INR4D1BWP30P140LVT U15137 ( .A1(inner_first_stage_valid_reg[29]), .B1(
        inner_first_stage_valid_reg[24]), .B2(inner_first_stage_valid_reg[25]), 
        .B3(n10386), .ZN(n11215) );
  NR4D0BWP30P140LVT U15138 ( .A1(inner_first_stage_valid_reg[24]), .A2(
        inner_first_stage_valid_reg[25]), .A3(inner_first_stage_valid_reg[29]), 
        .A4(n10382), .ZN(n10387) );
  INR3D2BWP30P140LVT U15139 ( .A1(inner_first_stage_valid_reg[31]), .B1(
        inner_first_stage_valid_reg[30]), .B2(n10384), .ZN(n11218) );
  INR3D2BWP30P140LVT U15140 ( .A1(inner_first_stage_valid_reg[30]), .B1(
        inner_first_stage_valid_reg[31]), .B2(n10384), .ZN(n11217) );
  NR4D0BWP30P140LVT U15141 ( .A1(n11216), .A2(n11215), .A3(n11218), .A4(n11217), .ZN(n10392) );
  INR4D1BWP30P140LVT U15142 ( .A1(inner_first_stage_valid_reg[25]), .B1(
        inner_first_stage_valid_reg[24]), .B2(inner_first_stage_valid_reg[29]), 
        .B3(n10386), .ZN(n11213) );
  NR4D0BWP30P140LVT U15143 ( .A1(n11214), .A2(n11213), .A3(n11212), .A4(n11211), .ZN(n10391) );
  ND2D1BWP30P140LVT U15144 ( .A1(n10392), .A2(n10391), .ZN(N7850) );
  OR4D1BWP30P140LVT U15145 ( .A1(n10396), .A2(n10395), .A3(n10394), .A4(n10393), .Z(N15200) );
  OR4D1BWP30P140LVT U15146 ( .A1(n10400), .A2(n10399), .A3(n10398), .A4(n10397), .Z(N14984) );
  OR4D1BWP30P140LVT U15147 ( .A1(n10404), .A2(n10403), .A3(n10402), .A4(n10401), .Z(N14768) );
  OR4D1BWP30P140LVT U15148 ( .A1(n10408), .A2(n10407), .A3(n10406), .A4(n10405), .Z(N14552) );
  OR4D1BWP30P140LVT U15149 ( .A1(n10412), .A2(n10411), .A3(n10410), .A4(n10409), .Z(N14336) );
  OR4D1BWP30P140LVT U15150 ( .A1(n10416), .A2(n10415), .A3(n10414), .A4(n10413), .Z(N14120) );
  OR4D1BWP30P140LVT U15151 ( .A1(n10420), .A2(n10419), .A3(n10418), .A4(n10417), .Z(N13904) );
  OR4D1BWP30P140LVT U15152 ( .A1(n10424), .A2(n10423), .A3(n10422), .A4(n10421), .Z(N13688) );
  OR4D1BWP30P140LVT U15153 ( .A1(n10428), .A2(n10427), .A3(n10426), .A4(n10425), .Z(N13326) );
  OR4D1BWP30P140LVT U15154 ( .A1(n10432), .A2(n10431), .A3(n10430), .A4(n10429), .Z(N13110) );
  OR4D1BWP30P140LVT U15155 ( .A1(n10436), .A2(n10435), .A3(n10434), .A4(n10433), .Z(N12894) );
  OR4D1BWP30P140LVT U15156 ( .A1(n10440), .A2(n10439), .A3(n10438), .A4(n10437), .Z(N12678) );
  OR4D1BWP30P140LVT U15157 ( .A1(n10444), .A2(n10443), .A3(n10442), .A4(n10441), .Z(N12462) );
  OR4D1BWP30P140LVT U15158 ( .A1(n10448), .A2(n10447), .A3(n10446), .A4(n10445), .Z(N12246) );
  OR4D1BWP30P140LVT U15159 ( .A1(n10452), .A2(n10451), .A3(n10450), .A4(n10449), .Z(N12030) );
  OR4D1BWP30P140LVT U15160 ( .A1(n10456), .A2(n10455), .A3(n10454), .A4(n10453), .Z(N11814) );
  OR4D1BWP30P140LVT U15161 ( .A1(n10460), .A2(n10459), .A3(n10458), .A4(n10457), .Z(N11452) );
  OR4D1BWP30P140LVT U15162 ( .A1(n10464), .A2(n10463), .A3(n10462), .A4(n10461), .Z(N11236) );
  OR4D1BWP30P140LVT U15163 ( .A1(n10468), .A2(n10467), .A3(n10466), .A4(n10465), .Z(N11020) );
  OR4D1BWP30P140LVT U15164 ( .A1(n10472), .A2(n10471), .A3(n10470), .A4(n10469), .Z(N10804) );
  OR4D1BWP30P140LVT U15165 ( .A1(n10476), .A2(n10475), .A3(n10474), .A4(n10473), .Z(N10588) );
  OR4D1BWP30P140LVT U15166 ( .A1(n10480), .A2(n10479), .A3(n10478), .A4(n10477), .Z(N10372) );
  OR4D1BWP30P140LVT U15167 ( .A1(n10484), .A2(n10483), .A3(n10482), .A4(n10481), .Z(N10156) );
  OR4D1BWP30P140LVT U15168 ( .A1(n10488), .A2(n10487), .A3(n10486), .A4(n10485), .Z(N9940) );
  OR4D1BWP30P140LVT U15169 ( .A1(n10492), .A2(n10491), .A3(n10490), .A4(n10489), .Z(N9578) );
  OR4D1BWP30P140LVT U15170 ( .A1(n10496), .A2(n10495), .A3(n10494), .A4(n10493), .Z(N9362) );
  OR4D1BWP30P140LVT U15171 ( .A1(n10500), .A2(n10499), .A3(n10498), .A4(n10497), .Z(N9146) );
  OR4D1BWP30P140LVT U15172 ( .A1(n10504), .A2(n10503), .A3(n10502), .A4(n10501), .Z(N8930) );
  OR4D1BWP30P140LVT U15173 ( .A1(n10508), .A2(n10507), .A3(n10506), .A4(n10505), .Z(N8714) );
  OR4D1BWP30P140LVT U15174 ( .A1(n10512), .A2(n10511), .A3(n10510), .A4(n10509), .Z(N8498) );
  OR4D1BWP30P140LVT U15175 ( .A1(n10516), .A2(n10515), .A3(n10514), .A4(n10513), .Z(N8282) );
  OR4D1BWP30P140LVT U15176 ( .A1(n10520), .A2(n10519), .A3(n10518), .A4(n10517), .Z(N8066) );
  OR4D1BWP30P140LVT U15177 ( .A1(n10524), .A2(n10523), .A3(n10522), .A4(n10521), .Z(N7704) );
  OR4D1BWP30P140LVT U15178 ( .A1(n10528), .A2(n10527), .A3(n10526), .A4(n10525), .Z(N7488) );
  OR4D1BWP30P140LVT U15179 ( .A1(n10532), .A2(n10531), .A3(n10530), .A4(n10529), .Z(N7272) );
  OR4D1BWP30P140LVT U15180 ( .A1(n10536), .A2(n10535), .A3(n10534), .A4(n10533), .Z(N7056) );
  OR4D1BWP30P140LVT U15181 ( .A1(n10540), .A2(n10539), .A3(n10538), .A4(n10537), .Z(N6840) );
  OR4D1BWP30P140LVT U15182 ( .A1(n10544), .A2(n10543), .A3(n10542), .A4(n10541), .Z(N6624) );
  OR4D1BWP30P140LVT U15183 ( .A1(n10548), .A2(n10547), .A3(n10546), .A4(n10545), .Z(N6408) );
  OR4D1BWP30P140LVT U15184 ( .A1(n10552), .A2(n10551), .A3(n10550), .A4(n10549), .Z(N6192) );
  OR4D1BWP30P140LVT U15185 ( .A1(n10556), .A2(n10555), .A3(n10554), .A4(n10553), .Z(N5830) );
  OR4D1BWP30P140LVT U15186 ( .A1(n10560), .A2(n10559), .A3(n10558), .A4(n10557), .Z(N5614) );
  OR4D1BWP30P140LVT U15187 ( .A1(n10564), .A2(n10563), .A3(n10562), .A4(n10561), .Z(N5398) );
  OR4D1BWP30P140LVT U15188 ( .A1(n10568), .A2(n10567), .A3(n10566), .A4(n10565), .Z(N5182) );
  OR4D1BWP30P140LVT U15189 ( .A1(n10572), .A2(n10571), .A3(n10570), .A4(n10569), .Z(N4966) );
  OR4D1BWP30P140LVT U15190 ( .A1(n10576), .A2(n10575), .A3(n10574), .A4(n10573), .Z(N4750) );
  OR4D1BWP30P140LVT U15191 ( .A1(n10580), .A2(n10579), .A3(n10578), .A4(n10577), .Z(N4534) );
  OR4D1BWP30P140LVT U15192 ( .A1(n10584), .A2(n10583), .A3(n10582), .A4(n10581), .Z(N4318) );
  OR4D1BWP30P140LVT U15193 ( .A1(n10588), .A2(n10587), .A3(n10586), .A4(n10585), .Z(N3956) );
  OR4D1BWP30P140LVT U15194 ( .A1(n10592), .A2(n10591), .A3(n10590), .A4(n10589), .Z(N3740) );
  OR4D1BWP30P140LVT U15195 ( .A1(n10596), .A2(n10595), .A3(n10594), .A4(n10593), .Z(N3524) );
  OR4D1BWP30P140LVT U15196 ( .A1(n10600), .A2(n10599), .A3(n10598), .A4(n10597), .Z(N3308) );
  OR4D1BWP30P140LVT U15197 ( .A1(n10604), .A2(n10603), .A3(n10602), .A4(n10601), .Z(N3092) );
  OR4D1BWP30P140LVT U15198 ( .A1(n10608), .A2(n10607), .A3(n10606), .A4(n10605), .Z(N2876) );
  OR4D1BWP30P140LVT U15199 ( .A1(n10612), .A2(n10611), .A3(n10610), .A4(n10609), .Z(N2660) );
  OR4D1BWP30P140LVT U15200 ( .A1(n10616), .A2(n10615), .A3(n10614), .A4(n10613), .Z(N2444) );
  OR4D1BWP30P140LVT U15201 ( .A1(n10620), .A2(n10619), .A3(n10618), .A4(n10617), .Z(N2082) );
  OR4D1BWP30P140LVT U15202 ( .A1(n10623), .A2(n10622), .A3(n10621), .A4(n9749), 
        .Z(N1862) );
  OR4D1BWP30P140LVT U15203 ( .A1(n10627), .A2(n10626), .A3(n10625), .A4(n10624), .Z(N1642) );
  OR4D1BWP30P140LVT U15204 ( .A1(n10631), .A2(n10630), .A3(n10629), .A4(n10628), .Z(N1422) );
  OR4D1BWP30P140LVT U15205 ( .A1(n10634), .A2(n10633), .A3(n10632), .A4(n9766), 
        .Z(N1202) );
  OR4D1BWP30P140LVT U15206 ( .A1(n10638), .A2(n10637), .A3(n10636), .A4(n10635), .Z(N982) );
  OR4D1BWP30P140LVT U15207 ( .A1(n10642), .A2(n10641), .A3(n10640), .A4(n10639), .Z(N762) );
  OR4D1BWP30P140LVT U15208 ( .A1(n10646), .A2(n10645), .A3(n10644), .A4(n10643), .Z(N542) );
  AOI22D1BWP30P140LVT U15209 ( .A1(n10803), .A2(
        inner_first_stage_data_reg[160]), .B1(n10802), .B2(
        inner_first_stage_data_reg[192]), .ZN(n10650) );
  AOI22D1BWP30P140LVT U15210 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[224]), .B1(n10808), .B2(
        inner_first_stage_data_reg[0]), .ZN(n10649) );
  AOI22D1BWP30P140LVT U15211 ( .A1(n10806), .A2(inner_first_stage_data_reg[96]), .B1(n10804), .B2(inner_first_stage_data_reg[128]), .ZN(n10648) );
  ND2D1BWP30P140LVT U15212 ( .A1(n10807), .A2(inner_first_stage_data_reg[32]), 
        .ZN(n10647) );
  ND4D1BWP30P140LVT U15213 ( .A1(n10650), .A2(n10649), .A3(n10648), .A4(n10647), .ZN(n10651) );
  AO21D1BWP30P140LVT U15214 ( .A1(n10814), .A2(inner_first_stage_data_reg[64]), 
        .B(n10651), .Z(N2229) );
  AOI22D1BWP30P140LVT U15215 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[225]), .B1(n10802), .B2(
        inner_first_stage_data_reg[193]), .ZN(n10655) );
  AOI22D1BWP30P140LVT U15216 ( .A1(n10803), .A2(
        inner_first_stage_data_reg[161]), .B1(n10807), .B2(
        inner_first_stage_data_reg[33]), .ZN(n10654) );
  AOI22D1BWP30P140LVT U15217 ( .A1(n10814), .A2(inner_first_stage_data_reg[65]), .B1(n10804), .B2(inner_first_stage_data_reg[129]), .ZN(n10653) );
  ND2D1BWP30P140LVT U15218 ( .A1(n10808), .A2(inner_first_stage_data_reg[1]), 
        .ZN(n10652) );
  ND4D1BWP30P140LVT U15219 ( .A1(n10655), .A2(n10654), .A3(n10653), .A4(n10652), .ZN(n10656) );
  AO21D1BWP30P140LVT U15220 ( .A1(n10806), .A2(inner_first_stage_data_reg[97]), 
        .B(n10656), .Z(N2230) );
  AOI22D1BWP30P140LVT U15221 ( .A1(n10803), .A2(
        inner_first_stage_data_reg[162]), .B1(n10802), .B2(
        inner_first_stage_data_reg[194]), .ZN(n10660) );
  AOI22D1BWP30P140LVT U15222 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[226]), .B1(n10807), .B2(
        inner_first_stage_data_reg[34]), .ZN(n10659) );
  AOI22D1BWP30P140LVT U15223 ( .A1(n10808), .A2(inner_first_stage_data_reg[2]), 
        .B1(n10804), .B2(inner_first_stage_data_reg[130]), .ZN(n10658) );
  ND2D1BWP30P140LVT U15224 ( .A1(n10806), .A2(inner_first_stage_data_reg[98]), 
        .ZN(n10657) );
  ND4D1BWP30P140LVT U15225 ( .A1(n10660), .A2(n10659), .A3(n10658), .A4(n10657), .ZN(n10661) );
  AO21D1BWP30P140LVT U15226 ( .A1(n10814), .A2(inner_first_stage_data_reg[66]), 
        .B(n10661), .Z(N2231) );
  AOI22D1BWP30P140LVT U15227 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[227]), .B1(n10803), .B2(
        inner_first_stage_data_reg[163]), .ZN(n10665) );
  AOI22D1BWP30P140LVT U15228 ( .A1(n10802), .A2(
        inner_first_stage_data_reg[195]), .B1(n10807), .B2(
        inner_first_stage_data_reg[35]), .ZN(n10664) );
  AOI22D1BWP30P140LVT U15229 ( .A1(n10808), .A2(inner_first_stage_data_reg[3]), 
        .B1(n10806), .B2(inner_first_stage_data_reg[99]), .ZN(n10663) );
  ND2D1BWP30P140LVT U15230 ( .A1(n10804), .A2(inner_first_stage_data_reg[131]), 
        .ZN(n10662) );
  ND4D1BWP30P140LVT U15231 ( .A1(n10665), .A2(n10664), .A3(n10663), .A4(n10662), .ZN(n10666) );
  AO21D1BWP30P140LVT U15232 ( .A1(n10814), .A2(inner_first_stage_data_reg[67]), 
        .B(n10666), .Z(N2232) );
  AOI22D1BWP30P140LVT U15233 ( .A1(n10803), .A2(
        inner_first_stage_data_reg[164]), .B1(n10802), .B2(
        inner_first_stage_data_reg[196]), .ZN(n10670) );
  AOI22D1BWP30P140LVT U15234 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[228]), .B1(n10808), .B2(
        inner_first_stage_data_reg[4]), .ZN(n10669) );
  AOI22D1BWP30P140LVT U15235 ( .A1(n10807), .A2(inner_first_stage_data_reg[36]), .B1(n10804), .B2(inner_first_stage_data_reg[132]), .ZN(n10668) );
  ND2D1BWP30P140LVT U15236 ( .A1(n10814), .A2(inner_first_stage_data_reg[68]), 
        .ZN(n10667) );
  ND4D1BWP30P140LVT U15237 ( .A1(n10670), .A2(n10669), .A3(n10668), .A4(n10667), .ZN(n10671) );
  AO21D1BWP30P140LVT U15238 ( .A1(n10806), .A2(inner_first_stage_data_reg[100]), .B(n10671), .Z(N2233) );
  AOI22D1BWP30P140LVT U15239 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[229]), .B1(n10803), .B2(
        inner_first_stage_data_reg[165]), .ZN(n10675) );
  AOI22D1BWP30P140LVT U15240 ( .A1(n10802), .A2(
        inner_first_stage_data_reg[197]), .B1(n10804), .B2(
        inner_first_stage_data_reg[133]), .ZN(n10674) );
  AOI22D1BWP30P140LVT U15241 ( .A1(n10808), .A2(inner_first_stage_data_reg[5]), 
        .B1(n10807), .B2(inner_first_stage_data_reg[37]), .ZN(n10673) );
  ND2D1BWP30P140LVT U15242 ( .A1(n10814), .A2(inner_first_stage_data_reg[69]), 
        .ZN(n10672) );
  ND4D1BWP30P140LVT U15243 ( .A1(n10675), .A2(n10674), .A3(n10673), .A4(n10672), .ZN(n10676) );
  AO21D1BWP30P140LVT U15244 ( .A1(n10806), .A2(inner_first_stage_data_reg[101]), .B(n10676), .Z(N2234) );
  AOI22D1BWP30P140LVT U15245 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[230]), .B1(n10803), .B2(
        inner_first_stage_data_reg[166]), .ZN(n10680) );
  AOI22D1BWP30P140LVT U15246 ( .A1(n10802), .A2(
        inner_first_stage_data_reg[198]), .B1(n10804), .B2(
        inner_first_stage_data_reg[134]), .ZN(n10679) );
  AOI22D1BWP30P140LVT U15247 ( .A1(n10814), .A2(inner_first_stage_data_reg[70]), .B1(n10807), .B2(inner_first_stage_data_reg[38]), .ZN(n10678) );
  ND2D1BWP30P140LVT U15248 ( .A1(n10808), .A2(inner_first_stage_data_reg[6]), 
        .ZN(n10677) );
  ND4D1BWP30P140LVT U15249 ( .A1(n10680), .A2(n10679), .A3(n10678), .A4(n10677), .ZN(n10681) );
  AO21D1BWP30P140LVT U15250 ( .A1(n10806), .A2(inner_first_stage_data_reg[102]), .B(n10681), .Z(N2235) );
  AOI22D1BWP30P140LVT U15251 ( .A1(n10803), .A2(
        inner_first_stage_data_reg[167]), .B1(n10802), .B2(
        inner_first_stage_data_reg[199]), .ZN(n10685) );
  AOI22D1BWP30P140LVT U15252 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[231]), .B1(n10804), .B2(
        inner_first_stage_data_reg[135]), .ZN(n10684) );
  AOI22D1BWP30P140LVT U15253 ( .A1(n10808), .A2(inner_first_stage_data_reg[7]), 
        .B1(n10807), .B2(inner_first_stage_data_reg[39]), .ZN(n10683) );
  ND2D1BWP30P140LVT U15254 ( .A1(n10806), .A2(inner_first_stage_data_reg[103]), 
        .ZN(n10682) );
  ND4D1BWP30P140LVT U15255 ( .A1(n10685), .A2(n10684), .A3(n10683), .A4(n10682), .ZN(n10686) );
  AO21D1BWP30P140LVT U15256 ( .A1(n10814), .A2(inner_first_stage_data_reg[71]), 
        .B(n10686), .Z(N2236) );
  AOI22D1BWP30P140LVT U15257 ( .A1(n10803), .A2(
        inner_first_stage_data_reg[168]), .B1(n10802), .B2(
        inner_first_stage_data_reg[200]), .ZN(n10690) );
  AOI22D1BWP30P140LVT U15258 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[232]), .B1(n10808), .B2(
        inner_first_stage_data_reg[8]), .ZN(n10689) );
  AOI22D1BWP30P140LVT U15259 ( .A1(n10807), .A2(inner_first_stage_data_reg[40]), .B1(n10804), .B2(inner_first_stage_data_reg[136]), .ZN(n10688) );
  ND2D1BWP30P140LVT U15260 ( .A1(n10814), .A2(inner_first_stage_data_reg[72]), 
        .ZN(n10687) );
  ND4D1BWP30P140LVT U15261 ( .A1(n10690), .A2(n10689), .A3(n10688), .A4(n10687), .ZN(n10691) );
  AO21D1BWP30P140LVT U15262 ( .A1(n10806), .A2(inner_first_stage_data_reg[104]), .B(n10691), .Z(N2237) );
  AOI22D1BWP30P140LVT U15263 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[233]), .B1(n10802), .B2(
        inner_first_stage_data_reg[201]), .ZN(n10695) );
  AOI22D1BWP30P140LVT U15264 ( .A1(n10803), .A2(
        inner_first_stage_data_reg[169]), .B1(n10807), .B2(
        inner_first_stage_data_reg[41]), .ZN(n10694) );
  AOI22D1BWP30P140LVT U15265 ( .A1(n10814), .A2(inner_first_stage_data_reg[73]), .B1(n10808), .B2(inner_first_stage_data_reg[9]), .ZN(n10693) );
  ND2D1BWP30P140LVT U15266 ( .A1(n10804), .A2(inner_first_stage_data_reg[137]), 
        .ZN(n10692) );
  ND4D1BWP30P140LVT U15267 ( .A1(n10695), .A2(n10694), .A3(n10693), .A4(n10692), .ZN(n10696) );
  AO21D1BWP30P140LVT U15268 ( .A1(n10806), .A2(inner_first_stage_data_reg[105]), .B(n10696), .Z(N2238) );
  AOI22D1BWP30P140LVT U15269 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[234]), .B1(n10802), .B2(
        inner_first_stage_data_reg[202]), .ZN(n10700) );
  AOI22D1BWP30P140LVT U15270 ( .A1(n10803), .A2(
        inner_first_stage_data_reg[170]), .B1(n10807), .B2(
        inner_first_stage_data_reg[42]), .ZN(n10699) );
  AOI22D1BWP30P140LVT U15271 ( .A1(n10814), .A2(inner_first_stage_data_reg[74]), .B1(n10804), .B2(inner_first_stage_data_reg[138]), .ZN(n10698) );
  ND2D1BWP30P140LVT U15272 ( .A1(n10808), .A2(inner_first_stage_data_reg[10]), 
        .ZN(n10697) );
  ND4D1BWP30P140LVT U15273 ( .A1(n10700), .A2(n10699), .A3(n10698), .A4(n10697), .ZN(n10701) );
  AO21D1BWP30P140LVT U15274 ( .A1(n10806), .A2(inner_first_stage_data_reg[106]), .B(n10701), .Z(N2239) );
  AOI22D1BWP30P140LVT U15275 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[235]), .B1(n10802), .B2(
        inner_first_stage_data_reg[203]), .ZN(n10705) );
  AOI22D1BWP30P140LVT U15276 ( .A1(n10803), .A2(
        inner_first_stage_data_reg[171]), .B1(n10807), .B2(
        inner_first_stage_data_reg[43]), .ZN(n10704) );
  AOI22D1BWP30P140LVT U15277 ( .A1(n10808), .A2(inner_first_stage_data_reg[11]), .B1(n10806), .B2(inner_first_stage_data_reg[107]), .ZN(n10703) );
  ND2D1BWP30P140LVT U15278 ( .A1(n10804), .A2(inner_first_stage_data_reg[139]), 
        .ZN(n10702) );
  ND4D1BWP30P140LVT U15279 ( .A1(n10705), .A2(n10704), .A3(n10703), .A4(n10702), .ZN(n10706) );
  AO21D1BWP30P140LVT U15280 ( .A1(n10814), .A2(inner_first_stage_data_reg[75]), 
        .B(n10706), .Z(N2240) );
  AOI22D1BWP30P140LVT U15281 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[236]), .B1(n10802), .B2(
        inner_first_stage_data_reg[204]), .ZN(n10710) );
  AOI22D1BWP30P140LVT U15282 ( .A1(n10808), .A2(inner_first_stage_data_reg[12]), .B1(n10803), .B2(inner_first_stage_data_reg[172]), .ZN(n10709) );
  AOI22D1BWP30P140LVT U15283 ( .A1(n10807), .A2(inner_first_stage_data_reg[44]), .B1(n10804), .B2(inner_first_stage_data_reg[140]), .ZN(n10708) );
  ND2D1BWP30P140LVT U15284 ( .A1(n10806), .A2(inner_first_stage_data_reg[108]), 
        .ZN(n10707) );
  ND4D1BWP30P140LVT U15285 ( .A1(n10710), .A2(n10709), .A3(n10708), .A4(n10707), .ZN(n10711) );
  AO21D1BWP30P140LVT U15286 ( .A1(n10814), .A2(inner_first_stage_data_reg[76]), 
        .B(n10711), .Z(N2241) );
  AOI22D1BWP30P140LVT U15287 ( .A1(n10803), .A2(
        inner_first_stage_data_reg[173]), .B1(n10802), .B2(
        inner_first_stage_data_reg[205]), .ZN(n10715) );
  AOI22D1BWP30P140LVT U15288 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[237]), .B1(n10808), .B2(
        inner_first_stage_data_reg[13]), .ZN(n10714) );
  AOI22D1BWP30P140LVT U15289 ( .A1(n10806), .A2(
        inner_first_stage_data_reg[109]), .B1(n10804), .B2(
        inner_first_stage_data_reg[141]), .ZN(n10713) );
  ND2D1BWP30P140LVT U15290 ( .A1(n10807), .A2(inner_first_stage_data_reg[45]), 
        .ZN(n10712) );
  ND4D1BWP30P140LVT U15291 ( .A1(n10715), .A2(n10714), .A3(n10713), .A4(n10712), .ZN(n10716) );
  AO21D1BWP30P140LVT U15292 ( .A1(n10814), .A2(inner_first_stage_data_reg[77]), 
        .B(n10716), .Z(N2242) );
  AOI22D1BWP30P140LVT U15293 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[238]), .B1(n10802), .B2(
        inner_first_stage_data_reg[206]), .ZN(n10720) );
  AOI22D1BWP30P140LVT U15294 ( .A1(n10803), .A2(
        inner_first_stage_data_reg[174]), .B1(n10804), .B2(
        inner_first_stage_data_reg[142]), .ZN(n10719) );
  AOI22D1BWP30P140LVT U15295 ( .A1(n10814), .A2(inner_first_stage_data_reg[78]), .B1(n10808), .B2(inner_first_stage_data_reg[14]), .ZN(n10718) );
  ND2D1BWP30P140LVT U15296 ( .A1(n10807), .A2(inner_first_stage_data_reg[46]), 
        .ZN(n10717) );
  ND4D1BWP30P140LVT U15297 ( .A1(n10720), .A2(n10719), .A3(n10718), .A4(n10717), .ZN(n10721) );
  AO21D1BWP30P140LVT U15298 ( .A1(n10806), .A2(inner_first_stage_data_reg[110]), .B(n10721), .Z(N2243) );
  AOI22D1BWP30P140LVT U15299 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[239]), .B1(n10802), .B2(
        inner_first_stage_data_reg[207]), .ZN(n10725) );
  AOI22D1BWP30P140LVT U15300 ( .A1(n10803), .A2(
        inner_first_stage_data_reg[175]), .B1(n10804), .B2(
        inner_first_stage_data_reg[143]), .ZN(n10724) );
  AOI22D1BWP30P140LVT U15301 ( .A1(n10808), .A2(inner_first_stage_data_reg[15]), .B1(n10806), .B2(inner_first_stage_data_reg[111]), .ZN(n10723) );
  ND2D1BWP30P140LVT U15302 ( .A1(n10807), .A2(inner_first_stage_data_reg[47]), 
        .ZN(n10722) );
  ND4D1BWP30P140LVT U15303 ( .A1(n10725), .A2(n10724), .A3(n10723), .A4(n10722), .ZN(n10726) );
  AO21D1BWP30P140LVT U15304 ( .A1(n10814), .A2(inner_first_stage_data_reg[79]), 
        .B(n10726), .Z(N2244) );
  AOI22D1BWP30P140LVT U15305 ( .A1(n10803), .A2(
        inner_first_stage_data_reg[176]), .B1(n10802), .B2(
        inner_first_stage_data_reg[208]), .ZN(n10730) );
  AOI22D1BWP30P140LVT U15306 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[240]), .B1(n10807), .B2(
        inner_first_stage_data_reg[48]), .ZN(n10729) );
  AOI22D1BWP30P140LVT U15307 ( .A1(n10814), .A2(inner_first_stage_data_reg[80]), .B1(n10808), .B2(inner_first_stage_data_reg[16]), .ZN(n10728) );
  ND2D1BWP30P140LVT U15308 ( .A1(n10804), .A2(inner_first_stage_data_reg[144]), 
        .ZN(n10727) );
  ND4D1BWP30P140LVT U15309 ( .A1(n10730), .A2(n10729), .A3(n10728), .A4(n10727), .ZN(n10731) );
  AO21D1BWP30P140LVT U15310 ( .A1(n10806), .A2(inner_first_stage_data_reg[112]), .B(n10731), .Z(N2245) );
  AOI22D1BWP30P140LVT U15311 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[241]), .B1(n10803), .B2(
        inner_first_stage_data_reg[177]), .ZN(n10735) );
  AOI22D1BWP30P140LVT U15312 ( .A1(n10802), .A2(
        inner_first_stage_data_reg[209]), .B1(n10807), .B2(
        inner_first_stage_data_reg[49]), .ZN(n10734) );
  AOI22D1BWP30P140LVT U15313 ( .A1(n10808), .A2(inner_first_stage_data_reg[17]), .B1(n10806), .B2(inner_first_stage_data_reg[113]), .ZN(n10733) );
  ND2D1BWP30P140LVT U15314 ( .A1(n10804), .A2(inner_first_stage_data_reg[145]), 
        .ZN(n10732) );
  ND4D1BWP30P140LVT U15315 ( .A1(n10735), .A2(n10734), .A3(n10733), .A4(n10732), .ZN(n10736) );
  AO21D1BWP30P140LVT U15316 ( .A1(n10814), .A2(inner_first_stage_data_reg[81]), 
        .B(n10736), .Z(N2246) );
  AOI22D1BWP30P140LVT U15317 ( .A1(n10803), .A2(
        inner_first_stage_data_reg[178]), .B1(n10802), .B2(
        inner_first_stage_data_reg[210]), .ZN(n10740) );
  AOI22D1BWP30P140LVT U15318 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[242]), .B1(n10808), .B2(
        inner_first_stage_data_reg[18]), .ZN(n10739) );
  AOI22D1BWP30P140LVT U15319 ( .A1(n10807), .A2(inner_first_stage_data_reg[50]), .B1(n10804), .B2(inner_first_stage_data_reg[146]), .ZN(n10738) );
  ND2D1BWP30P140LVT U15320 ( .A1(n10806), .A2(inner_first_stage_data_reg[114]), 
        .ZN(n10737) );
  ND4D1BWP30P140LVT U15321 ( .A1(n10740), .A2(n10739), .A3(n10738), .A4(n10737), .ZN(n10741) );
  AO21D1BWP30P140LVT U15322 ( .A1(n10814), .A2(inner_first_stage_data_reg[82]), 
        .B(n10741), .Z(N2247) );
  AOI22D1BWP30P140LVT U15323 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[243]), .B1(n10802), .B2(
        inner_first_stage_data_reg[211]), .ZN(n10745) );
  AOI22D1BWP30P140LVT U15324 ( .A1(n10803), .A2(
        inner_first_stage_data_reg[179]), .B1(n10804), .B2(
        inner_first_stage_data_reg[147]), .ZN(n10744) );
  AOI22D1BWP30P140LVT U15325 ( .A1(n10814), .A2(inner_first_stage_data_reg[83]), .B1(n10808), .B2(inner_first_stage_data_reg[19]), .ZN(n10743) );
  ND2D1BWP30P140LVT U15326 ( .A1(n10807), .A2(inner_first_stage_data_reg[51]), 
        .ZN(n10742) );
  ND4D1BWP30P140LVT U15327 ( .A1(n10745), .A2(n10744), .A3(n10743), .A4(n10742), .ZN(n10746) );
  AO21D1BWP30P140LVT U15328 ( .A1(n10806), .A2(inner_first_stage_data_reg[115]), .B(n10746), .Z(N2248) );
  AOI22D1BWP30P140LVT U15329 ( .A1(n10803), .A2(
        inner_first_stage_data_reg[180]), .B1(n10802), .B2(
        inner_first_stage_data_reg[212]), .ZN(n10750) );
  AOI22D1BWP30P140LVT U15330 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[244]), .B1(n10807), .B2(
        inner_first_stage_data_reg[52]), .ZN(n10749) );
  AOI22D1BWP30P140LVT U15331 ( .A1(n10814), .A2(inner_first_stage_data_reg[84]), .B1(n10804), .B2(inner_first_stage_data_reg[148]), .ZN(n10748) );
  ND2D1BWP30P140LVT U15332 ( .A1(n10808), .A2(inner_first_stage_data_reg[20]), 
        .ZN(n10747) );
  ND4D1BWP30P140LVT U15333 ( .A1(n10750), .A2(n10749), .A3(n10748), .A4(n10747), .ZN(n10751) );
  AO21D1BWP30P140LVT U15334 ( .A1(n10806), .A2(inner_first_stage_data_reg[116]), .B(n10751), .Z(N2249) );
  AOI22D1BWP30P140LVT U15335 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[245]), .B1(n10802), .B2(
        inner_first_stage_data_reg[213]), .ZN(n10755) );
  AOI22D1BWP30P140LVT U15336 ( .A1(n10803), .A2(
        inner_first_stage_data_reg[181]), .B1(n10804), .B2(
        inner_first_stage_data_reg[149]), .ZN(n10754) );
  AOI22D1BWP30P140LVT U15337 ( .A1(n10814), .A2(inner_first_stage_data_reg[85]), .B1(n10807), .B2(inner_first_stage_data_reg[53]), .ZN(n10753) );
  ND2D1BWP30P140LVT U15338 ( .A1(n10808), .A2(inner_first_stage_data_reg[21]), 
        .ZN(n10752) );
  ND4D1BWP30P140LVT U15339 ( .A1(n10755), .A2(n10754), .A3(n10753), .A4(n10752), .ZN(n10756) );
  AO21D1BWP30P140LVT U15340 ( .A1(n10806), .A2(inner_first_stage_data_reg[117]), .B(n10756), .Z(N2250) );
  AOI22D1BWP30P140LVT U15341 ( .A1(n10803), .A2(
        inner_first_stage_data_reg[182]), .B1(n10802), .B2(
        inner_first_stage_data_reg[214]), .ZN(n10760) );
  AOI22D1BWP30P140LVT U15342 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[246]), .B1(n10804), .B2(
        inner_first_stage_data_reg[150]), .ZN(n10759) );
  AOI22D1BWP30P140LVT U15343 ( .A1(n10808), .A2(inner_first_stage_data_reg[22]), .B1(n10806), .B2(inner_first_stage_data_reg[118]), .ZN(n10758) );
  ND2D1BWP30P140LVT U15344 ( .A1(n10807), .A2(inner_first_stage_data_reg[54]), 
        .ZN(n10757) );
  ND4D1BWP30P140LVT U15345 ( .A1(n10760), .A2(n10759), .A3(n10758), .A4(n10757), .ZN(n10761) );
  AO21D1BWP30P140LVT U15346 ( .A1(n10814), .A2(inner_first_stage_data_reg[86]), 
        .B(n10761), .Z(N2251) );
  AOI22D1BWP30P140LVT U15347 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[247]), .B1(n10802), .B2(
        inner_first_stage_data_reg[215]), .ZN(n10765) );
  AOI22D1BWP30P140LVT U15348 ( .A1(n10803), .A2(
        inner_first_stage_data_reg[183]), .B1(n10807), .B2(
        inner_first_stage_data_reg[55]), .ZN(n10764) );
  AOI22D1BWP30P140LVT U15349 ( .A1(n10806), .A2(
        inner_first_stage_data_reg[119]), .B1(n10804), .B2(
        inner_first_stage_data_reg[151]), .ZN(n10763) );
  ND2D1BWP30P140LVT U15350 ( .A1(n10808), .A2(inner_first_stage_data_reg[23]), 
        .ZN(n10762) );
  ND4D1BWP30P140LVT U15351 ( .A1(n10765), .A2(n10764), .A3(n10763), .A4(n10762), .ZN(n10766) );
  AO21D1BWP30P140LVT U15352 ( .A1(n10814), .A2(inner_first_stage_data_reg[87]), 
        .B(n10766), .Z(N2252) );
  AOI22D1BWP30P140LVT U15353 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[248]), .B1(n10803), .B2(
        inner_first_stage_data_reg[184]), .ZN(n10770) );
  AOI22D1BWP30P140LVT U15354 ( .A1(n10802), .A2(
        inner_first_stage_data_reg[216]), .B1(n10804), .B2(
        inner_first_stage_data_reg[152]), .ZN(n10769) );
  AOI22D1BWP30P140LVT U15355 ( .A1(n10808), .A2(inner_first_stage_data_reg[24]), .B1(n10807), .B2(inner_first_stage_data_reg[56]), .ZN(n10768) );
  ND2D1BWP30P140LVT U15356 ( .A1(n10806), .A2(inner_first_stage_data_reg[120]), 
        .ZN(n10767) );
  ND4D1BWP30P140LVT U15357 ( .A1(n10770), .A2(n10769), .A3(n10768), .A4(n10767), .ZN(n10771) );
  AO21D1BWP30P140LVT U15358 ( .A1(n10814), .A2(inner_first_stage_data_reg[88]), 
        .B(n10771), .Z(N2253) );
  AOI22D1BWP30P140LVT U15359 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[249]), .B1(n10803), .B2(
        inner_first_stage_data_reg[185]), .ZN(n10775) );
  AOI22D1BWP30P140LVT U15360 ( .A1(n10802), .A2(
        inner_first_stage_data_reg[217]), .B1(n10804), .B2(
        inner_first_stage_data_reg[153]), .ZN(n10774) );
  AOI22D1BWP30P140LVT U15361 ( .A1(n10814), .A2(inner_first_stage_data_reg[89]), .B1(n10807), .B2(inner_first_stage_data_reg[57]), .ZN(n10773) );
  ND2D1BWP30P140LVT U15362 ( .A1(n10808), .A2(inner_first_stage_data_reg[25]), 
        .ZN(n10772) );
  ND4D1BWP30P140LVT U15363 ( .A1(n10775), .A2(n10774), .A3(n10773), .A4(n10772), .ZN(n10776) );
  AO21D1BWP30P140LVT U15364 ( .A1(n10806), .A2(inner_first_stage_data_reg[121]), .B(n10776), .Z(N2254) );
  AOI22D1BWP30P140LVT U15365 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[250]), .B1(n10802), .B2(
        inner_first_stage_data_reg[218]), .ZN(n10780) );
  AOI22D1BWP30P140LVT U15366 ( .A1(n10808), .A2(inner_first_stage_data_reg[26]), .B1(n10803), .B2(inner_first_stage_data_reg[186]), .ZN(n10779) );
  AOI22D1BWP30P140LVT U15367 ( .A1(n10814), .A2(inner_first_stage_data_reg[90]), .B1(n10804), .B2(inner_first_stage_data_reg[154]), .ZN(n10778) );
  ND2D1BWP30P140LVT U15368 ( .A1(n10807), .A2(inner_first_stage_data_reg[58]), 
        .ZN(n10777) );
  ND4D1BWP30P140LVT U15369 ( .A1(n10780), .A2(n10779), .A3(n10778), .A4(n10777), .ZN(n10781) );
  AO21D1BWP30P140LVT U15370 ( .A1(n10806), .A2(inner_first_stage_data_reg[122]), .B(n10781), .Z(N2255) );
  AOI22D1BWP30P140LVT U15371 ( .A1(n10803), .A2(
        inner_first_stage_data_reg[187]), .B1(n10802), .B2(
        inner_first_stage_data_reg[219]), .ZN(n10785) );
  AOI22D1BWP30P140LVT U15372 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[251]), .B1(n10808), .B2(
        inner_first_stage_data_reg[27]), .ZN(n10784) );
  AOI22D1BWP30P140LVT U15373 ( .A1(n10806), .A2(
        inner_first_stage_data_reg[123]), .B1(n10804), .B2(
        inner_first_stage_data_reg[155]), .ZN(n10783) );
  ND2D1BWP30P140LVT U15374 ( .A1(n10807), .A2(inner_first_stage_data_reg[59]), 
        .ZN(n10782) );
  ND4D1BWP30P140LVT U15375 ( .A1(n10785), .A2(n10784), .A3(n10783), .A4(n10782), .ZN(n10786) );
  AO21D1BWP30P140LVT U15376 ( .A1(n10814), .A2(inner_first_stage_data_reg[91]), 
        .B(n10786), .Z(N2256) );
  AOI22D1BWP30P140LVT U15377 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[252]), .B1(n10802), .B2(
        inner_first_stage_data_reg[220]), .ZN(n10790) );
  AOI22D1BWP30P140LVT U15378 ( .A1(n10803), .A2(
        inner_first_stage_data_reg[188]), .B1(n10804), .B2(
        inner_first_stage_data_reg[156]), .ZN(n10789) );
  AOI22D1BWP30P140LVT U15379 ( .A1(n10814), .A2(inner_first_stage_data_reg[92]), .B1(n10808), .B2(inner_first_stage_data_reg[28]), .ZN(n10788) );
  ND2D1BWP30P140LVT U15380 ( .A1(n10807), .A2(inner_first_stage_data_reg[60]), 
        .ZN(n10787) );
  ND4D1BWP30P140LVT U15381 ( .A1(n10790), .A2(n10789), .A3(n10788), .A4(n10787), .ZN(n10791) );
  AO21D1BWP30P140LVT U15382 ( .A1(n10806), .A2(inner_first_stage_data_reg[124]), .B(n10791), .Z(N2257) );
  AOI22D1BWP30P140LVT U15383 ( .A1(n10803), .A2(
        inner_first_stage_data_reg[189]), .B1(n10802), .B2(
        inner_first_stage_data_reg[221]), .ZN(n10795) );
  AOI22D1BWP30P140LVT U15384 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[253]), .B1(n10808), .B2(
        inner_first_stage_data_reg[29]), .ZN(n10794) );
  AOI22D1BWP30P140LVT U15385 ( .A1(n10807), .A2(inner_first_stage_data_reg[61]), .B1(n10806), .B2(inner_first_stage_data_reg[125]), .ZN(n10793) );
  ND2D1BWP30P140LVT U15386 ( .A1(n10804), .A2(inner_first_stage_data_reg[157]), 
        .ZN(n10792) );
  ND4D1BWP30P140LVT U15387 ( .A1(n10795), .A2(n10794), .A3(n10793), .A4(n10792), .ZN(n10796) );
  AO21D1BWP30P140LVT U15388 ( .A1(n10814), .A2(inner_first_stage_data_reg[93]), 
        .B(n10796), .Z(N2258) );
  AOI22D1BWP30P140LVT U15389 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[254]), .B1(n10803), .B2(
        inner_first_stage_data_reg[190]), .ZN(n10800) );
  AOI22D1BWP30P140LVT U15390 ( .A1(n10802), .A2(
        inner_first_stage_data_reg[222]), .B1(n10807), .B2(
        inner_first_stage_data_reg[62]), .ZN(n10799) );
  AOI22D1BWP30P140LVT U15391 ( .A1(n10808), .A2(inner_first_stage_data_reg[30]), .B1(n10804), .B2(inner_first_stage_data_reg[158]), .ZN(n10798) );
  ND2D1BWP30P140LVT U15392 ( .A1(n10806), .A2(inner_first_stage_data_reg[126]), 
        .ZN(n10797) );
  ND4D1BWP30P140LVT U15393 ( .A1(n10800), .A2(n10799), .A3(n10798), .A4(n10797), .ZN(n10801) );
  AO21D1BWP30P140LVT U15394 ( .A1(n10814), .A2(inner_first_stage_data_reg[94]), 
        .B(n10801), .Z(N2259) );
  AOI22D1BWP30P140LVT U15395 ( .A1(n10803), .A2(
        inner_first_stage_data_reg[191]), .B1(n10802), .B2(
        inner_first_stage_data_reg[223]), .ZN(n10812) );
  AOI22D1BWP30P140LVT U15396 ( .A1(n10805), .A2(
        inner_first_stage_data_reg[255]), .B1(n10804), .B2(
        inner_first_stage_data_reg[159]), .ZN(n10811) );
  AOI22D1BWP30P140LVT U15397 ( .A1(n10807), .A2(inner_first_stage_data_reg[63]), .B1(n10806), .B2(inner_first_stage_data_reg[127]), .ZN(n10810) );
  ND2D1BWP30P140LVT U15398 ( .A1(n10808), .A2(inner_first_stage_data_reg[31]), 
        .ZN(n10809) );
  ND4D1BWP30P140LVT U15399 ( .A1(n10812), .A2(n10811), .A3(n10810), .A4(n10809), .ZN(n10813) );
  AO21D1BWP30P140LVT U15400 ( .A1(n10814), .A2(inner_first_stage_data_reg[95]), 
        .B(n10813), .Z(N2260) );
  AOI22D1BWP30P140LVT U15401 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[384]), .B1(n10939), .B2(
        inner_first_stage_data_reg[288]), .ZN(n10818) );
  AOI22D1BWP30P140LVT U15402 ( .A1(n10942), .A2(
        inner_first_stage_data_reg[256]), .B1(n10941), .B2(
        inner_first_stage_data_reg[416]), .ZN(n10817) );
  AOI22D1BWP30P140LVT U15403 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[352]), .B1(n10946), .B2(
        inner_first_stage_data_reg[480]), .ZN(n10816) );
  AOI22D1BWP30P140LVT U15404 ( .A1(n10943), .A2(
        inner_first_stage_data_reg[448]), .B1(n10945), .B2(
        inner_first_stage_data_reg[320]), .ZN(n10815) );
  ND4D1BWP30P140LVT U15405 ( .A1(n10818), .A2(n10817), .A3(n10816), .A4(n10815), .ZN(N4103) );
  AOI22D1BWP30P140LVT U15406 ( .A1(n10939), .A2(
        inner_first_stage_data_reg[289]), .B1(n10941), .B2(
        inner_first_stage_data_reg[417]), .ZN(n10822) );
  AOI22D1BWP30P140LVT U15407 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[385]), .B1(n10942), .B2(
        inner_first_stage_data_reg[257]), .ZN(n10821) );
  AOI22D1BWP30P140LVT U15408 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[353]), .B1(n10943), .B2(
        inner_first_stage_data_reg[449]), .ZN(n10820) );
  AOI22D1BWP30P140LVT U15409 ( .A1(n10946), .A2(
        inner_first_stage_data_reg[481]), .B1(n10945), .B2(
        inner_first_stage_data_reg[321]), .ZN(n10819) );
  ND4D1BWP30P140LVT U15410 ( .A1(n10822), .A2(n10821), .A3(n10820), .A4(n10819), .ZN(N4104) );
  AOI22D1BWP30P140LVT U15411 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[386]), .B1(n10942), .B2(
        inner_first_stage_data_reg[258]), .ZN(n10826) );
  AOI22D1BWP30P140LVT U15412 ( .A1(n10939), .A2(
        inner_first_stage_data_reg[290]), .B1(n10941), .B2(
        inner_first_stage_data_reg[418]), .ZN(n10825) );
  AOI22D1BWP30P140LVT U15413 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[354]), .B1(n10946), .B2(
        inner_first_stage_data_reg[482]), .ZN(n10824) );
  AOI22D1BWP30P140LVT U15414 ( .A1(n10943), .A2(
        inner_first_stage_data_reg[450]), .B1(n10945), .B2(
        inner_first_stage_data_reg[322]), .ZN(n10823) );
  ND4D1BWP30P140LVT U15415 ( .A1(n10826), .A2(n10825), .A3(n10824), .A4(n10823), .ZN(N4105) );
  AOI22D1BWP30P140LVT U15416 ( .A1(n10939), .A2(
        inner_first_stage_data_reg[291]), .B1(n10942), .B2(
        inner_first_stage_data_reg[259]), .ZN(n10830) );
  AOI22D1BWP30P140LVT U15417 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[387]), .B1(n10941), .B2(
        inner_first_stage_data_reg[419]), .ZN(n10829) );
  AOI22D1BWP30P140LVT U15418 ( .A1(n10943), .A2(
        inner_first_stage_data_reg[451]), .B1(n10945), .B2(
        inner_first_stage_data_reg[323]), .ZN(n10828) );
  AOI22D1BWP30P140LVT U15419 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[355]), .B1(n10946), .B2(
        inner_first_stage_data_reg[483]), .ZN(n10827) );
  ND4D1BWP30P140LVT U15420 ( .A1(n10830), .A2(n10829), .A3(n10828), .A4(n10827), .ZN(N4106) );
  AOI22D1BWP30P140LVT U15421 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[388]), .B1(n10942), .B2(
        inner_first_stage_data_reg[260]), .ZN(n10834) );
  AOI22D1BWP30P140LVT U15422 ( .A1(n10939), .A2(
        inner_first_stage_data_reg[292]), .B1(n10941), .B2(
        inner_first_stage_data_reg[420]), .ZN(n10833) );
  AOI22D1BWP30P140LVT U15423 ( .A1(n10946), .A2(
        inner_first_stage_data_reg[484]), .B1(n10943), .B2(
        inner_first_stage_data_reg[452]), .ZN(n10832) );
  AOI22D1BWP30P140LVT U15424 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[356]), .B1(n10945), .B2(
        inner_first_stage_data_reg[324]), .ZN(n10831) );
  ND4D1BWP30P140LVT U15425 ( .A1(n10834), .A2(n10833), .A3(n10832), .A4(n10831), .ZN(N4107) );
  AOI22D1BWP30P140LVT U15426 ( .A1(n10939), .A2(
        inner_first_stage_data_reg[293]), .B1(n10942), .B2(
        inner_first_stage_data_reg[261]), .ZN(n10838) );
  AOI22D1BWP30P140LVT U15427 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[389]), .B1(n10941), .B2(
        inner_first_stage_data_reg[421]), .ZN(n10837) );
  AOI22D1BWP30P140LVT U15428 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[357]), .B1(n10945), .B2(
        inner_first_stage_data_reg[325]), .ZN(n10836) );
  AOI22D1BWP30P140LVT U15429 ( .A1(n10946), .A2(
        inner_first_stage_data_reg[485]), .B1(n10943), .B2(
        inner_first_stage_data_reg[453]), .ZN(n10835) );
  ND4D1BWP30P140LVT U15430 ( .A1(n10838), .A2(n10837), .A3(n10836), .A4(n10835), .ZN(N4108) );
  AOI22D1BWP30P140LVT U15431 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[390]), .B1(n10939), .B2(
        inner_first_stage_data_reg[294]), .ZN(n10842) );
  AOI22D1BWP30P140LVT U15432 ( .A1(n10942), .A2(
        inner_first_stage_data_reg[262]), .B1(n10941), .B2(
        inner_first_stage_data_reg[422]), .ZN(n10841) );
  AOI22D1BWP30P140LVT U15433 ( .A1(n10946), .A2(
        inner_first_stage_data_reg[486]), .B1(n10945), .B2(
        inner_first_stage_data_reg[326]), .ZN(n10840) );
  AOI22D1BWP30P140LVT U15434 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[358]), .B1(n10943), .B2(
        inner_first_stage_data_reg[454]), .ZN(n10839) );
  ND4D1BWP30P140LVT U15435 ( .A1(n10842), .A2(n10841), .A3(n10840), .A4(n10839), .ZN(N4109) );
  AOI22D1BWP30P140LVT U15436 ( .A1(n10939), .A2(
        inner_first_stage_data_reg[295]), .B1(n10941), .B2(
        inner_first_stage_data_reg[423]), .ZN(n10846) );
  AOI22D1BWP30P140LVT U15437 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[391]), .B1(n10942), .B2(
        inner_first_stage_data_reg[263]), .ZN(n10845) );
  AOI22D1BWP30P140LVT U15438 ( .A1(n10946), .A2(
        inner_first_stage_data_reg[487]), .B1(n10943), .B2(
        inner_first_stage_data_reg[455]), .ZN(n10844) );
  AOI22D1BWP30P140LVT U15439 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[359]), .B1(n10945), .B2(
        inner_first_stage_data_reg[327]), .ZN(n10843) );
  ND4D1BWP30P140LVT U15440 ( .A1(n10846), .A2(n10845), .A3(n10844), .A4(n10843), .ZN(N4110) );
  AOI22D1BWP30P140LVT U15441 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[392]), .B1(n10942), .B2(
        inner_first_stage_data_reg[264]), .ZN(n10850) );
  AOI22D1BWP30P140LVT U15442 ( .A1(n10939), .A2(
        inner_first_stage_data_reg[296]), .B1(n10941), .B2(
        inner_first_stage_data_reg[424]), .ZN(n10849) );
  AOI22D1BWP30P140LVT U15443 ( .A1(n10946), .A2(
        inner_first_stage_data_reg[488]), .B1(n10943), .B2(
        inner_first_stage_data_reg[456]), .ZN(n10848) );
  AOI22D1BWP30P140LVT U15444 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[360]), .B1(n10945), .B2(
        inner_first_stage_data_reg[328]), .ZN(n10847) );
  ND4D1BWP30P140LVT U15445 ( .A1(n10850), .A2(n10849), .A3(n10848), .A4(n10847), .ZN(N4111) );
  AOI22D1BWP30P140LVT U15446 ( .A1(n10942), .A2(
        inner_first_stage_data_reg[265]), .B1(n10941), .B2(
        inner_first_stage_data_reg[425]), .ZN(n10854) );
  AOI22D1BWP30P140LVT U15447 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[393]), .B1(n10939), .B2(
        inner_first_stage_data_reg[297]), .ZN(n10853) );
  AOI22D1BWP30P140LVT U15448 ( .A1(n10946), .A2(
        inner_first_stage_data_reg[489]), .B1(n10945), .B2(
        inner_first_stage_data_reg[329]), .ZN(n10852) );
  AOI22D1BWP30P140LVT U15449 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[361]), .B1(n10943), .B2(
        inner_first_stage_data_reg[457]), .ZN(n10851) );
  ND4D1BWP30P140LVT U15450 ( .A1(n10854), .A2(n10853), .A3(n10852), .A4(n10851), .ZN(N4112) );
  AOI22D1BWP30P140LVT U15451 ( .A1(n10939), .A2(
        inner_first_stage_data_reg[298]), .B1(n10942), .B2(
        inner_first_stage_data_reg[266]), .ZN(n10858) );
  AOI22D1BWP30P140LVT U15452 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[394]), .B1(n10941), .B2(
        inner_first_stage_data_reg[426]), .ZN(n10857) );
  AOI22D1BWP30P140LVT U15453 ( .A1(n10943), .A2(
        inner_first_stage_data_reg[458]), .B1(n10945), .B2(
        inner_first_stage_data_reg[330]), .ZN(n10856) );
  AOI22D1BWP30P140LVT U15454 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[362]), .B1(n10946), .B2(
        inner_first_stage_data_reg[490]), .ZN(n10855) );
  ND4D1BWP30P140LVT U15455 ( .A1(n10858), .A2(n10857), .A3(n10856), .A4(n10855), .ZN(N4113) );
  AOI22D1BWP30P140LVT U15456 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[395]), .B1(n10941), .B2(
        inner_first_stage_data_reg[427]), .ZN(n10862) );
  AOI22D1BWP30P140LVT U15457 ( .A1(n10939), .A2(
        inner_first_stage_data_reg[299]), .B1(n10942), .B2(
        inner_first_stage_data_reg[267]), .ZN(n10861) );
  AOI22D1BWP30P140LVT U15458 ( .A1(n10946), .A2(
        inner_first_stage_data_reg[491]), .B1(n10943), .B2(
        inner_first_stage_data_reg[459]), .ZN(n10860) );
  AOI22D1BWP30P140LVT U15459 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[363]), .B1(n10945), .B2(
        inner_first_stage_data_reg[331]), .ZN(n10859) );
  ND4D1BWP30P140LVT U15460 ( .A1(n10862), .A2(n10861), .A3(n10860), .A4(n10859), .ZN(N4114) );
  AOI22D1BWP30P140LVT U15461 ( .A1(n10942), .A2(
        inner_first_stage_data_reg[268]), .B1(n10941), .B2(
        inner_first_stage_data_reg[428]), .ZN(n10866) );
  AOI22D1BWP30P140LVT U15462 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[396]), .B1(n10939), .B2(
        inner_first_stage_data_reg[300]), .ZN(n10865) );
  AOI22D1BWP30P140LVT U15463 ( .A1(n10943), .A2(
        inner_first_stage_data_reg[460]), .B1(n10945), .B2(
        inner_first_stage_data_reg[332]), .ZN(n10864) );
  AOI22D1BWP30P140LVT U15464 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[364]), .B1(n10946), .B2(
        inner_first_stage_data_reg[492]), .ZN(n10863) );
  ND4D1BWP30P140LVT U15465 ( .A1(n10866), .A2(n10865), .A3(n10864), .A4(n10863), .ZN(N4115) );
  AOI22D1BWP30P140LVT U15466 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[397]), .B1(n10941), .B2(
        inner_first_stage_data_reg[429]), .ZN(n10870) );
  AOI22D1BWP30P140LVT U15467 ( .A1(n10939), .A2(
        inner_first_stage_data_reg[301]), .B1(n10942), .B2(
        inner_first_stage_data_reg[269]), .ZN(n10869) );
  AOI22D1BWP30P140LVT U15468 ( .A1(n10943), .A2(
        inner_first_stage_data_reg[461]), .B1(n10945), .B2(
        inner_first_stage_data_reg[333]), .ZN(n10868) );
  AOI22D1BWP30P140LVT U15469 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[365]), .B1(n10946), .B2(
        inner_first_stage_data_reg[493]), .ZN(n10867) );
  ND4D1BWP30P140LVT U15470 ( .A1(n10870), .A2(n10869), .A3(n10868), .A4(n10867), .ZN(N4116) );
  AOI22D1BWP30P140LVT U15471 ( .A1(n10942), .A2(
        inner_first_stage_data_reg[270]), .B1(n10941), .B2(
        inner_first_stage_data_reg[430]), .ZN(n10874) );
  AOI22D1BWP30P140LVT U15472 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[398]), .B1(n10939), .B2(
        inner_first_stage_data_reg[302]), .ZN(n10873) );
  AOI22D1BWP30P140LVT U15473 ( .A1(n10943), .A2(
        inner_first_stage_data_reg[462]), .B1(n10945), .B2(
        inner_first_stage_data_reg[334]), .ZN(n10872) );
  AOI22D1BWP30P140LVT U15474 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[366]), .B1(n10946), .B2(
        inner_first_stage_data_reg[494]), .ZN(n10871) );
  ND4D1BWP30P140LVT U15475 ( .A1(n10874), .A2(n10873), .A3(n10872), .A4(n10871), .ZN(N4117) );
  AOI22D1BWP30P140LVT U15476 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[399]), .B1(n10941), .B2(
        inner_first_stage_data_reg[431]), .ZN(n10878) );
  AOI22D1BWP30P140LVT U15477 ( .A1(n10939), .A2(
        inner_first_stage_data_reg[303]), .B1(n10942), .B2(
        inner_first_stage_data_reg[271]), .ZN(n10877) );
  AOI22D1BWP30P140LVT U15478 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[367]), .B1(n10945), .B2(
        inner_first_stage_data_reg[335]), .ZN(n10876) );
  AOI22D1BWP30P140LVT U15479 ( .A1(n10946), .A2(
        inner_first_stage_data_reg[495]), .B1(n10943), .B2(
        inner_first_stage_data_reg[463]), .ZN(n10875) );
  ND4D1BWP30P140LVT U15480 ( .A1(n10878), .A2(n10877), .A3(n10876), .A4(n10875), .ZN(N4118) );
  AOI22D1BWP30P140LVT U15481 ( .A1(n10939), .A2(
        inner_first_stage_data_reg[304]), .B1(n10942), .B2(
        inner_first_stage_data_reg[272]), .ZN(n10882) );
  AOI22D1BWP30P140LVT U15482 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[400]), .B1(n10941), .B2(
        inner_first_stage_data_reg[432]), .ZN(n10881) );
  AOI22D1BWP30P140LVT U15483 ( .A1(n10943), .A2(
        inner_first_stage_data_reg[464]), .B1(n10945), .B2(
        inner_first_stage_data_reg[336]), .ZN(n10880) );
  AOI22D1BWP30P140LVT U15484 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[368]), .B1(n10946), .B2(
        inner_first_stage_data_reg[496]), .ZN(n10879) );
  ND4D1BWP30P140LVT U15485 ( .A1(n10882), .A2(n10881), .A3(n10880), .A4(n10879), .ZN(N4119) );
  AOI22D1BWP30P140LVT U15486 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[401]), .B1(n10942), .B2(
        inner_first_stage_data_reg[273]), .ZN(n10886) );
  AOI22D1BWP30P140LVT U15487 ( .A1(n10939), .A2(
        inner_first_stage_data_reg[305]), .B1(n10941), .B2(
        inner_first_stage_data_reg[433]), .ZN(n10885) );
  AOI22D1BWP30P140LVT U15488 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[369]), .B1(n10943), .B2(
        inner_first_stage_data_reg[465]), .ZN(n10884) );
  AOI22D1BWP30P140LVT U15489 ( .A1(n10946), .A2(
        inner_first_stage_data_reg[497]), .B1(n10945), .B2(
        inner_first_stage_data_reg[337]), .ZN(n10883) );
  ND4D1BWP30P140LVT U15490 ( .A1(n10886), .A2(n10885), .A3(n10884), .A4(n10883), .ZN(N4120) );
  AOI22D1BWP30P140LVT U15491 ( .A1(n10942), .A2(
        inner_first_stage_data_reg[274]), .B1(n10941), .B2(
        inner_first_stage_data_reg[434]), .ZN(n10890) );
  AOI22D1BWP30P140LVT U15492 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[402]), .B1(n10939), .B2(
        inner_first_stage_data_reg[306]), .ZN(n10889) );
  AOI22D1BWP30P140LVT U15493 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[370]), .B1(n10943), .B2(
        inner_first_stage_data_reg[466]), .ZN(n10888) );
  AOI22D1BWP30P140LVT U15494 ( .A1(n10946), .A2(
        inner_first_stage_data_reg[498]), .B1(n10945), .B2(
        inner_first_stage_data_reg[338]), .ZN(n10887) );
  ND4D1BWP30P140LVT U15495 ( .A1(n10890), .A2(n10889), .A3(n10888), .A4(n10887), .ZN(N4121) );
  AOI22D1BWP30P140LVT U15496 ( .A1(n10942), .A2(
        inner_first_stage_data_reg[275]), .B1(n10941), .B2(
        inner_first_stage_data_reg[435]), .ZN(n10894) );
  AOI22D1BWP30P140LVT U15497 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[403]), .B1(n10939), .B2(
        inner_first_stage_data_reg[307]), .ZN(n10893) );
  AOI22D1BWP30P140LVT U15498 ( .A1(n10946), .A2(
        inner_first_stage_data_reg[499]), .B1(n10945), .B2(
        inner_first_stage_data_reg[339]), .ZN(n10892) );
  AOI22D1BWP30P140LVT U15499 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[371]), .B1(n10943), .B2(
        inner_first_stage_data_reg[467]), .ZN(n10891) );
  ND4D1BWP30P140LVT U15500 ( .A1(n10894), .A2(n10893), .A3(n10892), .A4(n10891), .ZN(N4122) );
  AOI22D1BWP30P140LVT U15501 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[404]), .B1(n10939), .B2(
        inner_first_stage_data_reg[308]), .ZN(n10898) );
  AOI22D1BWP30P140LVT U15502 ( .A1(n10942), .A2(
        inner_first_stage_data_reg[276]), .B1(n10941), .B2(
        inner_first_stage_data_reg[436]), .ZN(n10897) );
  AOI22D1BWP30P140LVT U15503 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[372]), .B1(n10943), .B2(
        inner_first_stage_data_reg[468]), .ZN(n10896) );
  AOI22D1BWP30P140LVT U15504 ( .A1(n10946), .A2(
        inner_first_stage_data_reg[500]), .B1(n10945), .B2(
        inner_first_stage_data_reg[340]), .ZN(n10895) );
  ND4D1BWP30P140LVT U15505 ( .A1(n10898), .A2(n10897), .A3(n10896), .A4(n10895), .ZN(N4123) );
  AOI22D1BWP30P140LVT U15506 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[405]), .B1(n10939), .B2(
        inner_first_stage_data_reg[309]), .ZN(n10902) );
  AOI22D1BWP30P140LVT U15507 ( .A1(n10942), .A2(
        inner_first_stage_data_reg[277]), .B1(n10941), .B2(
        inner_first_stage_data_reg[437]), .ZN(n10901) );
  AOI22D1BWP30P140LVT U15508 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[373]), .B1(n10945), .B2(
        inner_first_stage_data_reg[341]), .ZN(n10900) );
  AOI22D1BWP30P140LVT U15509 ( .A1(n10946), .A2(
        inner_first_stage_data_reg[501]), .B1(n10943), .B2(
        inner_first_stage_data_reg[469]), .ZN(n10899) );
  ND4D1BWP30P140LVT U15510 ( .A1(n10902), .A2(n10901), .A3(n10900), .A4(n10899), .ZN(N4124) );
  AOI22D1BWP30P140LVT U15511 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[406]), .B1(n10942), .B2(
        inner_first_stage_data_reg[278]), .ZN(n10906) );
  AOI22D1BWP30P140LVT U15512 ( .A1(n10939), .A2(
        inner_first_stage_data_reg[310]), .B1(n10941), .B2(
        inner_first_stage_data_reg[438]), .ZN(n10905) );
  AOI22D1BWP30P140LVT U15513 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[374]), .B1(n10946), .B2(
        inner_first_stage_data_reg[502]), .ZN(n10904) );
  AOI22D1BWP30P140LVT U15514 ( .A1(n10943), .A2(
        inner_first_stage_data_reg[470]), .B1(n10945), .B2(
        inner_first_stage_data_reg[342]), .ZN(n10903) );
  ND4D1BWP30P140LVT U15515 ( .A1(n10906), .A2(n10905), .A3(n10904), .A4(n10903), .ZN(N4125) );
  AOI22D1BWP30P140LVT U15516 ( .A1(n10939), .A2(
        inner_first_stage_data_reg[311]), .B1(n10941), .B2(
        inner_first_stage_data_reg[439]), .ZN(n10910) );
  AOI22D1BWP30P140LVT U15517 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[407]), .B1(n10942), .B2(
        inner_first_stage_data_reg[279]), .ZN(n10909) );
  AOI22D1BWP30P140LVT U15518 ( .A1(n10943), .A2(
        inner_first_stage_data_reg[471]), .B1(n10945), .B2(
        inner_first_stage_data_reg[343]), .ZN(n10908) );
  AOI22D1BWP30P140LVT U15519 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[375]), .B1(n10946), .B2(
        inner_first_stage_data_reg[503]), .ZN(n10907) );
  ND4D1BWP30P140LVT U15520 ( .A1(n10910), .A2(n10909), .A3(n10908), .A4(n10907), .ZN(N4126) );
  AOI22D1BWP30P140LVT U15521 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[408]), .B1(n10941), .B2(
        inner_first_stage_data_reg[440]), .ZN(n10914) );
  AOI22D1BWP30P140LVT U15522 ( .A1(n10939), .A2(
        inner_first_stage_data_reg[312]), .B1(n10942), .B2(
        inner_first_stage_data_reg[280]), .ZN(n10913) );
  AOI22D1BWP30P140LVT U15523 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[376]), .B1(n10946), .B2(
        inner_first_stage_data_reg[504]), .ZN(n10912) );
  AOI22D1BWP30P140LVT U15524 ( .A1(n10943), .A2(
        inner_first_stage_data_reg[472]), .B1(n10945), .B2(
        inner_first_stage_data_reg[344]), .ZN(n10911) );
  ND4D1BWP30P140LVT U15525 ( .A1(n10914), .A2(n10913), .A3(n10912), .A4(n10911), .ZN(N4127) );
  AOI22D1BWP30P140LVT U15526 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[409]), .B1(n10941), .B2(
        inner_first_stage_data_reg[441]), .ZN(n10918) );
  AOI22D1BWP30P140LVT U15527 ( .A1(n10939), .A2(
        inner_first_stage_data_reg[313]), .B1(n10942), .B2(
        inner_first_stage_data_reg[281]), .ZN(n10917) );
  AOI22D1BWP30P140LVT U15528 ( .A1(n10946), .A2(
        inner_first_stage_data_reg[505]), .B1(n10945), .B2(
        inner_first_stage_data_reg[345]), .ZN(n10916) );
  AOI22D1BWP30P140LVT U15529 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[377]), .B1(n10943), .B2(
        inner_first_stage_data_reg[473]), .ZN(n10915) );
  ND4D1BWP30P140LVT U15530 ( .A1(n10918), .A2(n10917), .A3(n10916), .A4(n10915), .ZN(N4128) );
  AOI22D1BWP30P140LVT U15531 ( .A1(n10939), .A2(
        inner_first_stage_data_reg[314]), .B1(n10942), .B2(
        inner_first_stage_data_reg[282]), .ZN(n10922) );
  AOI22D1BWP30P140LVT U15532 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[410]), .B1(n10941), .B2(
        inner_first_stage_data_reg[442]), .ZN(n10921) );
  AOI22D1BWP30P140LVT U15533 ( .A1(n10946), .A2(
        inner_first_stage_data_reg[506]), .B1(n10945), .B2(
        inner_first_stage_data_reg[346]), .ZN(n10920) );
  AOI22D1BWP30P140LVT U15534 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[378]), .B1(n10943), .B2(
        inner_first_stage_data_reg[474]), .ZN(n10919) );
  ND4D1BWP30P140LVT U15535 ( .A1(n10922), .A2(n10921), .A3(n10920), .A4(n10919), .ZN(N4129) );
  AOI22D1BWP30P140LVT U15536 ( .A1(n10942), .A2(
        inner_first_stage_data_reg[283]), .B1(n10941), .B2(
        inner_first_stage_data_reg[443]), .ZN(n10926) );
  AOI22D1BWP30P140LVT U15537 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[411]), .B1(n10939), .B2(
        inner_first_stage_data_reg[315]), .ZN(n10925) );
  AOI22D1BWP30P140LVT U15538 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[379]), .B1(n10946), .B2(
        inner_first_stage_data_reg[507]), .ZN(n10924) );
  AOI22D1BWP30P140LVT U15539 ( .A1(n10943), .A2(
        inner_first_stage_data_reg[475]), .B1(n10945), .B2(
        inner_first_stage_data_reg[347]), .ZN(n10923) );
  ND4D1BWP30P140LVT U15540 ( .A1(n10926), .A2(n10925), .A3(n10924), .A4(n10923), .ZN(N4130) );
  AOI22D1BWP30P140LVT U15541 ( .A1(n10939), .A2(
        inner_first_stage_data_reg[316]), .B1(n10941), .B2(
        inner_first_stage_data_reg[444]), .ZN(n10930) );
  AOI22D1BWP30P140LVT U15542 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[412]), .B1(n10942), .B2(
        inner_first_stage_data_reg[284]), .ZN(n10929) );
  AOI22D1BWP30P140LVT U15543 ( .A1(n10946), .A2(
        inner_first_stage_data_reg[508]), .B1(n10945), .B2(
        inner_first_stage_data_reg[348]), .ZN(n10928) );
  AOI22D1BWP30P140LVT U15544 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[380]), .B1(n10943), .B2(
        inner_first_stage_data_reg[476]), .ZN(n10927) );
  ND4D1BWP30P140LVT U15545 ( .A1(n10930), .A2(n10929), .A3(n10928), .A4(n10927), .ZN(N4131) );
  AOI22D1BWP30P140LVT U15546 ( .A1(n10939), .A2(
        inner_first_stage_data_reg[317]), .B1(n10942), .B2(
        inner_first_stage_data_reg[285]), .ZN(n10934) );
  AOI22D1BWP30P140LVT U15547 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[413]), .B1(n10941), .B2(
        inner_first_stage_data_reg[445]), .ZN(n10933) );
  AOI22D1BWP30P140LVT U15548 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[381]), .B1(n10943), .B2(
        inner_first_stage_data_reg[477]), .ZN(n10932) );
  AOI22D1BWP30P140LVT U15549 ( .A1(n10946), .A2(
        inner_first_stage_data_reg[509]), .B1(n10945), .B2(
        inner_first_stage_data_reg[349]), .ZN(n10931) );
  ND4D1BWP30P140LVT U15550 ( .A1(n10934), .A2(n10933), .A3(n10932), .A4(n10931), .ZN(N4132) );
  AOI22D1BWP30P140LVT U15551 ( .A1(n10942), .A2(
        inner_first_stage_data_reg[286]), .B1(n10941), .B2(
        inner_first_stage_data_reg[446]), .ZN(n10938) );
  AOI22D1BWP30P140LVT U15552 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[414]), .B1(n10939), .B2(
        inner_first_stage_data_reg[318]), .ZN(n10937) );
  AOI22D1BWP30P140LVT U15553 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[382]), .B1(n10946), .B2(
        inner_first_stage_data_reg[510]), .ZN(n10936) );
  AOI22D1BWP30P140LVT U15554 ( .A1(n10943), .A2(
        inner_first_stage_data_reg[478]), .B1(n10945), .B2(
        inner_first_stage_data_reg[350]), .ZN(n10935) );
  ND4D1BWP30P140LVT U15555 ( .A1(n10938), .A2(n10937), .A3(n10936), .A4(n10935), .ZN(N4133) );
  AOI22D1BWP30P140LVT U15556 ( .A1(n10940), .A2(
        inner_first_stage_data_reg[415]), .B1(n10939), .B2(
        inner_first_stage_data_reg[319]), .ZN(n10950) );
  AOI22D1BWP30P140LVT U15557 ( .A1(n10942), .A2(
        inner_first_stage_data_reg[287]), .B1(n10941), .B2(
        inner_first_stage_data_reg[447]), .ZN(n10949) );
  AOI22D1BWP30P140LVT U15558 ( .A1(n10944), .A2(
        inner_first_stage_data_reg[383]), .B1(n10943), .B2(
        inner_first_stage_data_reg[479]), .ZN(n10948) );
  AOI22D1BWP30P140LVT U15559 ( .A1(n10946), .A2(
        inner_first_stage_data_reg[511]), .B1(n10945), .B2(
        inner_first_stage_data_reg[351]), .ZN(n10947) );
  ND4D1BWP30P140LVT U15560 ( .A1(n10950), .A2(n10949), .A3(n10948), .A4(n10947), .ZN(N4134) );
  AOI22D1BWP30P140LVT U15561 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[512]), .B1(n11076), .B2(
        inner_first_stage_data_reg[544]), .ZN(n10954) );
  AOI22D1BWP30P140LVT U15562 ( .A1(n11075), .A2(
        inner_first_stage_data_reg[640]), .B1(n11079), .B2(
        inner_first_stage_data_reg[672]), .ZN(n10953) );
  AOI22D1BWP30P140LVT U15563 ( .A1(n11078), .A2(
        inner_first_stage_data_reg[704]), .B1(n11077), .B2(
        inner_first_stage_data_reg[736]), .ZN(n10952) );
  AOI22D1BWP30P140LVT U15564 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[576]), .B1(n11081), .B2(
        inner_first_stage_data_reg[608]), .ZN(n10951) );
  ND4D1BWP30P140LVT U15565 ( .A1(n10954), .A2(n10953), .A3(n10952), .A4(n10951), .ZN(N5977) );
  AOI22D1BWP30P140LVT U15566 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[545]), .B1(n11079), .B2(
        inner_first_stage_data_reg[673]), .ZN(n10958) );
  AOI22D1BWP30P140LVT U15567 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[513]), .B1(n11077), .B2(
        inner_first_stage_data_reg[737]), .ZN(n10957) );
  AOI22D1BWP30P140LVT U15568 ( .A1(n11075), .A2(
        inner_first_stage_data_reg[641]), .B1(n11078), .B2(
        inner_first_stage_data_reg[705]), .ZN(n10956) );
  AOI22D1BWP30P140LVT U15569 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[577]), .B1(n11081), .B2(
        inner_first_stage_data_reg[609]), .ZN(n10955) );
  ND4D1BWP30P140LVT U15570 ( .A1(n10958), .A2(n10957), .A3(n10956), .A4(n10955), .ZN(N5978) );
  AOI22D1BWP30P140LVT U15571 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[514]), .B1(n11078), .B2(
        inner_first_stage_data_reg[706]), .ZN(n10962) );
  AOI22D1BWP30P140LVT U15572 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[546]), .B1(n11079), .B2(
        inner_first_stage_data_reg[674]), .ZN(n10961) );
  AOI22D1BWP30P140LVT U15573 ( .A1(n11075), .A2(
        inner_first_stage_data_reg[642]), .B1(n11077), .B2(
        inner_first_stage_data_reg[738]), .ZN(n10960) );
  AOI22D1BWP30P140LVT U15574 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[578]), .B1(n11081), .B2(
        inner_first_stage_data_reg[610]), .ZN(n10959) );
  ND4D1BWP30P140LVT U15575 ( .A1(n10962), .A2(n10961), .A3(n10960), .A4(n10959), .ZN(N5979) );
  AOI22D1BWP30P140LVT U15576 ( .A1(n11075), .A2(
        inner_first_stage_data_reg[643]), .B1(n11077), .B2(
        inner_first_stage_data_reg[739]), .ZN(n10966) );
  AOI22D1BWP30P140LVT U15577 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[515]), .B1(n11076), .B2(
        inner_first_stage_data_reg[547]), .ZN(n10965) );
  AOI22D1BWP30P140LVT U15578 ( .A1(n11079), .A2(
        inner_first_stage_data_reg[675]), .B1(n11078), .B2(
        inner_first_stage_data_reg[707]), .ZN(n10964) );
  AOI22D1BWP30P140LVT U15579 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[579]), .B1(n11081), .B2(
        inner_first_stage_data_reg[611]), .ZN(n10963) );
  ND4D1BWP30P140LVT U15580 ( .A1(n10966), .A2(n10965), .A3(n10964), .A4(n10963), .ZN(N5980) );
  AOI22D1BWP30P140LVT U15581 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[548]), .B1(n11077), .B2(
        inner_first_stage_data_reg[740]), .ZN(n10970) );
  AOI22D1BWP30P140LVT U15582 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[516]), .B1(n11078), .B2(
        inner_first_stage_data_reg[708]), .ZN(n10969) );
  AOI22D1BWP30P140LVT U15583 ( .A1(n11075), .A2(
        inner_first_stage_data_reg[644]), .B1(n11079), .B2(
        inner_first_stage_data_reg[676]), .ZN(n10968) );
  AOI22D1BWP30P140LVT U15584 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[580]), .B1(n11081), .B2(
        inner_first_stage_data_reg[612]), .ZN(n10967) );
  ND4D1BWP30P140LVT U15585 ( .A1(n10970), .A2(n10969), .A3(n10968), .A4(n10967), .ZN(N5981) );
  AOI22D1BWP30P140LVT U15586 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[549]), .B1(n11077), .B2(
        inner_first_stage_data_reg[741]), .ZN(n10974) );
  AOI22D1BWP30P140LVT U15587 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[517]), .B1(n11078), .B2(
        inner_first_stage_data_reg[709]), .ZN(n10973) );
  AOI22D1BWP30P140LVT U15588 ( .A1(n11075), .A2(
        inner_first_stage_data_reg[645]), .B1(n11079), .B2(
        inner_first_stage_data_reg[677]), .ZN(n10972) );
  AOI22D1BWP30P140LVT U15589 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[581]), .B1(n11081), .B2(
        inner_first_stage_data_reg[613]), .ZN(n10971) );
  ND4D1BWP30P140LVT U15590 ( .A1(n10974), .A2(n10973), .A3(n10972), .A4(n10971), .ZN(N5982) );
  AOI22D1BWP30P140LVT U15591 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[518]), .B1(n11077), .B2(
        inner_first_stage_data_reg[742]), .ZN(n10978) );
  AOI22D1BWP30P140LVT U15592 ( .A1(n11079), .A2(
        inner_first_stage_data_reg[678]), .B1(n11078), .B2(
        inner_first_stage_data_reg[710]), .ZN(n10977) );
  AOI22D1BWP30P140LVT U15593 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[550]), .B1(n11075), .B2(
        inner_first_stage_data_reg[646]), .ZN(n10976) );
  AOI22D1BWP30P140LVT U15594 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[582]), .B1(n11081), .B2(
        inner_first_stage_data_reg[614]), .ZN(n10975) );
  ND4D1BWP30P140LVT U15595 ( .A1(n10978), .A2(n10977), .A3(n10976), .A4(n10975), .ZN(N5983) );
  AOI22D1BWP30P140LVT U15596 ( .A1(n11079), .A2(
        inner_first_stage_data_reg[679]), .B1(n11078), .B2(
        inner_first_stage_data_reg[711]), .ZN(n10982) );
  AOI22D1BWP30P140LVT U15597 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[519]), .B1(n11075), .B2(
        inner_first_stage_data_reg[647]), .ZN(n10981) );
  AOI22D1BWP30P140LVT U15598 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[551]), .B1(n11077), .B2(
        inner_first_stage_data_reg[743]), .ZN(n10980) );
  AOI22D1BWP30P140LVT U15599 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[583]), .B1(n11081), .B2(
        inner_first_stage_data_reg[615]), .ZN(n10979) );
  ND4D1BWP30P140LVT U15600 ( .A1(n10982), .A2(n10981), .A3(n10980), .A4(n10979), .ZN(N5984) );
  AOI22D1BWP30P140LVT U15601 ( .A1(n11079), .A2(
        inner_first_stage_data_reg[680]), .B1(n11078), .B2(
        inner_first_stage_data_reg[712]), .ZN(n10986) );
  AOI22D1BWP30P140LVT U15602 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[520]), .B1(n11077), .B2(
        inner_first_stage_data_reg[744]), .ZN(n10985) );
  AOI22D1BWP30P140LVT U15603 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[552]), .B1(n11075), .B2(
        inner_first_stage_data_reg[648]), .ZN(n10984) );
  AOI22D1BWP30P140LVT U15604 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[584]), .B1(n11081), .B2(
        inner_first_stage_data_reg[616]), .ZN(n10983) );
  ND4D1BWP30P140LVT U15605 ( .A1(n10986), .A2(n10985), .A3(n10984), .A4(n10983), .ZN(N5985) );
  AOI22D1BWP30P140LVT U15606 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[553]), .B1(n11077), .B2(
        inner_first_stage_data_reg[745]), .ZN(n10990) );
  AOI22D1BWP30P140LVT U15607 ( .A1(n11079), .A2(
        inner_first_stage_data_reg[681]), .B1(n11078), .B2(
        inner_first_stage_data_reg[713]), .ZN(n10989) );
  AOI22D1BWP30P140LVT U15608 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[521]), .B1(n11075), .B2(
        inner_first_stage_data_reg[649]), .ZN(n10988) );
  AOI22D1BWP30P140LVT U15609 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[585]), .B1(n11081), .B2(
        inner_first_stage_data_reg[617]), .ZN(n10987) );
  ND4D1BWP30P140LVT U15610 ( .A1(n10990), .A2(n10989), .A3(n10988), .A4(n10987), .ZN(N5986) );
  AOI22D1BWP30P140LVT U15611 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[554]), .B1(n11077), .B2(
        inner_first_stage_data_reg[746]), .ZN(n10994) );
  AOI22D1BWP30P140LVT U15612 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[522]), .B1(n11078), .B2(
        inner_first_stage_data_reg[714]), .ZN(n10993) );
  AOI22D1BWP30P140LVT U15613 ( .A1(n11075), .A2(
        inner_first_stage_data_reg[650]), .B1(n11079), .B2(
        inner_first_stage_data_reg[682]), .ZN(n10992) );
  AOI22D1BWP30P140LVT U15614 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[586]), .B1(n11081), .B2(
        inner_first_stage_data_reg[618]), .ZN(n10991) );
  ND4D1BWP30P140LVT U15615 ( .A1(n10994), .A2(n10993), .A3(n10992), .A4(n10991), .ZN(N5987) );
  AOI22D1BWP30P140LVT U15616 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[523]), .B1(n11078), .B2(
        inner_first_stage_data_reg[715]), .ZN(n10998) );
  AOI22D1BWP30P140LVT U15617 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[555]), .B1(n11079), .B2(
        inner_first_stage_data_reg[683]), .ZN(n10997) );
  AOI22D1BWP30P140LVT U15618 ( .A1(n11075), .A2(
        inner_first_stage_data_reg[651]), .B1(n11077), .B2(
        inner_first_stage_data_reg[747]), .ZN(n10996) );
  AOI22D1BWP30P140LVT U15619 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[587]), .B1(n11081), .B2(
        inner_first_stage_data_reg[619]), .ZN(n10995) );
  ND4D1BWP30P140LVT U15620 ( .A1(n10998), .A2(n10997), .A3(n10996), .A4(n10995), .ZN(N5988) );
  AOI22D1BWP30P140LVT U15621 ( .A1(n11075), .A2(
        inner_first_stage_data_reg[652]), .B1(n11078), .B2(
        inner_first_stage_data_reg[716]), .ZN(n11002) );
  AOI22D1BWP30P140LVT U15622 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[524]), .B1(n11076), .B2(
        inner_first_stage_data_reg[556]), .ZN(n11001) );
  AOI22D1BWP30P140LVT U15623 ( .A1(n11079), .A2(
        inner_first_stage_data_reg[684]), .B1(n11077), .B2(
        inner_first_stage_data_reg[748]), .ZN(n11000) );
  AOI22D1BWP30P140LVT U15624 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[588]), .B1(n11081), .B2(
        inner_first_stage_data_reg[620]), .ZN(n10999) );
  ND4D1BWP30P140LVT U15625 ( .A1(n11002), .A2(n11001), .A3(n11000), .A4(n10999), .ZN(N5989) );
  AOI22D1BWP30P140LVT U15626 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[557]), .B1(n11077), .B2(
        inner_first_stage_data_reg[749]), .ZN(n11006) );
  AOI22D1BWP30P140LVT U15627 ( .A1(n11075), .A2(
        inner_first_stage_data_reg[653]), .B1(n11079), .B2(
        inner_first_stage_data_reg[685]), .ZN(n11005) );
  AOI22D1BWP30P140LVT U15628 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[525]), .B1(n11078), .B2(
        inner_first_stage_data_reg[717]), .ZN(n11004) );
  AOI22D1BWP30P140LVT U15629 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[589]), .B1(n11081), .B2(
        inner_first_stage_data_reg[621]), .ZN(n11003) );
  ND4D1BWP30P140LVT U15630 ( .A1(n11006), .A2(n11005), .A3(n11004), .A4(n11003), .ZN(N5990) );
  AOI22D1BWP30P140LVT U15631 ( .A1(n11078), .A2(
        inner_first_stage_data_reg[718]), .B1(n11077), .B2(
        inner_first_stage_data_reg[750]), .ZN(n11010) );
  AOI22D1BWP30P140LVT U15632 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[558]), .B1(n11079), .B2(
        inner_first_stage_data_reg[686]), .ZN(n11009) );
  AOI22D1BWP30P140LVT U15633 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[526]), .B1(n11075), .B2(
        inner_first_stage_data_reg[654]), .ZN(n11008) );
  AOI22D1BWP30P140LVT U15634 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[590]), .B1(n11081), .B2(
        inner_first_stage_data_reg[622]), .ZN(n11007) );
  ND4D1BWP30P140LVT U15635 ( .A1(n11010), .A2(n11009), .A3(n11008), .A4(n11007), .ZN(N5991) );
  AOI22D1BWP30P140LVT U15636 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[559]), .B1(n11079), .B2(
        inner_first_stage_data_reg[687]), .ZN(n11014) );
  AOI22D1BWP30P140LVT U15637 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[527]), .B1(n11075), .B2(
        inner_first_stage_data_reg[655]), .ZN(n11013) );
  AOI22D1BWP30P140LVT U15638 ( .A1(n11078), .A2(
        inner_first_stage_data_reg[719]), .B1(n11077), .B2(
        inner_first_stage_data_reg[751]), .ZN(n11012) );
  AOI22D1BWP30P140LVT U15639 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[591]), .B1(n11081), .B2(
        inner_first_stage_data_reg[623]), .ZN(n11011) );
  ND4D1BWP30P140LVT U15640 ( .A1(n11014), .A2(n11013), .A3(n11012), .A4(n11011), .ZN(N5992) );
  AOI22D1BWP30P140LVT U15641 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[528]), .B1(n11079), .B2(
        inner_first_stage_data_reg[688]), .ZN(n11018) );
  AOI22D1BWP30P140LVT U15642 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[560]), .B1(n11078), .B2(
        inner_first_stage_data_reg[720]), .ZN(n11017) );
  AOI22D1BWP30P140LVT U15643 ( .A1(n11075), .A2(
        inner_first_stage_data_reg[656]), .B1(n11077), .B2(
        inner_first_stage_data_reg[752]), .ZN(n11016) );
  AOI22D1BWP30P140LVT U15644 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[592]), .B1(n11081), .B2(
        inner_first_stage_data_reg[624]), .ZN(n11015) );
  ND4D1BWP30P140LVT U15645 ( .A1(n11018), .A2(n11017), .A3(n11016), .A4(n11015), .ZN(N5993) );
  AOI22D1BWP30P140LVT U15646 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[561]), .B1(n11075), .B2(
        inner_first_stage_data_reg[657]), .ZN(n11022) );
  AOI22D1BWP30P140LVT U15647 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[529]), .B1(n11078), .B2(
        inner_first_stage_data_reg[721]), .ZN(n11021) );
  AOI22D1BWP30P140LVT U15648 ( .A1(n11079), .A2(
        inner_first_stage_data_reg[689]), .B1(n11077), .B2(
        inner_first_stage_data_reg[753]), .ZN(n11020) );
  AOI22D1BWP30P140LVT U15649 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[593]), .B1(n11081), .B2(
        inner_first_stage_data_reg[625]), .ZN(n11019) );
  ND4D1BWP30P140LVT U15650 ( .A1(n11022), .A2(n11021), .A3(n11020), .A4(n11019), .ZN(N5994) );
  AOI22D1BWP30P140LVT U15651 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[530]), .B1(n11077), .B2(
        inner_first_stage_data_reg[754]), .ZN(n11026) );
  AOI22D1BWP30P140LVT U15652 ( .A1(n11079), .A2(
        inner_first_stage_data_reg[690]), .B1(n11078), .B2(
        inner_first_stage_data_reg[722]), .ZN(n11025) );
  AOI22D1BWP30P140LVT U15653 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[562]), .B1(n11075), .B2(
        inner_first_stage_data_reg[658]), .ZN(n11024) );
  AOI22D1BWP30P140LVT U15654 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[594]), .B1(n11081), .B2(
        inner_first_stage_data_reg[626]), .ZN(n11023) );
  ND4D1BWP30P140LVT U15655 ( .A1(n11026), .A2(n11025), .A3(n11024), .A4(n11023), .ZN(N5995) );
  AOI22D1BWP30P140LVT U15656 ( .A1(n11079), .A2(
        inner_first_stage_data_reg[691]), .B1(n11078), .B2(
        inner_first_stage_data_reg[723]), .ZN(n11030) );
  AOI22D1BWP30P140LVT U15657 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[563]), .B1(n11075), .B2(
        inner_first_stage_data_reg[659]), .ZN(n11029) );
  AOI22D1BWP30P140LVT U15658 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[531]), .B1(n11077), .B2(
        inner_first_stage_data_reg[755]), .ZN(n11028) );
  AOI22D1BWP30P140LVT U15659 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[595]), .B1(n11081), .B2(
        inner_first_stage_data_reg[627]), .ZN(n11027) );
  ND4D1BWP30P140LVT U15660 ( .A1(n11030), .A2(n11029), .A3(n11028), .A4(n11027), .ZN(N5996) );
  AOI22D1BWP30P140LVT U15661 ( .A1(n11075), .A2(
        inner_first_stage_data_reg[660]), .B1(n11078), .B2(
        inner_first_stage_data_reg[724]), .ZN(n11034) );
  AOI22D1BWP30P140LVT U15662 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[532]), .B1(n11077), .B2(
        inner_first_stage_data_reg[756]), .ZN(n11033) );
  AOI22D1BWP30P140LVT U15663 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[564]), .B1(n11079), .B2(
        inner_first_stage_data_reg[692]), .ZN(n11032) );
  AOI22D1BWP30P140LVT U15664 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[596]), .B1(n11081), .B2(
        inner_first_stage_data_reg[628]), .ZN(n11031) );
  ND4D1BWP30P140LVT U15665 ( .A1(n11034), .A2(n11033), .A3(n11032), .A4(n11031), .ZN(N5997) );
  AOI22D1BWP30P140LVT U15666 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[533]), .B1(n11076), .B2(
        inner_first_stage_data_reg[565]), .ZN(n11038) );
  AOI22D1BWP30P140LVT U15667 ( .A1(n11079), .A2(
        inner_first_stage_data_reg[693]), .B1(n11078), .B2(
        inner_first_stage_data_reg[725]), .ZN(n11037) );
  AOI22D1BWP30P140LVT U15668 ( .A1(n11075), .A2(
        inner_first_stage_data_reg[661]), .B1(n11077), .B2(
        inner_first_stage_data_reg[757]), .ZN(n11036) );
  AOI22D1BWP30P140LVT U15669 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[597]), .B1(n11081), .B2(
        inner_first_stage_data_reg[629]), .ZN(n11035) );
  ND4D1BWP30P140LVT U15670 ( .A1(n11038), .A2(n11037), .A3(n11036), .A4(n11035), .ZN(N5998) );
  AOI22D1BWP30P140LVT U15671 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[566]), .B1(n11079), .B2(
        inner_first_stage_data_reg[694]), .ZN(n11042) );
  AOI22D1BWP30P140LVT U15672 ( .A1(n11075), .A2(
        inner_first_stage_data_reg[662]), .B1(n11078), .B2(
        inner_first_stage_data_reg[726]), .ZN(n11041) );
  AOI22D1BWP30P140LVT U15673 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[534]), .B1(n11077), .B2(
        inner_first_stage_data_reg[758]), .ZN(n11040) );
  AOI22D1BWP30P140LVT U15674 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[598]), .B1(n11081), .B2(
        inner_first_stage_data_reg[630]), .ZN(n11039) );
  ND4D1BWP30P140LVT U15675 ( .A1(n11042), .A2(n11041), .A3(n11040), .A4(n11039), .ZN(N5999) );
  AOI22D1BWP30P140LVT U15676 ( .A1(n11078), .A2(
        inner_first_stage_data_reg[727]), .B1(n11077), .B2(
        inner_first_stage_data_reg[759]), .ZN(n11046) );
  AOI22D1BWP30P140LVT U15677 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[535]), .B1(n11075), .B2(
        inner_first_stage_data_reg[663]), .ZN(n11045) );
  AOI22D1BWP30P140LVT U15678 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[567]), .B1(n11079), .B2(
        inner_first_stage_data_reg[695]), .ZN(n11044) );
  AOI22D1BWP30P140LVT U15679 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[599]), .B1(n11081), .B2(
        inner_first_stage_data_reg[631]), .ZN(n11043) );
  ND4D1BWP30P140LVT U15680 ( .A1(n11046), .A2(n11045), .A3(n11044), .A4(n11043), .ZN(N6000) );
  AOI22D1BWP30P140LVT U15681 ( .A1(n11075), .A2(
        inner_first_stage_data_reg[664]), .B1(n11077), .B2(
        inner_first_stage_data_reg[760]), .ZN(n11050) );
  AOI22D1BWP30P140LVT U15682 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[536]), .B1(n11076), .B2(
        inner_first_stage_data_reg[568]), .ZN(n11049) );
  AOI22D1BWP30P140LVT U15683 ( .A1(n11079), .A2(
        inner_first_stage_data_reg[696]), .B1(n11078), .B2(
        inner_first_stage_data_reg[728]), .ZN(n11048) );
  AOI22D1BWP30P140LVT U15684 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[600]), .B1(n11081), .B2(
        inner_first_stage_data_reg[632]), .ZN(n11047) );
  ND4D1BWP30P140LVT U15685 ( .A1(n11050), .A2(n11049), .A3(n11048), .A4(n11047), .ZN(N6001) );
  AOI22D1BWP30P140LVT U15686 ( .A1(n11075), .A2(
        inner_first_stage_data_reg[665]), .B1(n11077), .B2(
        inner_first_stage_data_reg[761]), .ZN(n11054) );
  AOI22D1BWP30P140LVT U15687 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[537]), .B1(n11078), .B2(
        inner_first_stage_data_reg[729]), .ZN(n11053) );
  AOI22D1BWP30P140LVT U15688 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[569]), .B1(n11079), .B2(
        inner_first_stage_data_reg[697]), .ZN(n11052) );
  AOI22D1BWP30P140LVT U15689 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[601]), .B1(n11081), .B2(
        inner_first_stage_data_reg[633]), .ZN(n11051) );
  ND4D1BWP30P140LVT U15690 ( .A1(n11054), .A2(n11053), .A3(n11052), .A4(n11051), .ZN(N6002) );
  AOI22D1BWP30P140LVT U15691 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[538]), .B1(n11075), .B2(
        inner_first_stage_data_reg[666]), .ZN(n11058) );
  AOI22D1BWP30P140LVT U15692 ( .A1(n11078), .A2(
        inner_first_stage_data_reg[730]), .B1(n11077), .B2(
        inner_first_stage_data_reg[762]), .ZN(n11057) );
  AOI22D1BWP30P140LVT U15693 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[570]), .B1(n11079), .B2(
        inner_first_stage_data_reg[698]), .ZN(n11056) );
  AOI22D1BWP30P140LVT U15694 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[602]), .B1(n11081), .B2(
        inner_first_stage_data_reg[634]), .ZN(n11055) );
  ND4D1BWP30P140LVT U15695 ( .A1(n11058), .A2(n11057), .A3(n11056), .A4(n11055), .ZN(N6003) );
  AOI22D1BWP30P140LVT U15696 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[571]), .B1(n11077), .B2(
        inner_first_stage_data_reg[763]), .ZN(n11062) );
  AOI22D1BWP30P140LVT U15697 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[539]), .B1(n11075), .B2(
        inner_first_stage_data_reg[667]), .ZN(n11061) );
  AOI22D1BWP30P140LVT U15698 ( .A1(n11079), .A2(
        inner_first_stage_data_reg[699]), .B1(n11078), .B2(
        inner_first_stage_data_reg[731]), .ZN(n11060) );
  AOI22D1BWP30P140LVT U15699 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[603]), .B1(n11081), .B2(
        inner_first_stage_data_reg[635]), .ZN(n11059) );
  ND4D1BWP30P140LVT U15700 ( .A1(n11062), .A2(n11061), .A3(n11060), .A4(n11059), .ZN(N6004) );
  AOI22D1BWP30P140LVT U15701 ( .A1(n11079), .A2(
        inner_first_stage_data_reg[700]), .B1(n11078), .B2(
        inner_first_stage_data_reg[732]), .ZN(n11066) );
  AOI22D1BWP30P140LVT U15702 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[540]), .B1(n11077), .B2(
        inner_first_stage_data_reg[764]), .ZN(n11065) );
  AOI22D1BWP30P140LVT U15703 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[572]), .B1(n11075), .B2(
        inner_first_stage_data_reg[668]), .ZN(n11064) );
  AOI22D1BWP30P140LVT U15704 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[604]), .B1(n11081), .B2(
        inner_first_stage_data_reg[636]), .ZN(n11063) );
  ND4D1BWP30P140LVT U15705 ( .A1(n11066), .A2(n11065), .A3(n11064), .A4(n11063), .ZN(N6005) );
  AOI22D1BWP30P140LVT U15706 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[541]), .B1(n11075), .B2(
        inner_first_stage_data_reg[669]), .ZN(n11070) );
  AOI22D1BWP30P140LVT U15707 ( .A1(n11079), .A2(
        inner_first_stage_data_reg[701]), .B1(n11077), .B2(
        inner_first_stage_data_reg[765]), .ZN(n11069) );
  AOI22D1BWP30P140LVT U15708 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[573]), .B1(n11078), .B2(
        inner_first_stage_data_reg[733]), .ZN(n11068) );
  AOI22D1BWP30P140LVT U15709 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[605]), .B1(n11081), .B2(
        inner_first_stage_data_reg[637]), .ZN(n11067) );
  ND4D1BWP30P140LVT U15710 ( .A1(n11070), .A2(n11069), .A3(n11068), .A4(n11067), .ZN(N6006) );
  AOI22D1BWP30P140LVT U15711 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[574]), .B1(n11078), .B2(
        inner_first_stage_data_reg[734]), .ZN(n11074) );
  AOI22D1BWP30P140LVT U15712 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[542]), .B1(n11079), .B2(
        inner_first_stage_data_reg[702]), .ZN(n11073) );
  AOI22D1BWP30P140LVT U15713 ( .A1(n11075), .A2(
        inner_first_stage_data_reg[670]), .B1(n11077), .B2(
        inner_first_stage_data_reg[766]), .ZN(n11072) );
  AOI22D1BWP30P140LVT U15714 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[606]), .B1(n11081), .B2(
        inner_first_stage_data_reg[638]), .ZN(n11071) );
  ND4D1BWP30P140LVT U15715 ( .A1(n11074), .A2(n11073), .A3(n11072), .A4(n11071), .ZN(N6007) );
  AOI22D1BWP30P140LVT U15716 ( .A1(n11076), .A2(
        inner_first_stage_data_reg[575]), .B1(n11075), .B2(
        inner_first_stage_data_reg[671]), .ZN(n11086) );
  AOI22D1BWP30P140LVT U15717 ( .A1(n11078), .A2(
        inner_first_stage_data_reg[735]), .B1(n11077), .B2(
        inner_first_stage_data_reg[767]), .ZN(n11085) );
  AOI22D1BWP30P140LVT U15718 ( .A1(n11080), .A2(
        inner_first_stage_data_reg[543]), .B1(n11079), .B2(
        inner_first_stage_data_reg[703]), .ZN(n11084) );
  AOI22D1BWP30P140LVT U15719 ( .A1(n11082), .A2(
        inner_first_stage_data_reg[607]), .B1(n11081), .B2(
        inner_first_stage_data_reg[639]), .ZN(n11083) );
  ND4D1BWP30P140LVT U15720 ( .A1(n11086), .A2(n11085), .A3(n11084), .A4(n11083), .ZN(N6008) );
  AOI22D1BWP30P140LVT U15721 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[768]), .B1(n11216), .B2(
        inner_first_stage_data_reg[864]), .ZN(n11090) );
  AOI22D1BWP30P140LVT U15722 ( .A1(n11215), .A2(
        inner_first_stage_data_reg[928]), .B1(n11213), .B2(
        inner_first_stage_data_reg[800]), .ZN(n11089) );
  AOI22D1BWP30P140LVT U15723 ( .A1(n11212), .A2(
        inner_first_stage_data_reg[896]), .B1(n11211), .B2(
        inner_first_stage_data_reg[832]), .ZN(n11088) );
  AOI22D1BWP30P140LVT U15724 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[992]), .B1(n11217), .B2(
        inner_first_stage_data_reg[960]), .ZN(n11087) );
  ND4D1BWP30P140LVT U15725 ( .A1(n11090), .A2(n11089), .A3(n11088), .A4(n11087), .ZN(N7851) );
  AOI22D1BWP30P140LVT U15726 ( .A1(n11216), .A2(
        inner_first_stage_data_reg[865]), .B1(n11211), .B2(
        inner_first_stage_data_reg[833]), .ZN(n11094) );
  AOI22D1BWP30P140LVT U15727 ( .A1(n11213), .A2(
        inner_first_stage_data_reg[801]), .B1(n11212), .B2(
        inner_first_stage_data_reg[897]), .ZN(n11093) );
  AOI22D1BWP30P140LVT U15728 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[769]), .B1(n11215), .B2(
        inner_first_stage_data_reg[929]), .ZN(n11092) );
  AOI22D1BWP30P140LVT U15729 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[993]), .B1(n11217), .B2(
        inner_first_stage_data_reg[961]), .ZN(n11091) );
  ND4D1BWP30P140LVT U15730 ( .A1(n11094), .A2(n11093), .A3(n11092), .A4(n11091), .ZN(N7852) );
  AOI22D1BWP30P140LVT U15731 ( .A1(n11215), .A2(
        inner_first_stage_data_reg[930]), .B1(n11211), .B2(
        inner_first_stage_data_reg[834]), .ZN(n11098) );
  AOI22D1BWP30P140LVT U15732 ( .A1(n11213), .A2(
        inner_first_stage_data_reg[802]), .B1(n11212), .B2(
        inner_first_stage_data_reg[898]), .ZN(n11097) );
  AOI22D1BWP30P140LVT U15733 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[770]), .B1(n11216), .B2(
        inner_first_stage_data_reg[866]), .ZN(n11096) );
  AOI22D1BWP30P140LVT U15734 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[994]), .B1(n11217), .B2(
        inner_first_stage_data_reg[962]), .ZN(n11095) );
  ND4D1BWP30P140LVT U15735 ( .A1(n11098), .A2(n11097), .A3(n11096), .A4(n11095), .ZN(N7853) );
  AOI22D1BWP30P140LVT U15736 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[771]), .B1(n11216), .B2(
        inner_first_stage_data_reg[867]), .ZN(n11102) );
  AOI22D1BWP30P140LVT U15737 ( .A1(n11213), .A2(
        inner_first_stage_data_reg[803]), .B1(n11212), .B2(
        inner_first_stage_data_reg[899]), .ZN(n11101) );
  AOI22D1BWP30P140LVT U15738 ( .A1(n11215), .A2(
        inner_first_stage_data_reg[931]), .B1(n11211), .B2(
        inner_first_stage_data_reg[835]), .ZN(n11100) );
  AOI22D1BWP30P140LVT U15739 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[995]), .B1(n11217), .B2(
        inner_first_stage_data_reg[963]), .ZN(n11099) );
  ND4D1BWP30P140LVT U15740 ( .A1(n11102), .A2(n11101), .A3(n11100), .A4(n11099), .ZN(N7854) );
  AOI22D1BWP30P140LVT U15741 ( .A1(n11216), .A2(
        inner_first_stage_data_reg[868]), .B1(n11212), .B2(
        inner_first_stage_data_reg[900]), .ZN(n11106) );
  AOI22D1BWP30P140LVT U15742 ( .A1(n11213), .A2(
        inner_first_stage_data_reg[804]), .B1(n11211), .B2(
        inner_first_stage_data_reg[836]), .ZN(n11105) );
  AOI22D1BWP30P140LVT U15743 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[772]), .B1(n11215), .B2(
        inner_first_stage_data_reg[932]), .ZN(n11104) );
  AOI22D1BWP30P140LVT U15744 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[996]), .B1(n11217), .B2(
        inner_first_stage_data_reg[964]), .ZN(n11103) );
  ND4D1BWP30P140LVT U15745 ( .A1(n11106), .A2(n11105), .A3(n11104), .A4(n11103), .ZN(N7855) );
  AOI22D1BWP30P140LVT U15746 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[773]), .B1(n11216), .B2(
        inner_first_stage_data_reg[869]), .ZN(n11110) );
  AOI22D1BWP30P140LVT U15747 ( .A1(n11213), .A2(
        inner_first_stage_data_reg[805]), .B1(n11212), .B2(
        inner_first_stage_data_reg[901]), .ZN(n11109) );
  AOI22D1BWP30P140LVT U15748 ( .A1(n11215), .A2(
        inner_first_stage_data_reg[933]), .B1(n11211), .B2(
        inner_first_stage_data_reg[837]), .ZN(n11108) );
  AOI22D1BWP30P140LVT U15749 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[997]), .B1(n11217), .B2(
        inner_first_stage_data_reg[965]), .ZN(n11107) );
  ND4D1BWP30P140LVT U15750 ( .A1(n11110), .A2(n11109), .A3(n11108), .A4(n11107), .ZN(N7856) );
  AOI22D1BWP30P140LVT U15751 ( .A1(n11215), .A2(
        inner_first_stage_data_reg[934]), .B1(n11212), .B2(
        inner_first_stage_data_reg[902]), .ZN(n11114) );
  AOI22D1BWP30P140LVT U15752 ( .A1(n11216), .A2(
        inner_first_stage_data_reg[870]), .B1(n11213), .B2(
        inner_first_stage_data_reg[806]), .ZN(n11113) );
  AOI22D1BWP30P140LVT U15753 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[774]), .B1(n11211), .B2(
        inner_first_stage_data_reg[838]), .ZN(n11112) );
  AOI22D1BWP30P140LVT U15754 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[998]), .B1(n11217), .B2(
        inner_first_stage_data_reg[966]), .ZN(n11111) );
  ND4D1BWP30P140LVT U15755 ( .A1(n11114), .A2(n11113), .A3(n11112), .A4(n11111), .ZN(N7857) );
  AOI22D1BWP30P140LVT U15756 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[775]), .B1(n11212), .B2(
        inner_first_stage_data_reg[903]), .ZN(n11118) );
  AOI22D1BWP30P140LVT U15757 ( .A1(n11213), .A2(
        inner_first_stage_data_reg[807]), .B1(n11211), .B2(
        inner_first_stage_data_reg[839]), .ZN(n11117) );
  AOI22D1BWP30P140LVT U15758 ( .A1(n11216), .A2(
        inner_first_stage_data_reg[871]), .B1(n11215), .B2(
        inner_first_stage_data_reg[935]), .ZN(n11116) );
  AOI22D1BWP30P140LVT U15759 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[999]), .B1(n11217), .B2(
        inner_first_stage_data_reg[967]), .ZN(n11115) );
  ND4D1BWP30P140LVT U15760 ( .A1(n11118), .A2(n11117), .A3(n11116), .A4(n11115), .ZN(N7858) );
  AOI22D1BWP30P140LVT U15761 ( .A1(n11216), .A2(
        inner_first_stage_data_reg[872]), .B1(n11211), .B2(
        inner_first_stage_data_reg[840]), .ZN(n11122) );
  AOI22D1BWP30P140LVT U15762 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[776]), .B1(n11215), .B2(
        inner_first_stage_data_reg[936]), .ZN(n11121) );
  AOI22D1BWP30P140LVT U15763 ( .A1(n11213), .A2(
        inner_first_stage_data_reg[808]), .B1(n11212), .B2(
        inner_first_stage_data_reg[904]), .ZN(n11120) );
  AOI22D1BWP30P140LVT U15764 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[1000]), .B1(n11217), .B2(
        inner_first_stage_data_reg[968]), .ZN(n11119) );
  ND4D1BWP30P140LVT U15765 ( .A1(n11122), .A2(n11121), .A3(n11120), .A4(n11119), .ZN(N7859) );
  AOI22D1BWP30P140LVT U15766 ( .A1(n11213), .A2(
        inner_first_stage_data_reg[809]), .B1(n11211), .B2(
        inner_first_stage_data_reg[841]), .ZN(n11126) );
  AOI22D1BWP30P140LVT U15767 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[777]), .B1(n11215), .B2(
        inner_first_stage_data_reg[937]), .ZN(n11125) );
  AOI22D1BWP30P140LVT U15768 ( .A1(n11216), .A2(
        inner_first_stage_data_reg[873]), .B1(n11212), .B2(
        inner_first_stage_data_reg[905]), .ZN(n11124) );
  AOI22D1BWP30P140LVT U15769 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[1001]), .B1(n11217), .B2(
        inner_first_stage_data_reg[969]), .ZN(n11123) );
  ND4D1BWP30P140LVT U15770 ( .A1(n11126), .A2(n11125), .A3(n11124), .A4(n11123), .ZN(N7860) );
  AOI22D1BWP30P140LVT U15771 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[778]), .B1(n11216), .B2(
        inner_first_stage_data_reg[874]), .ZN(n11130) );
  AOI22D1BWP30P140LVT U15772 ( .A1(n11213), .A2(
        inner_first_stage_data_reg[810]), .B1(n11211), .B2(
        inner_first_stage_data_reg[842]), .ZN(n11129) );
  AOI22D1BWP30P140LVT U15773 ( .A1(n11215), .A2(
        inner_first_stage_data_reg[938]), .B1(n11212), .B2(
        inner_first_stage_data_reg[906]), .ZN(n11128) );
  AOI22D1BWP30P140LVT U15774 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[1002]), .B1(n11217), .B2(
        inner_first_stage_data_reg[970]), .ZN(n11127) );
  ND4D1BWP30P140LVT U15775 ( .A1(n11130), .A2(n11129), .A3(n11128), .A4(n11127), .ZN(N7861) );
  AOI22D1BWP30P140LVT U15776 ( .A1(n11215), .A2(
        inner_first_stage_data_reg[939]), .B1(n11211), .B2(
        inner_first_stage_data_reg[843]), .ZN(n11134) );
  AOI22D1BWP30P140LVT U15777 ( .A1(n11216), .A2(
        inner_first_stage_data_reg[875]), .B1(n11212), .B2(
        inner_first_stage_data_reg[907]), .ZN(n11133) );
  AOI22D1BWP30P140LVT U15778 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[779]), .B1(n11213), .B2(
        inner_first_stage_data_reg[811]), .ZN(n11132) );
  AOI22D1BWP30P140LVT U15779 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[1003]), .B1(n11217), .B2(
        inner_first_stage_data_reg[971]), .ZN(n11131) );
  ND4D1BWP30P140LVT U15780 ( .A1(n11134), .A2(n11133), .A3(n11132), .A4(n11131), .ZN(N7862) );
  AOI22D1BWP30P140LVT U15781 ( .A1(n11212), .A2(
        inner_first_stage_data_reg[908]), .B1(n11211), .B2(
        inner_first_stage_data_reg[844]), .ZN(n11138) );
  AOI22D1BWP30P140LVT U15782 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[780]), .B1(n11216), .B2(
        inner_first_stage_data_reg[876]), .ZN(n11137) );
  AOI22D1BWP30P140LVT U15783 ( .A1(n11215), .A2(
        inner_first_stage_data_reg[940]), .B1(n11213), .B2(
        inner_first_stage_data_reg[812]), .ZN(n11136) );
  AOI22D1BWP30P140LVT U15784 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[1004]), .B1(n11217), .B2(
        inner_first_stage_data_reg[972]), .ZN(n11135) );
  ND4D1BWP30P140LVT U15785 ( .A1(n11138), .A2(n11137), .A3(n11136), .A4(n11135), .ZN(N7863) );
  AOI22D1BWP30P140LVT U15786 ( .A1(n11215), .A2(
        inner_first_stage_data_reg[941]), .B1(n11212), .B2(
        inner_first_stage_data_reg[909]), .ZN(n11142) );
  AOI22D1BWP30P140LVT U15787 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[781]), .B1(n11213), .B2(
        inner_first_stage_data_reg[813]), .ZN(n11141) );
  AOI22D1BWP30P140LVT U15788 ( .A1(n11216), .A2(
        inner_first_stage_data_reg[877]), .B1(n11211), .B2(
        inner_first_stage_data_reg[845]), .ZN(n11140) );
  AOI22D1BWP30P140LVT U15789 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[1005]), .B1(n11217), .B2(
        inner_first_stage_data_reg[973]), .ZN(n11139) );
  ND4D1BWP30P140LVT U15790 ( .A1(n11142), .A2(n11141), .A3(n11140), .A4(n11139), .ZN(N7864) );
  AOI22D1BWP30P140LVT U15791 ( .A1(n11216), .A2(
        inner_first_stage_data_reg[878]), .B1(n11213), .B2(
        inner_first_stage_data_reg[814]), .ZN(n11146) );
  AOI22D1BWP30P140LVT U15792 ( .A1(n11215), .A2(
        inner_first_stage_data_reg[942]), .B1(n11211), .B2(
        inner_first_stage_data_reg[846]), .ZN(n11145) );
  AOI22D1BWP30P140LVT U15793 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[782]), .B1(n11212), .B2(
        inner_first_stage_data_reg[910]), .ZN(n11144) );
  AOI22D1BWP30P140LVT U15794 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[1006]), .B1(n11217), .B2(
        inner_first_stage_data_reg[974]), .ZN(n11143) );
  ND4D1BWP30P140LVT U15795 ( .A1(n11146), .A2(n11145), .A3(n11144), .A4(n11143), .ZN(N7865) );
  AOI22D1BWP30P140LVT U15796 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[783]), .B1(n11215), .B2(
        inner_first_stage_data_reg[943]), .ZN(n11150) );
  AOI22D1BWP30P140LVT U15797 ( .A1(n11216), .A2(
        inner_first_stage_data_reg[879]), .B1(n11212), .B2(
        inner_first_stage_data_reg[911]), .ZN(n11149) );
  AOI22D1BWP30P140LVT U15798 ( .A1(n11213), .A2(
        inner_first_stage_data_reg[815]), .B1(n11211), .B2(
        inner_first_stage_data_reg[847]), .ZN(n11148) );
  AOI22D1BWP30P140LVT U15799 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[1007]), .B1(n11217), .B2(
        inner_first_stage_data_reg[975]), .ZN(n11147) );
  ND4D1BWP30P140LVT U15800 ( .A1(n11150), .A2(n11149), .A3(n11148), .A4(n11147), .ZN(N7866) );
  AOI22D1BWP30P140LVT U15801 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[784]), .B1(n11215), .B2(
        inner_first_stage_data_reg[944]), .ZN(n11154) );
  AOI22D1BWP30P140LVT U15802 ( .A1(n11216), .A2(
        inner_first_stage_data_reg[880]), .B1(n11211), .B2(
        inner_first_stage_data_reg[848]), .ZN(n11153) );
  AOI22D1BWP30P140LVT U15803 ( .A1(n11213), .A2(
        inner_first_stage_data_reg[816]), .B1(n11212), .B2(
        inner_first_stage_data_reg[912]), .ZN(n11152) );
  AOI22D1BWP30P140LVT U15804 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[1008]), .B1(n11217), .B2(
        inner_first_stage_data_reg[976]), .ZN(n11151) );
  ND4D1BWP30P140LVT U15805 ( .A1(n11154), .A2(n11153), .A3(n11152), .A4(n11151), .ZN(N7867) );
  AOI22D1BWP30P140LVT U15806 ( .A1(n11216), .A2(
        inner_first_stage_data_reg[881]), .B1(n11213), .B2(
        inner_first_stage_data_reg[817]), .ZN(n11158) );
  AOI22D1BWP30P140LVT U15807 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[785]), .B1(n11215), .B2(
        inner_first_stage_data_reg[945]), .ZN(n11157) );
  AOI22D1BWP30P140LVT U15808 ( .A1(n11212), .A2(
        inner_first_stage_data_reg[913]), .B1(n11211), .B2(
        inner_first_stage_data_reg[849]), .ZN(n11156) );
  AOI22D1BWP30P140LVT U15809 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[1009]), .B1(n11217), .B2(
        inner_first_stage_data_reg[977]), .ZN(n11155) );
  ND4D1BWP30P140LVT U15810 ( .A1(n11158), .A2(n11157), .A3(n11156), .A4(n11155), .ZN(N7868) );
  AOI22D1BWP30P140LVT U15811 ( .A1(n11215), .A2(
        inner_first_stage_data_reg[946]), .B1(n11212), .B2(
        inner_first_stage_data_reg[914]), .ZN(n11162) );
  AOI22D1BWP30P140LVT U15812 ( .A1(n11213), .A2(
        inner_first_stage_data_reg[818]), .B1(n11211), .B2(
        inner_first_stage_data_reg[850]), .ZN(n11161) );
  AOI22D1BWP30P140LVT U15813 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[786]), .B1(n11216), .B2(
        inner_first_stage_data_reg[882]), .ZN(n11160) );
  AOI22D1BWP30P140LVT U15814 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[1010]), .B1(n11217), .B2(
        inner_first_stage_data_reg[978]), .ZN(n11159) );
  ND4D1BWP30P140LVT U15815 ( .A1(n11162), .A2(n11161), .A3(n11160), .A4(n11159), .ZN(N7869) );
  AOI22D1BWP30P140LVT U15816 ( .A1(n11213), .A2(
        inner_first_stage_data_reg[819]), .B1(n11212), .B2(
        inner_first_stage_data_reg[915]), .ZN(n11166) );
  AOI22D1BWP30P140LVT U15817 ( .A1(n11216), .A2(
        inner_first_stage_data_reg[883]), .B1(n11215), .B2(
        inner_first_stage_data_reg[947]), .ZN(n11165) );
  AOI22D1BWP30P140LVT U15818 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[787]), .B1(n11211), .B2(
        inner_first_stage_data_reg[851]), .ZN(n11164) );
  AOI22D1BWP30P140LVT U15819 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[1011]), .B1(n11217), .B2(
        inner_first_stage_data_reg[979]), .ZN(n11163) );
  ND4D1BWP30P140LVT U15820 ( .A1(n11166), .A2(n11165), .A3(n11164), .A4(n11163), .ZN(N7870) );
  AOI22D1BWP30P140LVT U15821 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[788]), .B1(n11213), .B2(
        inner_first_stage_data_reg[820]), .ZN(n11170) );
  AOI22D1BWP30P140LVT U15822 ( .A1(n11216), .A2(
        inner_first_stage_data_reg[884]), .B1(n11212), .B2(
        inner_first_stage_data_reg[916]), .ZN(n11169) );
  AOI22D1BWP30P140LVT U15823 ( .A1(n11215), .A2(
        inner_first_stage_data_reg[948]), .B1(n11211), .B2(
        inner_first_stage_data_reg[852]), .ZN(n11168) );
  AOI22D1BWP30P140LVT U15824 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[1012]), .B1(n11217), .B2(
        inner_first_stage_data_reg[980]), .ZN(n11167) );
  ND4D1BWP30P140LVT U15825 ( .A1(n11170), .A2(n11169), .A3(n11168), .A4(n11167), .ZN(N7871) );
  AOI22D1BWP30P140LVT U15826 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[789]), .B1(n11212), .B2(
        inner_first_stage_data_reg[917]), .ZN(n11174) );
  AOI22D1BWP30P140LVT U15827 ( .A1(n11215), .A2(
        inner_first_stage_data_reg[949]), .B1(n11211), .B2(
        inner_first_stage_data_reg[853]), .ZN(n11173) );
  AOI22D1BWP30P140LVT U15828 ( .A1(n11216), .A2(
        inner_first_stage_data_reg[885]), .B1(n11213), .B2(
        inner_first_stage_data_reg[821]), .ZN(n11172) );
  AOI22D1BWP30P140LVT U15829 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[1013]), .B1(n11217), .B2(
        inner_first_stage_data_reg[981]), .ZN(n11171) );
  ND4D1BWP30P140LVT U15830 ( .A1(n11174), .A2(n11173), .A3(n11172), .A4(n11171), .ZN(N7872) );
  AOI22D1BWP30P140LVT U15831 ( .A1(n11216), .A2(
        inner_first_stage_data_reg[886]), .B1(n11215), .B2(
        inner_first_stage_data_reg[950]), .ZN(n11178) );
  AOI22D1BWP30P140LVT U15832 ( .A1(n11212), .A2(
        inner_first_stage_data_reg[918]), .B1(n11211), .B2(
        inner_first_stage_data_reg[854]), .ZN(n11177) );
  AOI22D1BWP30P140LVT U15833 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[790]), .B1(n11213), .B2(
        inner_first_stage_data_reg[822]), .ZN(n11176) );
  AOI22D1BWP30P140LVT U15834 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[1014]), .B1(n11217), .B2(
        inner_first_stage_data_reg[982]), .ZN(n11175) );
  ND4D1BWP30P140LVT U15835 ( .A1(n11178), .A2(n11177), .A3(n11176), .A4(n11175), .ZN(N7873) );
  AOI22D1BWP30P140LVT U15836 ( .A1(n11216), .A2(
        inner_first_stage_data_reg[887]), .B1(n11211), .B2(
        inner_first_stage_data_reg[855]), .ZN(n11182) );
  AOI22D1BWP30P140LVT U15837 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[791]), .B1(n11213), .B2(
        inner_first_stage_data_reg[823]), .ZN(n11181) );
  AOI22D1BWP30P140LVT U15838 ( .A1(n11215), .A2(
        inner_first_stage_data_reg[951]), .B1(n11212), .B2(
        inner_first_stage_data_reg[919]), .ZN(n11180) );
  AOI22D1BWP30P140LVT U15839 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[1015]), .B1(n11217), .B2(
        inner_first_stage_data_reg[983]), .ZN(n11179) );
  ND4D1BWP30P140LVT U15840 ( .A1(n11182), .A2(n11181), .A3(n11180), .A4(n11179), .ZN(N7874) );
  AOI22D1BWP30P140LVT U15841 ( .A1(n11213), .A2(
        inner_first_stage_data_reg[824]), .B1(n11212), .B2(
        inner_first_stage_data_reg[920]), .ZN(n11186) );
  AOI22D1BWP30P140LVT U15842 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[792]), .B1(n11216), .B2(
        inner_first_stage_data_reg[888]), .ZN(n11185) );
  AOI22D1BWP30P140LVT U15843 ( .A1(n11215), .A2(
        inner_first_stage_data_reg[952]), .B1(n11211), .B2(
        inner_first_stage_data_reg[856]), .ZN(n11184) );
  AOI22D1BWP30P140LVT U15844 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[1016]), .B1(n11217), .B2(
        inner_first_stage_data_reg[984]), .ZN(n11183) );
  ND4D1BWP30P140LVT U15845 ( .A1(n11186), .A2(n11185), .A3(n11184), .A4(n11183), .ZN(N7875) );
  AOI22D1BWP30P140LVT U15846 ( .A1(n11216), .A2(
        inner_first_stage_data_reg[889]), .B1(n11211), .B2(
        inner_first_stage_data_reg[857]), .ZN(n11190) );
  AOI22D1BWP30P140LVT U15847 ( .A1(n11215), .A2(
        inner_first_stage_data_reg[953]), .B1(n11213), .B2(
        inner_first_stage_data_reg[825]), .ZN(n11189) );
  AOI22D1BWP30P140LVT U15848 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[793]), .B1(n11212), .B2(
        inner_first_stage_data_reg[921]), .ZN(n11188) );
  AOI22D1BWP30P140LVT U15849 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[1017]), .B1(n11217), .B2(
        inner_first_stage_data_reg[985]), .ZN(n11187) );
  ND4D1BWP30P140LVT U15850 ( .A1(n11190), .A2(n11189), .A3(n11188), .A4(n11187), .ZN(N7876) );
  AOI22D1BWP30P140LVT U15851 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[794]), .B1(n11215), .B2(
        inner_first_stage_data_reg[954]), .ZN(n11194) );
  AOI22D1BWP30P140LVT U15852 ( .A1(n11216), .A2(
        inner_first_stage_data_reg[890]), .B1(n11211), .B2(
        inner_first_stage_data_reg[858]), .ZN(n11193) );
  AOI22D1BWP30P140LVT U15853 ( .A1(n11213), .A2(
        inner_first_stage_data_reg[826]), .B1(n11212), .B2(
        inner_first_stage_data_reg[922]), .ZN(n11192) );
  AOI22D1BWP30P140LVT U15854 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[1018]), .B1(n11217), .B2(
        inner_first_stage_data_reg[986]), .ZN(n11191) );
  ND4D1BWP30P140LVT U15855 ( .A1(n11194), .A2(n11193), .A3(n11192), .A4(n11191), .ZN(N7877) );
  AOI22D1BWP30P140LVT U15856 ( .A1(n11216), .A2(
        inner_first_stage_data_reg[891]), .B1(n11213), .B2(
        inner_first_stage_data_reg[827]), .ZN(n11198) );
  AOI22D1BWP30P140LVT U15857 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[795]), .B1(n11215), .B2(
        inner_first_stage_data_reg[955]), .ZN(n11197) );
  AOI22D1BWP30P140LVT U15858 ( .A1(n11212), .A2(
        inner_first_stage_data_reg[923]), .B1(n11211), .B2(
        inner_first_stage_data_reg[859]), .ZN(n11196) );
  AOI22D1BWP30P140LVT U15859 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[1019]), .B1(n11217), .B2(
        inner_first_stage_data_reg[987]), .ZN(n11195) );
  ND4D1BWP30P140LVT U15860 ( .A1(n11198), .A2(n11197), .A3(n11196), .A4(n11195), .ZN(N7878) );
  AOI22D1BWP30P140LVT U15861 ( .A1(n11213), .A2(
        inner_first_stage_data_reg[828]), .B1(n11212), .B2(
        inner_first_stage_data_reg[924]), .ZN(n11202) );
  AOI22D1BWP30P140LVT U15862 ( .A1(n11216), .A2(
        inner_first_stage_data_reg[892]), .B1(n11211), .B2(
        inner_first_stage_data_reg[860]), .ZN(n11201) );
  AOI22D1BWP30P140LVT U15863 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[796]), .B1(n11215), .B2(
        inner_first_stage_data_reg[956]), .ZN(n11200) );
  AOI22D1BWP30P140LVT U15864 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[1020]), .B1(n11217), .B2(
        inner_first_stage_data_reg[988]), .ZN(n11199) );
  ND4D1BWP30P140LVT U15865 ( .A1(n11202), .A2(n11201), .A3(n11200), .A4(n11199), .ZN(N7879) );
  AOI22D1BWP30P140LVT U15866 ( .A1(n11215), .A2(
        inner_first_stage_data_reg[957]), .B1(n11212), .B2(
        inner_first_stage_data_reg[925]), .ZN(n11206) );
  AOI22D1BWP30P140LVT U15867 ( .A1(n11216), .A2(
        inner_first_stage_data_reg[893]), .B1(n11211), .B2(
        inner_first_stage_data_reg[861]), .ZN(n11205) );
  AOI22D1BWP30P140LVT U15868 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[797]), .B1(n11213), .B2(
        inner_first_stage_data_reg[829]), .ZN(n11204) );
  AOI22D1BWP30P140LVT U15869 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[1021]), .B1(n11217), .B2(
        inner_first_stage_data_reg[989]), .ZN(n11203) );
  ND4D1BWP30P140LVT U15870 ( .A1(n11206), .A2(n11205), .A3(n11204), .A4(n11203), .ZN(N7880) );
  AOI22D1BWP30P140LVT U15871 ( .A1(n11213), .A2(
        inner_first_stage_data_reg[830]), .B1(n11212), .B2(
        inner_first_stage_data_reg[926]), .ZN(n11210) );
  AOI22D1BWP30P140LVT U15872 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[798]), .B1(n11215), .B2(
        inner_first_stage_data_reg[958]), .ZN(n11209) );
  AOI22D1BWP30P140LVT U15873 ( .A1(n11216), .A2(
        inner_first_stage_data_reg[894]), .B1(n11211), .B2(
        inner_first_stage_data_reg[862]), .ZN(n11208) );
  AOI22D1BWP30P140LVT U15874 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[1022]), .B1(n11217), .B2(
        inner_first_stage_data_reg[990]), .ZN(n11207) );
  ND4D1BWP30P140LVT U15875 ( .A1(n11210), .A2(n11209), .A3(n11208), .A4(n11207), .ZN(N7881) );
  AOI22D1BWP30P140LVT U15876 ( .A1(n11212), .A2(
        inner_first_stage_data_reg[927]), .B1(n11211), .B2(
        inner_first_stage_data_reg[863]), .ZN(n11222) );
  AOI22D1BWP30P140LVT U15877 ( .A1(n11214), .A2(
        inner_first_stage_data_reg[799]), .B1(n11213), .B2(
        inner_first_stage_data_reg[831]), .ZN(n11221) );
  AOI22D1BWP30P140LVT U15878 ( .A1(n11216), .A2(
        inner_first_stage_data_reg[895]), .B1(n11215), .B2(
        inner_first_stage_data_reg[959]), .ZN(n11220) );
  AOI22D1BWP30P140LVT U15879 ( .A1(n11218), .A2(
        inner_first_stage_data_reg[1023]), .B1(n11217), .B2(
        inner_first_stage_data_reg[991]), .ZN(n11219) );
  ND4D1BWP30P140LVT U15880 ( .A1(n11222), .A2(n11221), .A3(n11220), .A4(n11219), .ZN(N7882) );
  AOI22D1BWP30P140LVT U15881 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1184]), .B1(n11350), .B2(
        inner_first_stage_data_reg[1024]), .ZN(n11226) );
  AOI22D1BWP30P140LVT U15882 ( .A1(n11349), .A2(
        inner_first_stage_data_reg[1152]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1056]), .ZN(n11225) );
  AOI22D1BWP30P140LVT U15883 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1248]), .B1(n11353), .B2(
        inner_first_stage_data_reg[1088]), .ZN(n11224) );
  AOI22D1BWP30P140LVT U15884 ( .A1(n11352), .A2(
        inner_first_stage_data_reg[1120]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1216]), .ZN(n11223) );
  ND4D1BWP30P140LVT U15885 ( .A1(n11226), .A2(n11225), .A3(n11224), .A4(n11223), .ZN(N9725) );
  AOI22D1BWP30P140LVT U15886 ( .A1(n11350), .A2(
        inner_first_stage_data_reg[1025]), .B1(n11349), .B2(
        inner_first_stage_data_reg[1153]), .ZN(n11230) );
  AOI22D1BWP30P140LVT U15887 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1185]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1057]), .ZN(n11229) );
  AOI22D1BWP30P140LVT U15888 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1249]), .B1(n11352), .B2(
        inner_first_stage_data_reg[1121]), .ZN(n11228) );
  AOI22D1BWP30P140LVT U15889 ( .A1(n11353), .A2(
        inner_first_stage_data_reg[1089]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1217]), .ZN(n11227) );
  ND4D1BWP30P140LVT U15890 ( .A1(n11230), .A2(n11229), .A3(n11228), .A4(n11227), .ZN(N9726) );
  AOI22D1BWP30P140LVT U15891 ( .A1(n11350), .A2(
        inner_first_stage_data_reg[1026]), .B1(n11349), .B2(
        inner_first_stage_data_reg[1154]), .ZN(n11234) );
  AOI22D1BWP30P140LVT U15892 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1186]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1058]), .ZN(n11233) );
  AOI22D1BWP30P140LVT U15893 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1250]), .B1(n11352), .B2(
        inner_first_stage_data_reg[1122]), .ZN(n11232) );
  AOI22D1BWP30P140LVT U15894 ( .A1(n11353), .A2(
        inner_first_stage_data_reg[1090]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1218]), .ZN(n11231) );
  ND4D1BWP30P140LVT U15895 ( .A1(n11234), .A2(n11233), .A3(n11232), .A4(n11231), .ZN(N9727) );
  AOI22D1BWP30P140LVT U15896 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1187]), .B1(n11349), .B2(
        inner_first_stage_data_reg[1155]), .ZN(n11238) );
  AOI22D1BWP30P140LVT U15897 ( .A1(n11350), .A2(
        inner_first_stage_data_reg[1027]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1059]), .ZN(n11237) );
  AOI22D1BWP30P140LVT U15898 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1251]), .B1(n11353), .B2(
        inner_first_stage_data_reg[1091]), .ZN(n11236) );
  AOI22D1BWP30P140LVT U15899 ( .A1(n11352), .A2(
        inner_first_stage_data_reg[1123]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1219]), .ZN(n11235) );
  ND4D1BWP30P140LVT U15900 ( .A1(n11238), .A2(n11237), .A3(n11236), .A4(n11235), .ZN(N9728) );
  AOI22D1BWP30P140LVT U15901 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1188]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1060]), .ZN(n11242) );
  AOI22D1BWP30P140LVT U15902 ( .A1(n11350), .A2(
        inner_first_stage_data_reg[1028]), .B1(n11349), .B2(
        inner_first_stage_data_reg[1156]), .ZN(n11241) );
  AOI22D1BWP30P140LVT U15903 ( .A1(n11353), .A2(
        inner_first_stage_data_reg[1092]), .B1(n11352), .B2(
        inner_first_stage_data_reg[1124]), .ZN(n11240) );
  AOI22D1BWP30P140LVT U15904 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1252]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1220]), .ZN(n11239) );
  ND4D1BWP30P140LVT U15905 ( .A1(n11242), .A2(n11241), .A3(n11240), .A4(n11239), .ZN(N9729) );
  AOI22D1BWP30P140LVT U15906 ( .A1(n11350), .A2(
        inner_first_stage_data_reg[1029]), .B1(n11349), .B2(
        inner_first_stage_data_reg[1157]), .ZN(n11246) );
  AOI22D1BWP30P140LVT U15907 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1189]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1061]), .ZN(n11245) );
  AOI22D1BWP30P140LVT U15908 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1253]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1221]), .ZN(n11244) );
  AOI22D1BWP30P140LVT U15909 ( .A1(n11353), .A2(
        inner_first_stage_data_reg[1093]), .B1(n11352), .B2(
        inner_first_stage_data_reg[1125]), .ZN(n11243) );
  ND4D1BWP30P140LVT U15910 ( .A1(n11246), .A2(n11245), .A3(n11244), .A4(n11243), .ZN(N9730) );
  AOI22D1BWP30P140LVT U15911 ( .A1(n11350), .A2(
        inner_first_stage_data_reg[1030]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1062]), .ZN(n11250) );
  AOI22D1BWP30P140LVT U15912 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1190]), .B1(n11349), .B2(
        inner_first_stage_data_reg[1158]), .ZN(n11249) );
  AOI22D1BWP30P140LVT U15913 ( .A1(n11353), .A2(
        inner_first_stage_data_reg[1094]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1222]), .ZN(n11248) );
  AOI22D1BWP30P140LVT U15914 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1254]), .B1(n11352), .B2(
        inner_first_stage_data_reg[1126]), .ZN(n11247) );
  ND4D1BWP30P140LVT U15915 ( .A1(n11250), .A2(n11249), .A3(n11248), .A4(n11247), .ZN(N9731) );
  AOI22D1BWP30P140LVT U15916 ( .A1(n11349), .A2(
        inner_first_stage_data_reg[1159]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1063]), .ZN(n11254) );
  AOI22D1BWP30P140LVT U15917 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1191]), .B1(n11350), .B2(
        inner_first_stage_data_reg[1031]), .ZN(n11253) );
  AOI22D1BWP30P140LVT U15918 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1255]), .B1(n11352), .B2(
        inner_first_stage_data_reg[1127]), .ZN(n11252) );
  AOI22D1BWP30P140LVT U15919 ( .A1(n11353), .A2(
        inner_first_stage_data_reg[1095]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1223]), .ZN(n11251) );
  ND4D1BWP30P140LVT U15920 ( .A1(n11254), .A2(n11253), .A3(n11252), .A4(n11251), .ZN(N9732) );
  AOI22D1BWP30P140LVT U15921 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1192]), .B1(n11350), .B2(
        inner_first_stage_data_reg[1032]), .ZN(n11258) );
  AOI22D1BWP30P140LVT U15922 ( .A1(n11349), .A2(
        inner_first_stage_data_reg[1160]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1064]), .ZN(n11257) );
  AOI22D1BWP30P140LVT U15923 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1256]), .B1(n11352), .B2(
        inner_first_stage_data_reg[1128]), .ZN(n11256) );
  AOI22D1BWP30P140LVT U15924 ( .A1(n11353), .A2(
        inner_first_stage_data_reg[1096]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1224]), .ZN(n11255) );
  ND4D1BWP30P140LVT U15925 ( .A1(n11258), .A2(n11257), .A3(n11256), .A4(n11255), .ZN(N9733) );
  AOI22D1BWP30P140LVT U15926 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1193]), .B1(n11350), .B2(
        inner_first_stage_data_reg[1033]), .ZN(n11262) );
  AOI22D1BWP30P140LVT U15927 ( .A1(n11349), .A2(
        inner_first_stage_data_reg[1161]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1065]), .ZN(n11261) );
  AOI22D1BWP30P140LVT U15928 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1257]), .B1(n11352), .B2(
        inner_first_stage_data_reg[1129]), .ZN(n11260) );
  AOI22D1BWP30P140LVT U15929 ( .A1(n11353), .A2(
        inner_first_stage_data_reg[1097]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1225]), .ZN(n11259) );
  ND4D1BWP30P140LVT U15930 ( .A1(n11262), .A2(n11261), .A3(n11260), .A4(n11259), .ZN(N9734) );
  AOI22D1BWP30P140LVT U15931 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1194]), .B1(n11349), .B2(
        inner_first_stage_data_reg[1162]), .ZN(n11266) );
  AOI22D1BWP30P140LVT U15932 ( .A1(n11350), .A2(
        inner_first_stage_data_reg[1034]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1066]), .ZN(n11265) );
  AOI22D1BWP30P140LVT U15933 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1258]), .B1(n11353), .B2(
        inner_first_stage_data_reg[1098]), .ZN(n11264) );
  AOI22D1BWP30P140LVT U15934 ( .A1(n11352), .A2(
        inner_first_stage_data_reg[1130]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1226]), .ZN(n11263) );
  ND4D1BWP30P140LVT U15935 ( .A1(n11266), .A2(n11265), .A3(n11264), .A4(n11263), .ZN(N9735) );
  AOI22D1BWP30P140LVT U15936 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1195]), .B1(n11350), .B2(
        inner_first_stage_data_reg[1035]), .ZN(n11270) );
  AOI22D1BWP30P140LVT U15937 ( .A1(n11349), .A2(
        inner_first_stage_data_reg[1163]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1067]), .ZN(n11269) );
  AOI22D1BWP30P140LVT U15938 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1259]), .B1(n11353), .B2(
        inner_first_stage_data_reg[1099]), .ZN(n11268) );
  AOI22D1BWP30P140LVT U15939 ( .A1(n11352), .A2(
        inner_first_stage_data_reg[1131]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1227]), .ZN(n11267) );
  ND4D1BWP30P140LVT U15940 ( .A1(n11270), .A2(n11269), .A3(n11268), .A4(n11267), .ZN(N9736) );
  AOI22D1BWP30P140LVT U15941 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1196]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1068]), .ZN(n11274) );
  AOI22D1BWP30P140LVT U15942 ( .A1(n11350), .A2(
        inner_first_stage_data_reg[1036]), .B1(n11349), .B2(
        inner_first_stage_data_reg[1164]), .ZN(n11273) );
  AOI22D1BWP30P140LVT U15943 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1260]), .B1(n11353), .B2(
        inner_first_stage_data_reg[1100]), .ZN(n11272) );
  AOI22D1BWP30P140LVT U15944 ( .A1(n11352), .A2(
        inner_first_stage_data_reg[1132]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1228]), .ZN(n11271) );
  ND4D1BWP30P140LVT U15945 ( .A1(n11274), .A2(n11273), .A3(n11272), .A4(n11271), .ZN(N9737) );
  AOI22D1BWP30P140LVT U15946 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1197]), .B1(n11349), .B2(
        inner_first_stage_data_reg[1165]), .ZN(n11278) );
  AOI22D1BWP30P140LVT U15947 ( .A1(n11350), .A2(
        inner_first_stage_data_reg[1037]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1069]), .ZN(n11277) );
  AOI22D1BWP30P140LVT U15948 ( .A1(n11353), .A2(
        inner_first_stage_data_reg[1101]), .B1(n11352), .B2(
        inner_first_stage_data_reg[1133]), .ZN(n11276) );
  AOI22D1BWP30P140LVT U15949 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1261]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1229]), .ZN(n11275) );
  ND4D1BWP30P140LVT U15950 ( .A1(n11278), .A2(n11277), .A3(n11276), .A4(n11275), .ZN(N9738) );
  AOI22D1BWP30P140LVT U15951 ( .A1(n11350), .A2(
        inner_first_stage_data_reg[1038]), .B1(n11349), .B2(
        inner_first_stage_data_reg[1166]), .ZN(n11282) );
  AOI22D1BWP30P140LVT U15952 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1198]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1070]), .ZN(n11281) );
  AOI22D1BWP30P140LVT U15953 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1262]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1230]), .ZN(n11280) );
  AOI22D1BWP30P140LVT U15954 ( .A1(n11353), .A2(
        inner_first_stage_data_reg[1102]), .B1(n11352), .B2(
        inner_first_stage_data_reg[1134]), .ZN(n11279) );
  ND4D1BWP30P140LVT U15955 ( .A1(n11282), .A2(n11281), .A3(n11280), .A4(n11279), .ZN(N9739) );
  AOI22D1BWP30P140LVT U15956 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1199]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1071]), .ZN(n11286) );
  AOI22D1BWP30P140LVT U15957 ( .A1(n11350), .A2(
        inner_first_stage_data_reg[1039]), .B1(n11349), .B2(
        inner_first_stage_data_reg[1167]), .ZN(n11285) );
  AOI22D1BWP30P140LVT U15958 ( .A1(n11353), .A2(
        inner_first_stage_data_reg[1103]), .B1(n11352), .B2(
        inner_first_stage_data_reg[1135]), .ZN(n11284) );
  AOI22D1BWP30P140LVT U15959 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1263]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1231]), .ZN(n11283) );
  ND4D1BWP30P140LVT U15960 ( .A1(n11286), .A2(n11285), .A3(n11284), .A4(n11283), .ZN(N9740) );
  AOI22D1BWP30P140LVT U15961 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1200]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1072]), .ZN(n11290) );
  AOI22D1BWP30P140LVT U15962 ( .A1(n11350), .A2(
        inner_first_stage_data_reg[1040]), .B1(n11349), .B2(
        inner_first_stage_data_reg[1168]), .ZN(n11289) );
  AOI22D1BWP30P140LVT U15963 ( .A1(n11353), .A2(
        inner_first_stage_data_reg[1104]), .B1(n11352), .B2(
        inner_first_stage_data_reg[1136]), .ZN(n11288) );
  AOI22D1BWP30P140LVT U15964 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1264]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1232]), .ZN(n11287) );
  ND4D1BWP30P140LVT U15965 ( .A1(n11290), .A2(n11289), .A3(n11288), .A4(n11287), .ZN(N9741) );
  AOI22D1BWP30P140LVT U15966 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1201]), .B1(n11350), .B2(
        inner_first_stage_data_reg[1041]), .ZN(n11294) );
  AOI22D1BWP30P140LVT U15967 ( .A1(n11349), .A2(
        inner_first_stage_data_reg[1169]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1073]), .ZN(n11293) );
  AOI22D1BWP30P140LVT U15968 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1265]), .B1(n11353), .B2(
        inner_first_stage_data_reg[1105]), .ZN(n11292) );
  AOI22D1BWP30P140LVT U15969 ( .A1(n11352), .A2(
        inner_first_stage_data_reg[1137]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1233]), .ZN(n11291) );
  ND4D1BWP30P140LVT U15970 ( .A1(n11294), .A2(n11293), .A3(n11292), .A4(n11291), .ZN(N9742) );
  AOI22D1BWP30P140LVT U15971 ( .A1(n11350), .A2(
        inner_first_stage_data_reg[1042]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1074]), .ZN(n11298) );
  AOI22D1BWP30P140LVT U15972 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1202]), .B1(n11349), .B2(
        inner_first_stage_data_reg[1170]), .ZN(n11297) );
  AOI22D1BWP30P140LVT U15973 ( .A1(n11352), .A2(
        inner_first_stage_data_reg[1138]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1234]), .ZN(n11296) );
  AOI22D1BWP30P140LVT U15974 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1266]), .B1(n11353), .B2(
        inner_first_stage_data_reg[1106]), .ZN(n11295) );
  ND4D1BWP30P140LVT U15975 ( .A1(n11298), .A2(n11297), .A3(n11296), .A4(n11295), .ZN(N9743) );
  AOI22D1BWP30P140LVT U15976 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1203]), .B1(n11350), .B2(
        inner_first_stage_data_reg[1043]), .ZN(n11302) );
  AOI22D1BWP30P140LVT U15977 ( .A1(n11349), .A2(
        inner_first_stage_data_reg[1171]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1075]), .ZN(n11301) );
  AOI22D1BWP30P140LVT U15978 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1267]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1235]), .ZN(n11300) );
  AOI22D1BWP30P140LVT U15979 ( .A1(n11353), .A2(
        inner_first_stage_data_reg[1107]), .B1(n11352), .B2(
        inner_first_stage_data_reg[1139]), .ZN(n11299) );
  ND4D1BWP30P140LVT U15980 ( .A1(n11302), .A2(n11301), .A3(n11300), .A4(n11299), .ZN(N9744) );
  AOI22D1BWP30P140LVT U15981 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1204]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1076]), .ZN(n11306) );
  AOI22D1BWP30P140LVT U15982 ( .A1(n11350), .A2(
        inner_first_stage_data_reg[1044]), .B1(n11349), .B2(
        inner_first_stage_data_reg[1172]), .ZN(n11305) );
  AOI22D1BWP30P140LVT U15983 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1268]), .B1(n11353), .B2(
        inner_first_stage_data_reg[1108]), .ZN(n11304) );
  AOI22D1BWP30P140LVT U15984 ( .A1(n11352), .A2(
        inner_first_stage_data_reg[1140]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1236]), .ZN(n11303) );
  ND4D1BWP30P140LVT U15985 ( .A1(n11306), .A2(n11305), .A3(n11304), .A4(n11303), .ZN(N9745) );
  AOI22D1BWP30P140LVT U15986 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1205]), .B1(n11350), .B2(
        inner_first_stage_data_reg[1045]), .ZN(n11310) );
  AOI22D1BWP30P140LVT U15987 ( .A1(n11349), .A2(
        inner_first_stage_data_reg[1173]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1077]), .ZN(n11309) );
  AOI22D1BWP30P140LVT U15988 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1269]), .B1(n11353), .B2(
        inner_first_stage_data_reg[1109]), .ZN(n11308) );
  AOI22D1BWP30P140LVT U15989 ( .A1(n11352), .A2(
        inner_first_stage_data_reg[1141]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1237]), .ZN(n11307) );
  ND4D1BWP30P140LVT U15990 ( .A1(n11310), .A2(n11309), .A3(n11308), .A4(n11307), .ZN(N9746) );
  AOI22D1BWP30P140LVT U15991 ( .A1(n11349), .A2(
        inner_first_stage_data_reg[1174]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1078]), .ZN(n11314) );
  AOI22D1BWP30P140LVT U15992 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1206]), .B1(n11350), .B2(
        inner_first_stage_data_reg[1046]), .ZN(n11313) );
  AOI22D1BWP30P140LVT U15993 ( .A1(n11353), .A2(
        inner_first_stage_data_reg[1110]), .B1(n11352), .B2(
        inner_first_stage_data_reg[1142]), .ZN(n11312) );
  AOI22D1BWP30P140LVT U15994 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1270]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1238]), .ZN(n11311) );
  ND4D1BWP30P140LVT U15995 ( .A1(n11314), .A2(n11313), .A3(n11312), .A4(n11311), .ZN(N9747) );
  AOI22D1BWP30P140LVT U15996 ( .A1(n11350), .A2(
        inner_first_stage_data_reg[1047]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1079]), .ZN(n11318) );
  AOI22D1BWP30P140LVT U15997 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1207]), .B1(n11349), .B2(
        inner_first_stage_data_reg[1175]), .ZN(n11317) );
  AOI22D1BWP30P140LVT U15998 ( .A1(n11353), .A2(
        inner_first_stage_data_reg[1111]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1239]), .ZN(n11316) );
  AOI22D1BWP30P140LVT U15999 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1271]), .B1(n11352), .B2(
        inner_first_stage_data_reg[1143]), .ZN(n11315) );
  ND4D1BWP30P140LVT U16000 ( .A1(n11318), .A2(n11317), .A3(n11316), .A4(n11315), .ZN(N9748) );
  AOI22D1BWP30P140LVT U16001 ( .A1(n11349), .A2(
        inner_first_stage_data_reg[1176]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1080]), .ZN(n11322) );
  AOI22D1BWP30P140LVT U16002 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1208]), .B1(n11350), .B2(
        inner_first_stage_data_reg[1048]), .ZN(n11321) );
  AOI22D1BWP30P140LVT U16003 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1272]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1240]), .ZN(n11320) );
  AOI22D1BWP30P140LVT U16004 ( .A1(n11353), .A2(
        inner_first_stage_data_reg[1112]), .B1(n11352), .B2(
        inner_first_stage_data_reg[1144]), .ZN(n11319) );
  ND4D1BWP30P140LVT U16005 ( .A1(n11322), .A2(n11321), .A3(n11320), .A4(n11319), .ZN(N9749) );
  AOI22D1BWP30P140LVT U16006 ( .A1(n11350), .A2(
        inner_first_stage_data_reg[1049]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1081]), .ZN(n11326) );
  AOI22D1BWP30P140LVT U16007 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1209]), .B1(n11349), .B2(
        inner_first_stage_data_reg[1177]), .ZN(n11325) );
  AOI22D1BWP30P140LVT U16008 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1273]), .B1(n11353), .B2(
        inner_first_stage_data_reg[1113]), .ZN(n11324) );
  AOI22D1BWP30P140LVT U16009 ( .A1(n11352), .A2(
        inner_first_stage_data_reg[1145]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1241]), .ZN(n11323) );
  ND4D1BWP30P140LVT U16010 ( .A1(n11326), .A2(n11325), .A3(n11324), .A4(n11323), .ZN(N9750) );
  AOI22D1BWP30P140LVT U16011 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1210]), .B1(n11350), .B2(
        inner_first_stage_data_reg[1050]), .ZN(n11330) );
  AOI22D1BWP30P140LVT U16012 ( .A1(n11349), .A2(
        inner_first_stage_data_reg[1178]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1082]), .ZN(n11329) );
  AOI22D1BWP30P140LVT U16013 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1274]), .B1(n11352), .B2(
        inner_first_stage_data_reg[1146]), .ZN(n11328) );
  AOI22D1BWP30P140LVT U16014 ( .A1(n11353), .A2(
        inner_first_stage_data_reg[1114]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1242]), .ZN(n11327) );
  ND4D1BWP30P140LVT U16015 ( .A1(n11330), .A2(n11329), .A3(n11328), .A4(n11327), .ZN(N9751) );
  AOI22D1BWP30P140LVT U16016 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1211]), .B1(n11350), .B2(
        inner_first_stage_data_reg[1051]), .ZN(n11334) );
  AOI22D1BWP30P140LVT U16017 ( .A1(n11349), .A2(
        inner_first_stage_data_reg[1179]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1083]), .ZN(n11333) );
  AOI22D1BWP30P140LVT U16018 ( .A1(n11353), .A2(
        inner_first_stage_data_reg[1115]), .B1(n11352), .B2(
        inner_first_stage_data_reg[1147]), .ZN(n11332) );
  AOI22D1BWP30P140LVT U16019 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1275]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1243]), .ZN(n11331) );
  ND4D1BWP30P140LVT U16020 ( .A1(n11334), .A2(n11333), .A3(n11332), .A4(n11331), .ZN(N9752) );
  AOI22D1BWP30P140LVT U16021 ( .A1(n11350), .A2(
        inner_first_stage_data_reg[1052]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1084]), .ZN(n11338) );
  AOI22D1BWP30P140LVT U16022 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1212]), .B1(n11349), .B2(
        inner_first_stage_data_reg[1180]), .ZN(n11337) );
  AOI22D1BWP30P140LVT U16023 ( .A1(n11353), .A2(
        inner_first_stage_data_reg[1116]), .B1(n11352), .B2(
        inner_first_stage_data_reg[1148]), .ZN(n11336) );
  AOI22D1BWP30P140LVT U16024 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1276]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1244]), .ZN(n11335) );
  ND4D1BWP30P140LVT U16025 ( .A1(n11338), .A2(n11337), .A3(n11336), .A4(n11335), .ZN(N9753) );
  AOI22D1BWP30P140LVT U16026 ( .A1(n11350), .A2(
        inner_first_stage_data_reg[1053]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1085]), .ZN(n11343) );
  AOI22D1BWP30P140LVT U16027 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1213]), .B1(n11349), .B2(
        inner_first_stage_data_reg[1181]), .ZN(n11342) );
  AOI22D1BWP30P140LVT U16028 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1277]), .B1(n11352), .B2(
        inner_first_stage_data_reg[1149]), .ZN(n11341) );
  AOI22D1BWP30P140LVT U16029 ( .A1(n11353), .A2(
        inner_first_stage_data_reg[1117]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1245]), .ZN(n11340) );
  ND4D1BWP30P140LVT U16030 ( .A1(n11343), .A2(n11342), .A3(n11341), .A4(n11340), .ZN(N9754) );
  AOI22D1BWP30P140LVT U16031 ( .A1(n11350), .A2(
        inner_first_stage_data_reg[1054]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1086]), .ZN(n11347) );
  AOI22D1BWP30P140LVT U16032 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1214]), .B1(n11349), .B2(
        inner_first_stage_data_reg[1182]), .ZN(n11346) );
  AOI22D1BWP30P140LVT U16033 ( .A1(n11353), .A2(
        inner_first_stage_data_reg[1118]), .B1(n11352), .B2(
        inner_first_stage_data_reg[1150]), .ZN(n11345) );
  AOI22D1BWP30P140LVT U16034 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1278]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1246]), .ZN(n11344) );
  ND4D1BWP30P140LVT U16035 ( .A1(n11347), .A2(n11346), .A3(n11345), .A4(n11344), .ZN(N9755) );
  AOI22D1BWP30P140LVT U16036 ( .A1(n11348), .A2(
        inner_first_stage_data_reg[1215]), .B1(n11339), .B2(
        inner_first_stage_data_reg[1087]), .ZN(n11358) );
  AOI22D1BWP30P140LVT U16037 ( .A1(n11350), .A2(
        inner_first_stage_data_reg[1055]), .B1(n11349), .B2(
        inner_first_stage_data_reg[1183]), .ZN(n11357) );
  AOI22D1BWP30P140LVT U16038 ( .A1(n11352), .A2(
        inner_first_stage_data_reg[1151]), .B1(n11351), .B2(
        inner_first_stage_data_reg[1247]), .ZN(n11356) );
  AOI22D1BWP30P140LVT U16039 ( .A1(n11354), .A2(
        inner_first_stage_data_reg[1279]), .B1(n11353), .B2(
        inner_first_stage_data_reg[1119]), .ZN(n11355) );
  ND4D1BWP30P140LVT U16040 ( .A1(n11358), .A2(n11357), .A3(n11356), .A4(n11355), .ZN(N9756) );
  AOI22D1BWP30P140LVT U16041 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1440]), .B1(n11484), .B2(
        inner_first_stage_data_reg[1504]), .ZN(n11362) );
  AOI22D1BWP30P140LVT U16042 ( .A1(n11488), .A2(
        inner_first_stage_data_reg[1472]), .B1(n11485), .B2(
        inner_first_stage_data_reg[1408]), .ZN(n11361) );
  AOI22D1BWP30P140LVT U16043 ( .A1(n11487), .A2(
        inner_first_stage_data_reg[1312]), .B1(n11483), .B2(
        inner_first_stage_data_reg[1280]), .ZN(n11360) );
  AOI22D1BWP30P140LVT U16044 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1376]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1344]), .ZN(n11359) );
  ND4D1BWP30P140LVT U16045 ( .A1(n11362), .A2(n11361), .A3(n11360), .A4(n11359), .ZN(N11599) );
  AOI22D1BWP30P140LVT U16046 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1505]), .B1(n11485), .B2(
        inner_first_stage_data_reg[1409]), .ZN(n11366) );
  AOI22D1BWP30P140LVT U16047 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1441]), .B1(n11488), .B2(
        inner_first_stage_data_reg[1473]), .ZN(n11365) );
  AOI22D1BWP30P140LVT U16048 ( .A1(n11487), .A2(
        inner_first_stage_data_reg[1313]), .B1(n11483), .B2(
        inner_first_stage_data_reg[1281]), .ZN(n11364) );
  AOI22D1BWP30P140LVT U16049 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1377]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1345]), .ZN(n11363) );
  ND4D1BWP30P140LVT U16050 ( .A1(n11366), .A2(n11365), .A3(n11364), .A4(n11363), .ZN(N11600) );
  AOI22D1BWP30P140LVT U16051 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1506]), .B1(n11488), .B2(
        inner_first_stage_data_reg[1474]), .ZN(n11370) );
  AOI22D1BWP30P140LVT U16052 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1442]), .B1(n5893), .B2(
        inner_first_stage_data_reg[1282]), .ZN(n11369) );
  AOI22D1BWP30P140LVT U16053 ( .A1(n11485), .A2(
        inner_first_stage_data_reg[1410]), .B1(n11487), .B2(
        inner_first_stage_data_reg[1314]), .ZN(n11368) );
  AOI22D1BWP30P140LVT U16054 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1378]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1346]), .ZN(n11367) );
  ND4D1BWP30P140LVT U16055 ( .A1(n11370), .A2(n11369), .A3(n11368), .A4(n11367), .ZN(N11601) );
  AOI22D1BWP30P140LVT U16056 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1507]), .B1(n11488), .B2(
        inner_first_stage_data_reg[1475]), .ZN(n11374) );
  AOI22D1BWP30P140LVT U16057 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1443]), .B1(n11485), .B2(
        inner_first_stage_data_reg[1411]), .ZN(n11373) );
  AOI22D1BWP30P140LVT U16058 ( .A1(n11487), .A2(
        inner_first_stage_data_reg[1315]), .B1(n11483), .B2(
        inner_first_stage_data_reg[1283]), .ZN(n11372) );
  AOI22D1BWP30P140LVT U16059 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1379]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1347]), .ZN(n11371) );
  ND4D1BWP30P140LVT U16060 ( .A1(n11374), .A2(n11373), .A3(n11372), .A4(n11371), .ZN(N11602) );
  AOI22D1BWP30P140LVT U16061 ( .A1(n11488), .A2(
        inner_first_stage_data_reg[1476]), .B1(n11485), .B2(
        inner_first_stage_data_reg[1412]), .ZN(n11378) );
  AOI22D1BWP30P140LVT U16062 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1444]), .B1(n5892), .B2(
        inner_first_stage_data_reg[1284]), .ZN(n11377) );
  AOI22D1BWP30P140LVT U16063 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1508]), .B1(n11487), .B2(
        inner_first_stage_data_reg[1316]), .ZN(n11376) );
  AOI22D1BWP30P140LVT U16064 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1380]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1348]), .ZN(n11375) );
  ND4D1BWP30P140LVT U16065 ( .A1(n11378), .A2(n11377), .A3(n11376), .A4(n11375), .ZN(N11603) );
  AOI22D1BWP30P140LVT U16066 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1445]), .B1(n11485), .B2(
        inner_first_stage_data_reg[1413]), .ZN(n11382) );
  AOI22D1BWP30P140LVT U16067 ( .A1(n11488), .A2(
        inner_first_stage_data_reg[1477]), .B1(n11487), .B2(
        inner_first_stage_data_reg[1317]), .ZN(n11381) );
  AOI22D1BWP30P140LVT U16068 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1509]), .B1(n11483), .B2(
        inner_first_stage_data_reg[1285]), .ZN(n11380) );
  AOI22D1BWP30P140LVT U16069 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1381]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1349]), .ZN(n11379) );
  ND4D1BWP30P140LVT U16070 ( .A1(n11382), .A2(n11381), .A3(n11380), .A4(n11379), .ZN(N11604) );
  AOI22D1BWP30P140LVT U16071 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1510]), .B1(n11487), .B2(
        inner_first_stage_data_reg[1318]), .ZN(n11386) );
  AOI22D1BWP30P140LVT U16072 ( .A1(n11485), .A2(
        inner_first_stage_data_reg[1414]), .B1(n5893), .B2(
        inner_first_stage_data_reg[1286]), .ZN(n11385) );
  AOI22D1BWP30P140LVT U16073 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1446]), .B1(n11488), .B2(
        inner_first_stage_data_reg[1478]), .ZN(n11384) );
  AOI22D1BWP30P140LVT U16074 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1382]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1350]), .ZN(n11383) );
  ND4D1BWP30P140LVT U16075 ( .A1(n11386), .A2(n11385), .A3(n11384), .A4(n11383), .ZN(N11605) );
  AOI22D1BWP30P140LVT U16076 ( .A1(n11485), .A2(
        inner_first_stage_data_reg[1415]), .B1(n5893), .B2(
        inner_first_stage_data_reg[1287]), .ZN(n11390) );
  AOI22D1BWP30P140LVT U16077 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1447]), .B1(n11487), .B2(
        inner_first_stage_data_reg[1319]), .ZN(n11389) );
  AOI22D1BWP30P140LVT U16078 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1511]), .B1(n11488), .B2(
        inner_first_stage_data_reg[1479]), .ZN(n11388) );
  AOI22D1BWP30P140LVT U16079 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1383]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1351]), .ZN(n11387) );
  ND4D1BWP30P140LVT U16080 ( .A1(n11390), .A2(n11389), .A3(n11388), .A4(n11387), .ZN(N11606) );
  AOI22D1BWP30P140LVT U16081 ( .A1(n11488), .A2(
        inner_first_stage_data_reg[1480]), .B1(n5892), .B2(
        inner_first_stage_data_reg[1288]), .ZN(n11394) );
  AOI22D1BWP30P140LVT U16082 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1512]), .B1(n11487), .B2(
        inner_first_stage_data_reg[1320]), .ZN(n11393) );
  AOI22D1BWP30P140LVT U16083 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1448]), .B1(n11485), .B2(
        inner_first_stage_data_reg[1416]), .ZN(n11392) );
  AOI22D1BWP30P140LVT U16084 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1384]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1352]), .ZN(n11391) );
  ND4D1BWP30P140LVT U16085 ( .A1(n11394), .A2(n11393), .A3(n11392), .A4(n11391), .ZN(N11607) );
  AOI22D1BWP30P140LVT U16086 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1513]), .B1(n11488), .B2(
        inner_first_stage_data_reg[1481]), .ZN(n11398) );
  AOI22D1BWP30P140LVT U16087 ( .A1(n11487), .A2(
        inner_first_stage_data_reg[1321]), .B1(n5893), .B2(
        inner_first_stage_data_reg[1289]), .ZN(n11397) );
  AOI22D1BWP30P140LVT U16088 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1449]), .B1(n11485), .B2(
        inner_first_stage_data_reg[1417]), .ZN(n11396) );
  AOI22D1BWP30P140LVT U16089 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1385]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1353]), .ZN(n11395) );
  ND4D1BWP30P140LVT U16090 ( .A1(n11398), .A2(n11397), .A3(n11396), .A4(n11395), .ZN(N11608) );
  AOI22D1BWP30P140LVT U16091 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1450]), .B1(n11487), .B2(
        inner_first_stage_data_reg[1322]), .ZN(n11402) );
  AOI22D1BWP30P140LVT U16092 ( .A1(n11488), .A2(
        inner_first_stage_data_reg[1482]), .B1(n5892), .B2(
        inner_first_stage_data_reg[1290]), .ZN(n11401) );
  AOI22D1BWP30P140LVT U16093 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1514]), .B1(n11485), .B2(
        inner_first_stage_data_reg[1418]), .ZN(n11400) );
  AOI22D1BWP30P140LVT U16094 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1386]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1354]), .ZN(n11399) );
  ND4D1BWP30P140LVT U16095 ( .A1(n11402), .A2(n11401), .A3(n11400), .A4(n11399), .ZN(N11609) );
  AOI22D1BWP30P140LVT U16096 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1451]), .B1(n11488), .B2(
        inner_first_stage_data_reg[1483]), .ZN(n11406) );
  AOI22D1BWP30P140LVT U16097 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1515]), .B1(n5893), .B2(
        inner_first_stage_data_reg[1291]), .ZN(n11405) );
  AOI22D1BWP30P140LVT U16098 ( .A1(n11485), .A2(
        inner_first_stage_data_reg[1419]), .B1(n11487), .B2(
        inner_first_stage_data_reg[1323]), .ZN(n11404) );
  AOI22D1BWP30P140LVT U16099 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1387]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1355]), .ZN(n11403) );
  ND4D1BWP30P140LVT U16100 ( .A1(n11406), .A2(n11405), .A3(n11404), .A4(n11403), .ZN(N11610) );
  AOI22D1BWP30P140LVT U16101 ( .A1(n11487), .A2(
        inner_first_stage_data_reg[1324]), .B1(n5893), .B2(
        inner_first_stage_data_reg[1292]), .ZN(n11410) );
  AOI22D1BWP30P140LVT U16102 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1452]), .B1(n11484), .B2(
        inner_first_stage_data_reg[1516]), .ZN(n11409) );
  AOI22D1BWP30P140LVT U16103 ( .A1(n11488), .A2(
        inner_first_stage_data_reg[1484]), .B1(n11485), .B2(
        inner_first_stage_data_reg[1420]), .ZN(n11408) );
  AOI22D1BWP30P140LVT U16104 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1388]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1356]), .ZN(n11407) );
  ND4D1BWP30P140LVT U16105 ( .A1(n11410), .A2(n11409), .A3(n11408), .A4(n11407), .ZN(N11611) );
  AOI22D1BWP30P140LVT U16106 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1453]), .B1(n11487), .B2(
        inner_first_stage_data_reg[1325]), .ZN(n11414) );
  AOI22D1BWP30P140LVT U16107 ( .A1(n11485), .A2(
        inner_first_stage_data_reg[1421]), .B1(n5892), .B2(
        inner_first_stage_data_reg[1293]), .ZN(n11413) );
  AOI22D1BWP30P140LVT U16108 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1517]), .B1(n11488), .B2(
        inner_first_stage_data_reg[1485]), .ZN(n11412) );
  AOI22D1BWP30P140LVT U16109 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1389]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1357]), .ZN(n11411) );
  ND4D1BWP30P140LVT U16110 ( .A1(n11414), .A2(n11413), .A3(n11412), .A4(n11411), .ZN(N11612) );
  AOI22D1BWP30P140LVT U16111 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1454]), .B1(n11485), .B2(
        inner_first_stage_data_reg[1422]), .ZN(n11418) );
  AOI22D1BWP30P140LVT U16112 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1518]), .B1(n11488), .B2(
        inner_first_stage_data_reg[1486]), .ZN(n11417) );
  AOI22D1BWP30P140LVT U16113 ( .A1(n11487), .A2(
        inner_first_stage_data_reg[1326]), .B1(n11483), .B2(
        inner_first_stage_data_reg[1294]), .ZN(n11416) );
  AOI22D1BWP30P140LVT U16114 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1390]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1358]), .ZN(n11415) );
  ND4D1BWP30P140LVT U16115 ( .A1(n11418), .A2(n11417), .A3(n11416), .A4(n11415), .ZN(N11613) );
  AOI22D1BWP30P140LVT U16116 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1519]), .B1(n11488), .B2(
        inner_first_stage_data_reg[1487]), .ZN(n11422) );
  AOI22D1BWP30P140LVT U16117 ( .A1(n11485), .A2(
        inner_first_stage_data_reg[1423]), .B1(n11487), .B2(
        inner_first_stage_data_reg[1327]), .ZN(n11421) );
  AOI22D1BWP30P140LVT U16118 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1455]), .B1(n11483), .B2(
        inner_first_stage_data_reg[1295]), .ZN(n11420) );
  AOI22D1BWP30P140LVT U16119 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1391]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1359]), .ZN(n11419) );
  ND4D1BWP30P140LVT U16120 ( .A1(n11422), .A2(n11421), .A3(n11420), .A4(n11419), .ZN(N11614) );
  AOI22D1BWP30P140LVT U16121 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1520]), .B1(n11487), .B2(
        inner_first_stage_data_reg[1328]), .ZN(n11426) );
  AOI22D1BWP30P140LVT U16122 ( .A1(n11485), .A2(
        inner_first_stage_data_reg[1424]), .B1(n5892), .B2(
        inner_first_stage_data_reg[1296]), .ZN(n11425) );
  AOI22D1BWP30P140LVT U16123 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1456]), .B1(n11488), .B2(
        inner_first_stage_data_reg[1488]), .ZN(n11424) );
  AOI22D1BWP30P140LVT U16124 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1392]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1360]), .ZN(n11423) );
  ND4D1BWP30P140LVT U16125 ( .A1(n11426), .A2(n11425), .A3(n11424), .A4(n11423), .ZN(N11615) );
  AOI22D1BWP30P140LVT U16126 ( .A1(n11485), .A2(
        inner_first_stage_data_reg[1425]), .B1(n11487), .B2(
        inner_first_stage_data_reg[1329]), .ZN(n11430) );
  AOI22D1BWP30P140LVT U16127 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1521]), .B1(n5892), .B2(
        inner_first_stage_data_reg[1297]), .ZN(n11429) );
  AOI22D1BWP30P140LVT U16128 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1457]), .B1(n11488), .B2(
        inner_first_stage_data_reg[1489]), .ZN(n11428) );
  AOI22D1BWP30P140LVT U16129 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1393]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1361]), .ZN(n11427) );
  ND4D1BWP30P140LVT U16130 ( .A1(n11430), .A2(n11429), .A3(n11428), .A4(n11427), .ZN(N11616) );
  AOI22D1BWP30P140LVT U16131 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1458]), .B1(n11485), .B2(
        inner_first_stage_data_reg[1426]), .ZN(n11434) );
  AOI22D1BWP30P140LVT U16132 ( .A1(n11488), .A2(
        inner_first_stage_data_reg[1490]), .B1(n11487), .B2(
        inner_first_stage_data_reg[1330]), .ZN(n11433) );
  AOI22D1BWP30P140LVT U16133 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1522]), .B1(n11483), .B2(
        inner_first_stage_data_reg[1298]), .ZN(n11432) );
  AOI22D1BWP30P140LVT U16134 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1394]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1362]), .ZN(n11431) );
  ND4D1BWP30P140LVT U16135 ( .A1(n11434), .A2(n11433), .A3(n11432), .A4(n11431), .ZN(N11617) );
  AOI22D1BWP30P140LVT U16136 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1523]), .B1(n11485), .B2(
        inner_first_stage_data_reg[1427]), .ZN(n11438) );
  AOI22D1BWP30P140LVT U16137 ( .A1(n11487), .A2(
        inner_first_stage_data_reg[1331]), .B1(n5892), .B2(
        inner_first_stage_data_reg[1299]), .ZN(n11437) );
  AOI22D1BWP30P140LVT U16138 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1459]), .B1(n11488), .B2(
        inner_first_stage_data_reg[1491]), .ZN(n11436) );
  AOI22D1BWP30P140LVT U16139 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1395]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1363]), .ZN(n11435) );
  ND4D1BWP30P140LVT U16140 ( .A1(n11438), .A2(n11437), .A3(n11436), .A4(n11435), .ZN(N11618) );
  AOI22D1BWP30P140LVT U16141 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1460]), .B1(n11487), .B2(
        inner_first_stage_data_reg[1332]), .ZN(n11442) );
  AOI22D1BWP30P140LVT U16142 ( .A1(n11488), .A2(
        inner_first_stage_data_reg[1492]), .B1(n5892), .B2(
        inner_first_stage_data_reg[1300]), .ZN(n11441) );
  AOI22D1BWP30P140LVT U16143 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1524]), .B1(n11485), .B2(
        inner_first_stage_data_reg[1428]), .ZN(n11440) );
  AOI22D1BWP30P140LVT U16144 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1396]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1364]), .ZN(n11439) );
  ND4D1BWP30P140LVT U16145 ( .A1(n11442), .A2(n11441), .A3(n11440), .A4(n11439), .ZN(N11619) );
  AOI22D1BWP30P140LVT U16146 ( .A1(n11488), .A2(
        inner_first_stage_data_reg[1493]), .B1(n11485), .B2(
        inner_first_stage_data_reg[1429]), .ZN(n11446) );
  AOI22D1BWP30P140LVT U16147 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1461]), .B1(n5893), .B2(
        inner_first_stage_data_reg[1301]), .ZN(n11445) );
  AOI22D1BWP30P140LVT U16148 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1525]), .B1(n11487), .B2(
        inner_first_stage_data_reg[1333]), .ZN(n11444) );
  AOI22D1BWP30P140LVT U16149 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1397]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1365]), .ZN(n11443) );
  ND4D1BWP30P140LVT U16150 ( .A1(n11446), .A2(n11445), .A3(n11444), .A4(n11443), .ZN(N11620) );
  AOI22D1BWP30P140LVT U16151 ( .A1(n11485), .A2(
        inner_first_stage_data_reg[1430]), .B1(n5892), .B2(
        inner_first_stage_data_reg[1302]), .ZN(n11450) );
  AOI22D1BWP30P140LVT U16152 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1462]), .B1(n11487), .B2(
        inner_first_stage_data_reg[1334]), .ZN(n11449) );
  AOI22D1BWP30P140LVT U16153 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1526]), .B1(n11488), .B2(
        inner_first_stage_data_reg[1494]), .ZN(n11448) );
  AOI22D1BWP30P140LVT U16154 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1398]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1366]), .ZN(n11447) );
  ND4D1BWP30P140LVT U16155 ( .A1(n11450), .A2(n11449), .A3(n11448), .A4(n11447), .ZN(N11621) );
  AOI22D1BWP30P140LVT U16156 ( .A1(n11488), .A2(
        inner_first_stage_data_reg[1495]), .B1(n11487), .B2(
        inner_first_stage_data_reg[1335]), .ZN(n11454) );
  AOI22D1BWP30P140LVT U16157 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1463]), .B1(n11484), .B2(
        inner_first_stage_data_reg[1527]), .ZN(n11453) );
  AOI22D1BWP30P140LVT U16158 ( .A1(n11485), .A2(
        inner_first_stage_data_reg[1431]), .B1(n11483), .B2(
        inner_first_stage_data_reg[1303]), .ZN(n11452) );
  AOI22D1BWP30P140LVT U16159 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1399]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1367]), .ZN(n11451) );
  ND4D1BWP30P140LVT U16160 ( .A1(n11454), .A2(n11453), .A3(n11452), .A4(n11451), .ZN(N11622) );
  AOI22D1BWP30P140LVT U16161 ( .A1(n11485), .A2(
        inner_first_stage_data_reg[1432]), .B1(n11487), .B2(
        inner_first_stage_data_reg[1336]), .ZN(n11458) );
  AOI22D1BWP30P140LVT U16162 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1528]), .B1(n11488), .B2(
        inner_first_stage_data_reg[1496]), .ZN(n11457) );
  AOI22D1BWP30P140LVT U16163 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1464]), .B1(n11483), .B2(
        inner_first_stage_data_reg[1304]), .ZN(n11456) );
  AOI22D1BWP30P140LVT U16164 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1400]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1368]), .ZN(n11455) );
  ND4D1BWP30P140LVT U16165 ( .A1(n11458), .A2(n11457), .A3(n11456), .A4(n11455), .ZN(N11623) );
  AOI22D1BWP30P140LVT U16166 ( .A1(n11485), .A2(
        inner_first_stage_data_reg[1433]), .B1(n11487), .B2(
        inner_first_stage_data_reg[1337]), .ZN(n11462) );
  AOI22D1BWP30P140LVT U16167 ( .A1(n11488), .A2(
        inner_first_stage_data_reg[1497]), .B1(n5893), .B2(
        inner_first_stage_data_reg[1305]), .ZN(n11461) );
  AOI22D1BWP30P140LVT U16168 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1465]), .B1(n11484), .B2(
        inner_first_stage_data_reg[1529]), .ZN(n11460) );
  AOI22D1BWP30P140LVT U16169 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1401]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1369]), .ZN(n11459) );
  ND4D1BWP30P140LVT U16170 ( .A1(n11462), .A2(n11461), .A3(n11460), .A4(n11459), .ZN(N11624) );
  AOI22D1BWP30P140LVT U16171 ( .A1(n11485), .A2(
        inner_first_stage_data_reg[1434]), .B1(n11487), .B2(
        inner_first_stage_data_reg[1338]), .ZN(n11466) );
  AOI22D1BWP30P140LVT U16172 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1466]), .B1(n11484), .B2(
        inner_first_stage_data_reg[1530]), .ZN(n11465) );
  AOI22D1BWP30P140LVT U16173 ( .A1(n11488), .A2(
        inner_first_stage_data_reg[1498]), .B1(n11483), .B2(
        inner_first_stage_data_reg[1306]), .ZN(n11464) );
  AOI22D1BWP30P140LVT U16174 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1402]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1370]), .ZN(n11463) );
  ND4D1BWP30P140LVT U16175 ( .A1(n11466), .A2(n11465), .A3(n11464), .A4(n11463), .ZN(N11625) );
  AOI22D1BWP30P140LVT U16176 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1467]), .B1(n5892), .B2(
        inner_first_stage_data_reg[1307]), .ZN(n11470) );
  AOI22D1BWP30P140LVT U16177 ( .A1(n11485), .A2(
        inner_first_stage_data_reg[1435]), .B1(n11487), .B2(
        inner_first_stage_data_reg[1339]), .ZN(n11469) );
  AOI22D1BWP30P140LVT U16178 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1531]), .B1(n11488), .B2(
        inner_first_stage_data_reg[1499]), .ZN(n11468) );
  AOI22D1BWP30P140LVT U16179 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1403]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1371]), .ZN(n11467) );
  ND4D1BWP30P140LVT U16180 ( .A1(n11470), .A2(n11469), .A3(n11468), .A4(n11467), .ZN(N11626) );
  AOI22D1BWP30P140LVT U16181 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1532]), .B1(n11487), .B2(
        inner_first_stage_data_reg[1340]), .ZN(n11474) );
  AOI22D1BWP30P140LVT U16182 ( .A1(n11488), .A2(
        inner_first_stage_data_reg[1500]), .B1(n5893), .B2(
        inner_first_stage_data_reg[1308]), .ZN(n11473) );
  AOI22D1BWP30P140LVT U16183 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1468]), .B1(n11485), .B2(
        inner_first_stage_data_reg[1436]), .ZN(n11472) );
  AOI22D1BWP30P140LVT U16184 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1404]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1372]), .ZN(n11471) );
  ND4D1BWP30P140LVT U16185 ( .A1(n11474), .A2(n11473), .A3(n11472), .A4(n11471), .ZN(N11627) );
  AOI22D1BWP30P140LVT U16186 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1533]), .B1(n11485), .B2(
        inner_first_stage_data_reg[1437]), .ZN(n11478) );
  AOI22D1BWP30P140LVT U16187 ( .A1(n11488), .A2(
        inner_first_stage_data_reg[1501]), .B1(n5892), .B2(
        inner_first_stage_data_reg[1309]), .ZN(n11477) );
  AOI22D1BWP30P140LVT U16188 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1469]), .B1(n11487), .B2(
        inner_first_stage_data_reg[1341]), .ZN(n11476) );
  AOI22D1BWP30P140LVT U16189 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1405]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1373]), .ZN(n11475) );
  ND4D1BWP30P140LVT U16190 ( .A1(n11478), .A2(n11477), .A3(n11476), .A4(n11475), .ZN(N11628) );
  AOI22D1BWP30P140LVT U16191 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1534]), .B1(n11485), .B2(
        inner_first_stage_data_reg[1438]), .ZN(n11482) );
  AOI22D1BWP30P140LVT U16192 ( .A1(n11488), .A2(
        inner_first_stage_data_reg[1502]), .B1(n11487), .B2(
        inner_first_stage_data_reg[1342]), .ZN(n11481) );
  AOI22D1BWP30P140LVT U16193 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1470]), .B1(n11483), .B2(
        inner_first_stage_data_reg[1310]), .ZN(n11480) );
  AOI22D1BWP30P140LVT U16194 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1406]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1374]), .ZN(n11479) );
  ND4D1BWP30P140LVT U16195 ( .A1(n11482), .A2(n11481), .A3(n11480), .A4(n11479), .ZN(N11629) );
  AOI22D1BWP30P140LVT U16196 ( .A1(n11484), .A2(
        inner_first_stage_data_reg[1535]), .B1(n5893), .B2(
        inner_first_stage_data_reg[1311]), .ZN(n11494) );
  AOI22D1BWP30P140LVT U16197 ( .A1(n11486), .A2(
        inner_first_stage_data_reg[1471]), .B1(n11485), .B2(
        inner_first_stage_data_reg[1439]), .ZN(n11493) );
  AOI22D1BWP30P140LVT U16198 ( .A1(n11488), .A2(
        inner_first_stage_data_reg[1503]), .B1(n11487), .B2(
        inner_first_stage_data_reg[1343]), .ZN(n11492) );
  AOI22D1BWP30P140LVT U16199 ( .A1(n11490), .A2(
        inner_first_stage_data_reg[1407]), .B1(n11489), .B2(
        inner_first_stage_data_reg[1375]), .ZN(n11491) );
  ND4D1BWP30P140LVT U16200 ( .A1(n11494), .A2(n11493), .A3(n11492), .A4(n11491), .ZN(N11630) );
  AOI22D1BWP30P140LVT U16201 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1632]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1664]), .ZN(n11498) );
  AOI22D1BWP30P140LVT U16202 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1536]), .B1(n11621), .B2(
        inner_first_stage_data_reg[1696]), .ZN(n11497) );
  AOI22D1BWP30P140LVT U16203 ( .A1(n11624), .A2(
        inner_first_stage_data_reg[1600]), .B1(n11626), .B2(
        inner_first_stage_data_reg[1728]), .ZN(n11496) );
  AOI22D1BWP30P140LVT U16204 ( .A1(n11625), .A2(
        inner_first_stage_data_reg[1760]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1568]), .ZN(n11495) );
  ND4D1BWP30P140LVT U16205 ( .A1(n11498), .A2(n11497), .A3(n11496), .A4(n11495), .ZN(N13473) );
  AOI22D1BWP30P140LVT U16206 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1633]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1665]), .ZN(n11502) );
  AOI22D1BWP30P140LVT U16207 ( .A1(n11626), .A2(
        inner_first_stage_data_reg[1729]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1569]), .ZN(n11501) );
  AOI22D1BWP30P140LVT U16208 ( .A1(n11624), .A2(
        inner_first_stage_data_reg[1601]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1761]), .ZN(n11500) );
  AOI22D1BWP30P140LVT U16209 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1537]), .B1(n11621), .B2(
        inner_first_stage_data_reg[1697]), .ZN(n11499) );
  ND4D1BWP30P140LVT U16210 ( .A1(n11502), .A2(n11501), .A3(n11500), .A4(n11499), .ZN(N13474) );
  AOI22D1BWP30P140LVT U16211 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1634]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1666]), .ZN(n11506) );
  AOI22D1BWP30P140LVT U16212 ( .A1(n11621), .A2(
        inner_first_stage_data_reg[1698]), .B1(n11624), .B2(
        inner_first_stage_data_reg[1602]), .ZN(n11505) );
  AOI22D1BWP30P140LVT U16213 ( .A1(n11625), .A2(
        inner_first_stage_data_reg[1762]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1570]), .ZN(n11504) );
  AOI22D1BWP30P140LVT U16214 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1538]), .B1(n11626), .B2(
        inner_first_stage_data_reg[1730]), .ZN(n11503) );
  ND4D1BWP30P140LVT U16215 ( .A1(n11506), .A2(n11505), .A3(n11504), .A4(n11503), .ZN(N13475) );
  AOI22D1BWP30P140LVT U16216 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1635]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1667]), .ZN(n11510) );
  AOI22D1BWP30P140LVT U16217 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1539]), .B1(n11626), .B2(
        inner_first_stage_data_reg[1731]), .ZN(n11509) );
  AOI22D1BWP30P140LVT U16218 ( .A1(n11624), .A2(
        inner_first_stage_data_reg[1603]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1763]), .ZN(n11508) );
  AOI22D1BWP30P140LVT U16219 ( .A1(n11621), .A2(
        inner_first_stage_data_reg[1699]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1571]), .ZN(n11507) );
  ND4D1BWP30P140LVT U16220 ( .A1(n11510), .A2(n11509), .A3(n11508), .A4(n11507), .ZN(N13476) );
  AOI22D1BWP30P140LVT U16221 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1636]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1668]), .ZN(n11514) );
  AOI22D1BWP30P140LVT U16222 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1540]), .B1(n11624), .B2(
        inner_first_stage_data_reg[1604]), .ZN(n11513) );
  AOI22D1BWP30P140LVT U16223 ( .A1(n11625), .A2(
        inner_first_stage_data_reg[1764]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1572]), .ZN(n11512) );
  AOI22D1BWP30P140LVT U16224 ( .A1(n11621), .A2(
        inner_first_stage_data_reg[1700]), .B1(n11626), .B2(
        inner_first_stage_data_reg[1732]), .ZN(n11511) );
  ND4D1BWP30P140LVT U16225 ( .A1(n11514), .A2(n11513), .A3(n11512), .A4(n11511), .ZN(N13477) );
  AOI22D1BWP30P140LVT U16226 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1637]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1669]), .ZN(n11518) );
  AOI22D1BWP30P140LVT U16227 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1541]), .B1(n11624), .B2(
        inner_first_stage_data_reg[1605]), .ZN(n11517) );
  AOI22D1BWP30P140LVT U16228 ( .A1(n11626), .A2(
        inner_first_stage_data_reg[1733]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1765]), .ZN(n11516) );
  AOI22D1BWP30P140LVT U16229 ( .A1(n11621), .A2(
        inner_first_stage_data_reg[1701]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1573]), .ZN(n11515) );
  ND4D1BWP30P140LVT U16230 ( .A1(n11518), .A2(n11517), .A3(n11516), .A4(n11515), .ZN(N13478) );
  AOI22D1BWP30P140LVT U16231 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1638]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1670]), .ZN(n11522) );
  AOI22D1BWP30P140LVT U16232 ( .A1(n11626), .A2(
        inner_first_stage_data_reg[1734]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1574]), .ZN(n11521) );
  AOI22D1BWP30P140LVT U16233 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1542]), .B1(n11621), .B2(
        inner_first_stage_data_reg[1702]), .ZN(n11520) );
  AOI22D1BWP30P140LVT U16234 ( .A1(n11624), .A2(
        inner_first_stage_data_reg[1606]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1766]), .ZN(n11519) );
  ND4D1BWP30P140LVT U16235 ( .A1(n11522), .A2(n11521), .A3(n11520), .A4(n11519), .ZN(N13479) );
  AOI22D1BWP30P140LVT U16236 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1639]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1671]), .ZN(n11526) );
  AOI22D1BWP30P140LVT U16237 ( .A1(n11626), .A2(
        inner_first_stage_data_reg[1735]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1575]), .ZN(n11525) );
  AOI22D1BWP30P140LVT U16238 ( .A1(n11624), .A2(
        inner_first_stage_data_reg[1607]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1767]), .ZN(n11524) );
  AOI22D1BWP30P140LVT U16239 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1543]), .B1(n11621), .B2(
        inner_first_stage_data_reg[1703]), .ZN(n11523) );
  ND4D1BWP30P140LVT U16240 ( .A1(n11526), .A2(n11525), .A3(n11524), .A4(n11523), .ZN(N13480) );
  AOI22D1BWP30P140LVT U16241 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1640]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1672]), .ZN(n11530) );
  AOI22D1BWP30P140LVT U16242 ( .A1(n11621), .A2(
        inner_first_stage_data_reg[1704]), .B1(n11624), .B2(
        inner_first_stage_data_reg[1608]), .ZN(n11529) );
  AOI22D1BWP30P140LVT U16243 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1544]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1768]), .ZN(n11528) );
  AOI22D1BWP30P140LVT U16244 ( .A1(n11626), .A2(
        inner_first_stage_data_reg[1736]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1576]), .ZN(n11527) );
  ND4D1BWP30P140LVT U16245 ( .A1(n11530), .A2(n11529), .A3(n11528), .A4(n11527), .ZN(N13481) );
  AOI22D1BWP30P140LVT U16246 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1641]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1673]), .ZN(n11534) );
  AOI22D1BWP30P140LVT U16247 ( .A1(n11621), .A2(
        inner_first_stage_data_reg[1705]), .B1(n11624), .B2(
        inner_first_stage_data_reg[1609]), .ZN(n11533) );
  AOI22D1BWP30P140LVT U16248 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1545]), .B1(n11626), .B2(
        inner_first_stage_data_reg[1737]), .ZN(n11532) );
  AOI22D1BWP30P140LVT U16249 ( .A1(n11625), .A2(
        inner_first_stage_data_reg[1769]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1577]), .ZN(n11531) );
  ND4D1BWP30P140LVT U16250 ( .A1(n11534), .A2(n11533), .A3(n11532), .A4(n11531), .ZN(N13482) );
  AOI22D1BWP30P140LVT U16251 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1642]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1674]), .ZN(n11538) );
  AOI22D1BWP30P140LVT U16252 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1546]), .B1(n11626), .B2(
        inner_first_stage_data_reg[1738]), .ZN(n11537) );
  AOI22D1BWP30P140LVT U16253 ( .A1(n11624), .A2(
        inner_first_stage_data_reg[1610]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1770]), .ZN(n11536) );
  AOI22D1BWP30P140LVT U16254 ( .A1(n11621), .A2(
        inner_first_stage_data_reg[1706]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1578]), .ZN(n11535) );
  ND4D1BWP30P140LVT U16255 ( .A1(n11538), .A2(n11537), .A3(n11536), .A4(n11535), .ZN(N13483) );
  AOI22D1BWP30P140LVT U16256 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1643]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1675]), .ZN(n11542) );
  AOI22D1BWP30P140LVT U16257 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1547]), .B1(n11624), .B2(
        inner_first_stage_data_reg[1611]), .ZN(n11541) );
  AOI22D1BWP30P140LVT U16258 ( .A1(n11626), .A2(
        inner_first_stage_data_reg[1739]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1771]), .ZN(n11540) );
  AOI22D1BWP30P140LVT U16259 ( .A1(n11621), .A2(
        inner_first_stage_data_reg[1707]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1579]), .ZN(n11539) );
  ND4D1BWP30P140LVT U16260 ( .A1(n11542), .A2(n11541), .A3(n11540), .A4(n11539), .ZN(N13484) );
  AOI22D1BWP30P140LVT U16261 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1644]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1676]), .ZN(n11546) );
  AOI22D1BWP30P140LVT U16262 ( .A1(n11625), .A2(
        inner_first_stage_data_reg[1772]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1580]), .ZN(n11545) );
  AOI22D1BWP30P140LVT U16263 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1548]), .B1(n11621), .B2(
        inner_first_stage_data_reg[1708]), .ZN(n11544) );
  AOI22D1BWP30P140LVT U16264 ( .A1(n11624), .A2(
        inner_first_stage_data_reg[1612]), .B1(n11626), .B2(
        inner_first_stage_data_reg[1740]), .ZN(n11543) );
  ND4D1BWP30P140LVT U16265 ( .A1(n11546), .A2(n11545), .A3(n11544), .A4(n11543), .ZN(N13485) );
  AOI22D1BWP30P140LVT U16266 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1645]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1677]), .ZN(n11550) );
  AOI22D1BWP30P140LVT U16267 ( .A1(n11624), .A2(
        inner_first_stage_data_reg[1613]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1773]), .ZN(n11549) );
  AOI22D1BWP30P140LVT U16268 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1549]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1581]), .ZN(n11548) );
  AOI22D1BWP30P140LVT U16269 ( .A1(n11621), .A2(
        inner_first_stage_data_reg[1709]), .B1(n11626), .B2(
        inner_first_stage_data_reg[1741]), .ZN(n11547) );
  ND4D1BWP30P140LVT U16270 ( .A1(n11550), .A2(n11549), .A3(n11548), .A4(n11547), .ZN(N13486) );
  AOI22D1BWP30P140LVT U16271 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1646]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1678]), .ZN(n11554) );
  AOI22D1BWP30P140LVT U16272 ( .A1(n11624), .A2(
        inner_first_stage_data_reg[1614]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1582]), .ZN(n11553) );
  AOI22D1BWP30P140LVT U16273 ( .A1(n11621), .A2(
        inner_first_stage_data_reg[1710]), .B1(n11626), .B2(
        inner_first_stage_data_reg[1742]), .ZN(n11552) );
  AOI22D1BWP30P140LVT U16274 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1550]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1774]), .ZN(n11551) );
  ND4D1BWP30P140LVT U16275 ( .A1(n11554), .A2(n11553), .A3(n11552), .A4(n11551), .ZN(N13487) );
  AOI22D1BWP30P140LVT U16276 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1647]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1679]), .ZN(n11558) );
  AOI22D1BWP30P140LVT U16277 ( .A1(n11621), .A2(
        inner_first_stage_data_reg[1711]), .B1(n11624), .B2(
        inner_first_stage_data_reg[1615]), .ZN(n11557) );
  AOI22D1BWP30P140LVT U16278 ( .A1(n11626), .A2(
        inner_first_stage_data_reg[1743]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1583]), .ZN(n11556) );
  AOI22D1BWP30P140LVT U16279 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1551]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1775]), .ZN(n11555) );
  ND4D1BWP30P140LVT U16280 ( .A1(n11558), .A2(n11557), .A3(n11556), .A4(n11555), .ZN(N13488) );
  AOI22D1BWP30P140LVT U16281 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1648]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1680]), .ZN(n11562) );
  AOI22D1BWP30P140LVT U16282 ( .A1(n11624), .A2(
        inner_first_stage_data_reg[1616]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1776]), .ZN(n11561) );
  AOI22D1BWP30P140LVT U16283 ( .A1(n11621), .A2(
        inner_first_stage_data_reg[1712]), .B1(n11626), .B2(
        inner_first_stage_data_reg[1744]), .ZN(n11560) );
  AOI22D1BWP30P140LVT U16284 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1552]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1584]), .ZN(n11559) );
  ND4D1BWP30P140LVT U16285 ( .A1(n11562), .A2(n11561), .A3(n11560), .A4(n11559), .ZN(N13489) );
  AOI22D1BWP30P140LVT U16286 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1649]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1681]), .ZN(n11566) );
  AOI22D1BWP30P140LVT U16287 ( .A1(n11624), .A2(
        inner_first_stage_data_reg[1617]), .B1(n11626), .B2(
        inner_first_stage_data_reg[1745]), .ZN(n11565) );
  AOI22D1BWP30P140LVT U16288 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1553]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1585]), .ZN(n11564) );
  AOI22D1BWP30P140LVT U16289 ( .A1(n11621), .A2(
        inner_first_stage_data_reg[1713]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1777]), .ZN(n11563) );
  ND4D1BWP30P140LVT U16290 ( .A1(n11566), .A2(n11565), .A3(n11564), .A4(n11563), .ZN(N13490) );
  AOI22D1BWP30P140LVT U16291 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1650]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1682]), .ZN(n11570) );
  AOI22D1BWP30P140LVT U16292 ( .A1(n11621), .A2(
        inner_first_stage_data_reg[1714]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1778]), .ZN(n11569) );
  AOI22D1BWP30P140LVT U16293 ( .A1(n11624), .A2(
        inner_first_stage_data_reg[1618]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1586]), .ZN(n11568) );
  AOI22D1BWP30P140LVT U16294 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1554]), .B1(n11626), .B2(
        inner_first_stage_data_reg[1746]), .ZN(n11567) );
  ND4D1BWP30P140LVT U16295 ( .A1(n11570), .A2(n11569), .A3(n11568), .A4(n11567), .ZN(N13491) );
  AOI22D1BWP30P140LVT U16296 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1651]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1683]), .ZN(n11574) );
  AOI22D1BWP30P140LVT U16297 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1555]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1779]), .ZN(n11573) );
  AOI22D1BWP30P140LVT U16298 ( .A1(n11621), .A2(
        inner_first_stage_data_reg[1715]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1587]), .ZN(n11572) );
  AOI22D1BWP30P140LVT U16299 ( .A1(n11624), .A2(
        inner_first_stage_data_reg[1619]), .B1(n11626), .B2(
        inner_first_stage_data_reg[1747]), .ZN(n11571) );
  ND4D1BWP30P140LVT U16300 ( .A1(n11574), .A2(n11573), .A3(n11572), .A4(n11571), .ZN(N13492) );
  AOI22D1BWP30P140LVT U16301 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1652]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1684]), .ZN(n11578) );
  AOI22D1BWP30P140LVT U16302 ( .A1(n11621), .A2(
        inner_first_stage_data_reg[1716]), .B1(n11624), .B2(
        inner_first_stage_data_reg[1620]), .ZN(n11577) );
  AOI22D1BWP30P140LVT U16303 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1556]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1780]), .ZN(n11576) );
  AOI22D1BWP30P140LVT U16304 ( .A1(n11626), .A2(
        inner_first_stage_data_reg[1748]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1588]), .ZN(n11575) );
  ND4D1BWP30P140LVT U16305 ( .A1(n11578), .A2(n11577), .A3(n11576), .A4(n11575), .ZN(N13493) );
  AOI22D1BWP30P140LVT U16306 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1653]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1685]), .ZN(n11582) );
  AOI22D1BWP30P140LVT U16307 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1557]), .B1(n11626), .B2(
        inner_first_stage_data_reg[1749]), .ZN(n11581) );
  AOI22D1BWP30P140LVT U16308 ( .A1(n11624), .A2(
        inner_first_stage_data_reg[1621]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1781]), .ZN(n11580) );
  AOI22D1BWP30P140LVT U16309 ( .A1(n11621), .A2(
        inner_first_stage_data_reg[1717]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1589]), .ZN(n11579) );
  ND4D1BWP30P140LVT U16310 ( .A1(n11582), .A2(n11581), .A3(n11580), .A4(n11579), .ZN(N13494) );
  AOI22D1BWP30P140LVT U16311 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1654]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1686]), .ZN(n11586) );
  AOI22D1BWP30P140LVT U16312 ( .A1(n11621), .A2(
        inner_first_stage_data_reg[1718]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1782]), .ZN(n11585) );
  AOI22D1BWP30P140LVT U16313 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1558]), .B1(n11626), .B2(
        inner_first_stage_data_reg[1750]), .ZN(n11584) );
  AOI22D1BWP30P140LVT U16314 ( .A1(n11624), .A2(
        inner_first_stage_data_reg[1622]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1590]), .ZN(n11583) );
  ND4D1BWP30P140LVT U16315 ( .A1(n11586), .A2(n11585), .A3(n11584), .A4(n11583), .ZN(N13495) );
  AOI22D1BWP30P140LVT U16316 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1655]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1687]), .ZN(n11590) );
  AOI22D1BWP30P140LVT U16317 ( .A1(n11624), .A2(
        inner_first_stage_data_reg[1623]), .B1(n11626), .B2(
        inner_first_stage_data_reg[1751]), .ZN(n11589) );
  AOI22D1BWP30P140LVT U16318 ( .A1(n11621), .A2(
        inner_first_stage_data_reg[1719]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1783]), .ZN(n11588) );
  AOI22D1BWP30P140LVT U16319 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1559]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1591]), .ZN(n11587) );
  ND4D1BWP30P140LVT U16320 ( .A1(n11590), .A2(n11589), .A3(n11588), .A4(n11587), .ZN(N13496) );
  AOI22D1BWP30P140LVT U16321 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1656]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1688]), .ZN(n11594) );
  AOI22D1BWP30P140LVT U16322 ( .A1(n11624), .A2(
        inner_first_stage_data_reg[1624]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1592]), .ZN(n11593) );
  AOI22D1BWP30P140LVT U16323 ( .A1(n11621), .A2(
        inner_first_stage_data_reg[1720]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1784]), .ZN(n11592) );
  AOI22D1BWP30P140LVT U16324 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1560]), .B1(n11626), .B2(
        inner_first_stage_data_reg[1752]), .ZN(n11591) );
  ND4D1BWP30P140LVT U16325 ( .A1(n11594), .A2(n11593), .A3(n11592), .A4(n11591), .ZN(N13497) );
  AOI22D1BWP30P140LVT U16326 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1657]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1689]), .ZN(n11598) );
  AOI22D1BWP30P140LVT U16327 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1561]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1593]), .ZN(n11597) );
  AOI22D1BWP30P140LVT U16328 ( .A1(n11624), .A2(
        inner_first_stage_data_reg[1625]), .B1(n11626), .B2(
        inner_first_stage_data_reg[1753]), .ZN(n11596) );
  AOI22D1BWP30P140LVT U16329 ( .A1(n11621), .A2(
        inner_first_stage_data_reg[1721]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1785]), .ZN(n11595) );
  ND4D1BWP30P140LVT U16330 ( .A1(n11598), .A2(n11597), .A3(n11596), .A4(n11595), .ZN(N13498) );
  AOI22D1BWP30P140LVT U16331 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1658]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1690]), .ZN(n11602) );
  AOI22D1BWP30P140LVT U16332 ( .A1(n11621), .A2(
        inner_first_stage_data_reg[1722]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1786]), .ZN(n11601) );
  AOI22D1BWP30P140LVT U16333 ( .A1(n11624), .A2(
        inner_first_stage_data_reg[1626]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1594]), .ZN(n11600) );
  AOI22D1BWP30P140LVT U16334 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1562]), .B1(n11626), .B2(
        inner_first_stage_data_reg[1754]), .ZN(n11599) );
  ND4D1BWP30P140LVT U16335 ( .A1(n11602), .A2(n11601), .A3(n11600), .A4(n11599), .ZN(N13499) );
  AOI22D1BWP30P140LVT U16336 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1659]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1691]), .ZN(n11606) );
  AOI22D1BWP30P140LVT U16337 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1563]), .B1(n11624), .B2(
        inner_first_stage_data_reg[1627]), .ZN(n11605) );
  AOI22D1BWP30P140LVT U16338 ( .A1(n11621), .A2(
        inner_first_stage_data_reg[1723]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1787]), .ZN(n11604) );
  AOI22D1BWP30P140LVT U16339 ( .A1(n11626), .A2(
        inner_first_stage_data_reg[1755]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1595]), .ZN(n11603) );
  ND4D1BWP30P140LVT U16340 ( .A1(n11606), .A2(n11605), .A3(n11604), .A4(n11603), .ZN(N13500) );
  AOI22D1BWP30P140LVT U16341 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1660]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1692]), .ZN(n11610) );
  AOI22D1BWP30P140LVT U16342 ( .A1(n11621), .A2(
        inner_first_stage_data_reg[1724]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1596]), .ZN(n11609) );
  AOI22D1BWP30P140LVT U16343 ( .A1(n11624), .A2(
        inner_first_stage_data_reg[1628]), .B1(n11626), .B2(
        inner_first_stage_data_reg[1756]), .ZN(n11608) );
  AOI22D1BWP30P140LVT U16344 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1564]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1788]), .ZN(n11607) );
  ND4D1BWP30P140LVT U16345 ( .A1(n11610), .A2(n11609), .A3(n11608), .A4(n11607), .ZN(N13501) );
  AOI22D1BWP30P140LVT U16346 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1661]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1693]), .ZN(n11614) );
  AOI22D1BWP30P140LVT U16347 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1565]), .B1(n11621), .B2(
        inner_first_stage_data_reg[1725]), .ZN(n11613) );
  AOI22D1BWP30P140LVT U16348 ( .A1(n11624), .A2(
        inner_first_stage_data_reg[1629]), .B1(n11626), .B2(
        inner_first_stage_data_reg[1757]), .ZN(n11612) );
  AOI22D1BWP30P140LVT U16349 ( .A1(n11625), .A2(
        inner_first_stage_data_reg[1789]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1597]), .ZN(n11611) );
  ND4D1BWP30P140LVT U16350 ( .A1(n11614), .A2(n11613), .A3(n11612), .A4(n11611), .ZN(N13502) );
  AOI22D1BWP30P140LVT U16351 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1662]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1694]), .ZN(n11618) );
  AOI22D1BWP30P140LVT U16352 ( .A1(n11624), .A2(
        inner_first_stage_data_reg[1630]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1790]), .ZN(n11617) );
  AOI22D1BWP30P140LVT U16353 ( .A1(n11621), .A2(
        inner_first_stage_data_reg[1726]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1598]), .ZN(n11616) );
  AOI22D1BWP30P140LVT U16354 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1566]), .B1(n11626), .B2(
        inner_first_stage_data_reg[1758]), .ZN(n11615) );
  ND4D1BWP30P140LVT U16355 ( .A1(n11618), .A2(n11617), .A3(n11616), .A4(n11615), .ZN(N13503) );
  AOI22D1BWP30P140LVT U16356 ( .A1(n11620), .A2(
        inner_first_stage_data_reg[1663]), .B1(n11619), .B2(
        inner_first_stage_data_reg[1695]), .ZN(n11630) );
  AOI22D1BWP30P140LVT U16357 ( .A1(n11622), .A2(
        inner_first_stage_data_reg[1567]), .B1(n11621), .B2(
        inner_first_stage_data_reg[1727]), .ZN(n11629) );
  AOI22D1BWP30P140LVT U16358 ( .A1(n11624), .A2(
        inner_first_stage_data_reg[1631]), .B1(n11623), .B2(
        inner_first_stage_data_reg[1599]), .ZN(n11628) );
  AOI22D1BWP30P140LVT U16359 ( .A1(n11626), .A2(
        inner_first_stage_data_reg[1759]), .B1(n11625), .B2(
        inner_first_stage_data_reg[1791]), .ZN(n11627) );
  ND4D1BWP30P140LVT U16360 ( .A1(n11630), .A2(n11629), .A3(n11628), .A4(n11627), .ZN(N13504) );
  AOI22D1BWP30P140LVT U16361 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1952]), .B1(n11758), .B2(
        inner_first_stage_data_reg[1792]), .ZN(n11634) );
  AOI22D1BWP30P140LVT U16362 ( .A1(n11760), .A2(
        inner_first_stage_data_reg[1856]), .B1(n11757), .B2(
        inner_first_stage_data_reg[1920]), .ZN(n11633) );
  AOI22D1BWP30P140LVT U16363 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[1888]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1824]), .ZN(n11632) );
  AOI22D1BWP30P140LVT U16364 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[1984]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2016]), .ZN(n11631) );
  ND4D1BWP30P140LVT U16365 ( .A1(n11634), .A2(n11633), .A3(n11632), .A4(n11631), .ZN(N15347) );
  AOI22D1BWP30P140LVT U16366 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1953]), .B1(n11757), .B2(
        inner_first_stage_data_reg[1921]), .ZN(n11638) );
  AOI22D1BWP30P140LVT U16367 ( .A1(n11760), .A2(
        inner_first_stage_data_reg[1857]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1825]), .ZN(n11637) );
  AOI22D1BWP30P140LVT U16368 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1793]), .B1(n11755), .B2(
        inner_first_stage_data_reg[1889]), .ZN(n11636) );
  AOI22D1BWP30P140LVT U16369 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[1985]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2017]), .ZN(n11635) );
  ND4D1BWP30P140LVT U16370 ( .A1(n11638), .A2(n11637), .A3(n11636), .A4(n11635), .ZN(N15348) );
  AOI22D1BWP30P140LVT U16371 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1794]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1826]), .ZN(n11642) );
  AOI22D1BWP30P140LVT U16372 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1954]), .B1(n11760), .B2(
        inner_first_stage_data_reg[1858]), .ZN(n11641) );
  AOI22D1BWP30P140LVT U16373 ( .A1(n11757), .A2(
        inner_first_stage_data_reg[1922]), .B1(n11755), .B2(
        inner_first_stage_data_reg[1890]), .ZN(n11640) );
  AOI22D1BWP30P140LVT U16374 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[1986]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2018]), .ZN(n11639) );
  ND4D1BWP30P140LVT U16375 ( .A1(n11642), .A2(n11641), .A3(n11640), .A4(n11639), .ZN(N15349) );
  AOI22D1BWP30P140LVT U16376 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[1891]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1827]), .ZN(n11646) );
  AOI22D1BWP30P140LVT U16377 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1955]), .B1(n11757), .B2(
        inner_first_stage_data_reg[1923]), .ZN(n11645) );
  AOI22D1BWP30P140LVT U16378 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1795]), .B1(n11760), .B2(
        inner_first_stage_data_reg[1859]), .ZN(n11644) );
  AOI22D1BWP30P140LVT U16379 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[1987]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2019]), .ZN(n11643) );
  ND4D1BWP30P140LVT U16380 ( .A1(n11646), .A2(n11645), .A3(n11644), .A4(n11643), .ZN(N15350) );
  AOI22D1BWP30P140LVT U16381 ( .A1(n11757), .A2(
        inner_first_stage_data_reg[1924]), .B1(n11755), .B2(
        inner_first_stage_data_reg[1892]), .ZN(n11650) );
  AOI22D1BWP30P140LVT U16382 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1956]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1828]), .ZN(n11649) );
  AOI22D1BWP30P140LVT U16383 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1796]), .B1(n11760), .B2(
        inner_first_stage_data_reg[1860]), .ZN(n11648) );
  AOI22D1BWP30P140LVT U16384 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[1988]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2020]), .ZN(n11647) );
  ND4D1BWP30P140LVT U16385 ( .A1(n11650), .A2(n11649), .A3(n11648), .A4(n11647), .ZN(N15351) );
  AOI22D1BWP30P140LVT U16386 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1957]), .B1(n11755), .B2(
        inner_first_stage_data_reg[1893]), .ZN(n11654) );
  AOI22D1BWP30P140LVT U16387 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1797]), .B1(n11757), .B2(
        inner_first_stage_data_reg[1925]), .ZN(n11653) );
  AOI22D1BWP30P140LVT U16388 ( .A1(n11760), .A2(
        inner_first_stage_data_reg[1861]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1829]), .ZN(n11652) );
  AOI22D1BWP30P140LVT U16389 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[1989]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2021]), .ZN(n11651) );
  ND4D1BWP30P140LVT U16390 ( .A1(n11654), .A2(n11653), .A3(n11652), .A4(n11651), .ZN(N15352) );
  AOI22D1BWP30P140LVT U16391 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1958]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1830]), .ZN(n11658) );
  AOI22D1BWP30P140LVT U16392 ( .A1(n11757), .A2(
        inner_first_stage_data_reg[1926]), .B1(n11755), .B2(
        inner_first_stage_data_reg[1894]), .ZN(n11657) );
  AOI22D1BWP30P140LVT U16393 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1798]), .B1(n11760), .B2(
        inner_first_stage_data_reg[1862]), .ZN(n11656) );
  AOI22D1BWP30P140LVT U16394 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[1990]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2022]), .ZN(n11655) );
  ND4D1BWP30P140LVT U16395 ( .A1(n11658), .A2(n11657), .A3(n11656), .A4(n11655), .ZN(N15353) );
  AOI22D1BWP30P140LVT U16396 ( .A1(n11760), .A2(
        inner_first_stage_data_reg[1863]), .B1(n11757), .B2(
        inner_first_stage_data_reg[1927]), .ZN(n11662) );
  AOI22D1BWP30P140LVT U16397 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1799]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1831]), .ZN(n11661) );
  AOI22D1BWP30P140LVT U16398 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1959]), .B1(n11755), .B2(
        inner_first_stage_data_reg[1895]), .ZN(n11660) );
  AOI22D1BWP30P140LVT U16399 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[1991]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2023]), .ZN(n11659) );
  ND4D1BWP30P140LVT U16400 ( .A1(n11662), .A2(n11661), .A3(n11660), .A4(n11659), .ZN(N15354) );
  AOI22D1BWP30P140LVT U16401 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[1896]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1832]), .ZN(n11666) );
  AOI22D1BWP30P140LVT U16402 ( .A1(n11760), .A2(
        inner_first_stage_data_reg[1864]), .B1(n11757), .B2(
        inner_first_stage_data_reg[1928]), .ZN(n11665) );
  AOI22D1BWP30P140LVT U16403 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1960]), .B1(n11758), .B2(
        inner_first_stage_data_reg[1800]), .ZN(n11664) );
  AOI22D1BWP30P140LVT U16404 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[1992]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2024]), .ZN(n11663) );
  ND4D1BWP30P140LVT U16405 ( .A1(n11666), .A2(n11665), .A3(n11664), .A4(n11663), .ZN(N15355) );
  AOI22D1BWP30P140LVT U16406 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1801]), .B1(n11757), .B2(
        inner_first_stage_data_reg[1929]), .ZN(n11670) );
  AOI22D1BWP30P140LVT U16407 ( .A1(n11760), .A2(
        inner_first_stage_data_reg[1865]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1833]), .ZN(n11669) );
  AOI22D1BWP30P140LVT U16408 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1961]), .B1(n11755), .B2(
        inner_first_stage_data_reg[1897]), .ZN(n11668) );
  AOI22D1BWP30P140LVT U16409 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[1993]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2025]), .ZN(n11667) );
  ND4D1BWP30P140LVT U16410 ( .A1(n11670), .A2(n11669), .A3(n11668), .A4(n11667), .ZN(N15356) );
  AOI22D1BWP30P140LVT U16411 ( .A1(n11757), .A2(
        inner_first_stage_data_reg[1930]), .B1(n11755), .B2(
        inner_first_stage_data_reg[1898]), .ZN(n11674) );
  AOI22D1BWP30P140LVT U16412 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1962]), .B1(n11760), .B2(
        inner_first_stage_data_reg[1866]), .ZN(n11673) );
  AOI22D1BWP30P140LVT U16413 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1802]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1834]), .ZN(n11672) );
  AOI22D1BWP30P140LVT U16414 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[1994]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2026]), .ZN(n11671) );
  ND4D1BWP30P140LVT U16415 ( .A1(n11674), .A2(n11673), .A3(n11672), .A4(n11671), .ZN(N15357) );
  AOI22D1BWP30P140LVT U16416 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1803]), .B1(n11755), .B2(
        inner_first_stage_data_reg[1899]), .ZN(n11678) );
  AOI22D1BWP30P140LVT U16417 ( .A1(n11760), .A2(
        inner_first_stage_data_reg[1867]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1835]), .ZN(n11677) );
  AOI22D1BWP30P140LVT U16418 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1963]), .B1(n11757), .B2(
        inner_first_stage_data_reg[1931]), .ZN(n11676) );
  AOI22D1BWP30P140LVT U16419 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[1995]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2027]), .ZN(n11675) );
  ND4D1BWP30P140LVT U16420 ( .A1(n11678), .A2(n11677), .A3(n11676), .A4(n11675), .ZN(N15358) );
  AOI22D1BWP30P140LVT U16421 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1964]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1836]), .ZN(n11682) );
  AOI22D1BWP30P140LVT U16422 ( .A1(n11760), .A2(
        inner_first_stage_data_reg[1868]), .B1(n11757), .B2(
        inner_first_stage_data_reg[1932]), .ZN(n11681) );
  AOI22D1BWP30P140LVT U16423 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1804]), .B1(n11755), .B2(
        inner_first_stage_data_reg[1900]), .ZN(n11680) );
  AOI22D1BWP30P140LVT U16424 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[1996]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2028]), .ZN(n11679) );
  ND4D1BWP30P140LVT U16425 ( .A1(n11682), .A2(n11681), .A3(n11680), .A4(n11679), .ZN(N15359) );
  AOI22D1BWP30P140LVT U16426 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1805]), .B1(n11760), .B2(
        inner_first_stage_data_reg[1869]), .ZN(n11686) );
  AOI22D1BWP30P140LVT U16427 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[1901]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1837]), .ZN(n11685) );
  AOI22D1BWP30P140LVT U16428 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1965]), .B1(n11757), .B2(
        inner_first_stage_data_reg[1933]), .ZN(n11684) );
  AOI22D1BWP30P140LVT U16429 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[1997]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2029]), .ZN(n11683) );
  ND4D1BWP30P140LVT U16430 ( .A1(n11686), .A2(n11685), .A3(n11684), .A4(n11683), .ZN(N15360) );
  AOI22D1BWP30P140LVT U16431 ( .A1(n11760), .A2(
        inner_first_stage_data_reg[1870]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1838]), .ZN(n11690) );
  AOI22D1BWP30P140LVT U16432 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1966]), .B1(n11757), .B2(
        inner_first_stage_data_reg[1934]), .ZN(n11689) );
  AOI22D1BWP30P140LVT U16433 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1806]), .B1(n11755), .B2(
        inner_first_stage_data_reg[1902]), .ZN(n11688) );
  AOI22D1BWP30P140LVT U16434 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[1998]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2030]), .ZN(n11687) );
  ND4D1BWP30P140LVT U16435 ( .A1(n11690), .A2(n11689), .A3(n11688), .A4(n11687), .ZN(N15361) );
  AOI22D1BWP30P140LVT U16436 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1807]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1839]), .ZN(n11694) );
  AOI22D1BWP30P140LVT U16437 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1967]), .B1(n11760), .B2(
        inner_first_stage_data_reg[1871]), .ZN(n11693) );
  AOI22D1BWP30P140LVT U16438 ( .A1(n11757), .A2(
        inner_first_stage_data_reg[1935]), .B1(n11755), .B2(
        inner_first_stage_data_reg[1903]), .ZN(n11692) );
  AOI22D1BWP30P140LVT U16439 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[1999]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2031]), .ZN(n11691) );
  ND4D1BWP30P140LVT U16440 ( .A1(n11694), .A2(n11693), .A3(n11692), .A4(n11691), .ZN(N15362) );
  AOI22D1BWP30P140LVT U16441 ( .A1(n11760), .A2(
        inner_first_stage_data_reg[1872]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1840]), .ZN(n11698) );
  AOI22D1BWP30P140LVT U16442 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1968]), .B1(n11755), .B2(
        inner_first_stage_data_reg[1904]), .ZN(n11697) );
  AOI22D1BWP30P140LVT U16443 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1808]), .B1(n11757), .B2(
        inner_first_stage_data_reg[1936]), .ZN(n11696) );
  AOI22D1BWP30P140LVT U16444 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[2000]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2032]), .ZN(n11695) );
  ND4D1BWP30P140LVT U16445 ( .A1(n11698), .A2(n11697), .A3(n11696), .A4(n11695), .ZN(N15363) );
  AOI22D1BWP30P140LVT U16446 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[1905]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1841]), .ZN(n11702) );
  AOI22D1BWP30P140LVT U16447 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1809]), .B1(n11760), .B2(
        inner_first_stage_data_reg[1873]), .ZN(n11701) );
  AOI22D1BWP30P140LVT U16448 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1969]), .B1(n11757), .B2(
        inner_first_stage_data_reg[1937]), .ZN(n11700) );
  AOI22D1BWP30P140LVT U16449 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[2001]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2033]), .ZN(n11699) );
  ND4D1BWP30P140LVT U16450 ( .A1(n11702), .A2(n11701), .A3(n11700), .A4(n11699), .ZN(N15364) );
  AOI22D1BWP30P140LVT U16451 ( .A1(n11757), .A2(
        inner_first_stage_data_reg[1938]), .B1(n11755), .B2(
        inner_first_stage_data_reg[1906]), .ZN(n11706) );
  AOI22D1BWP30P140LVT U16452 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1810]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1842]), .ZN(n11705) );
  AOI22D1BWP30P140LVT U16453 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1970]), .B1(n11760), .B2(
        inner_first_stage_data_reg[1874]), .ZN(n11704) );
  AOI22D1BWP30P140LVT U16454 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[2002]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2034]), .ZN(n11703) );
  ND4D1BWP30P140LVT U16455 ( .A1(n11706), .A2(n11705), .A3(n11704), .A4(n11703), .ZN(N15365) );
  AOI22D1BWP30P140LVT U16456 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1971]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1843]), .ZN(n11710) );
  AOI22D1BWP30P140LVT U16457 ( .A1(n11760), .A2(
        inner_first_stage_data_reg[1875]), .B1(n11757), .B2(
        inner_first_stage_data_reg[1939]), .ZN(n11709) );
  AOI22D1BWP30P140LVT U16458 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1811]), .B1(n11755), .B2(
        inner_first_stage_data_reg[1907]), .ZN(n11708) );
  AOI22D1BWP30P140LVT U16459 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[2003]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2035]), .ZN(n11707) );
  ND4D1BWP30P140LVT U16460 ( .A1(n11710), .A2(n11709), .A3(n11708), .A4(n11707), .ZN(N15366) );
  AOI22D1BWP30P140LVT U16461 ( .A1(n11760), .A2(
        inner_first_stage_data_reg[1876]), .B1(n11757), .B2(
        inner_first_stage_data_reg[1940]), .ZN(n11714) );
  AOI22D1BWP30P140LVT U16462 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1812]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1844]), .ZN(n11713) );
  AOI22D1BWP30P140LVT U16463 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1972]), .B1(n11755), .B2(
        inner_first_stage_data_reg[1908]), .ZN(n11712) );
  AOI22D1BWP30P140LVT U16464 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[2004]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2036]), .ZN(n11711) );
  ND4D1BWP30P140LVT U16465 ( .A1(n11714), .A2(n11713), .A3(n11712), .A4(n11711), .ZN(N15367) );
  AOI22D1BWP30P140LVT U16466 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1813]), .B1(n11757), .B2(
        inner_first_stage_data_reg[1941]), .ZN(n11718) );
  AOI22D1BWP30P140LVT U16467 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1973]), .B1(n11760), .B2(
        inner_first_stage_data_reg[1877]), .ZN(n11717) );
  AOI22D1BWP30P140LVT U16468 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[1909]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1845]), .ZN(n11716) );
  AOI22D1BWP30P140LVT U16469 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[2005]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2037]), .ZN(n11715) );
  ND4D1BWP30P140LVT U16470 ( .A1(n11718), .A2(n11717), .A3(n11716), .A4(n11715), .ZN(N15368) );
  AOI22D1BWP30P140LVT U16471 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1814]), .B1(n11757), .B2(
        inner_first_stage_data_reg[1942]), .ZN(n11722) );
  AOI22D1BWP30P140LVT U16472 ( .A1(n11760), .A2(
        inner_first_stage_data_reg[1878]), .B1(n11755), .B2(
        inner_first_stage_data_reg[1910]), .ZN(n11721) );
  AOI22D1BWP30P140LVT U16473 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1974]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1846]), .ZN(n11720) );
  AOI22D1BWP30P140LVT U16474 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[2006]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2038]), .ZN(n11719) );
  ND4D1BWP30P140LVT U16475 ( .A1(n11722), .A2(n11721), .A3(n11720), .A4(n11719), .ZN(N15369) );
  AOI22D1BWP30P140LVT U16476 ( .A1(n11757), .A2(
        inner_first_stage_data_reg[1943]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1847]), .ZN(n11726) );
  AOI22D1BWP30P140LVT U16477 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1975]), .B1(n11758), .B2(
        inner_first_stage_data_reg[1815]), .ZN(n11725) );
  AOI22D1BWP30P140LVT U16478 ( .A1(n11760), .A2(
        inner_first_stage_data_reg[1879]), .B1(n11755), .B2(
        inner_first_stage_data_reg[1911]), .ZN(n11724) );
  AOI22D1BWP30P140LVT U16479 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[2007]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2039]), .ZN(n11723) );
  ND4D1BWP30P140LVT U16480 ( .A1(n11726), .A2(n11725), .A3(n11724), .A4(n11723), .ZN(N15370) );
  AOI22D1BWP30P140LVT U16481 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[1912]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1848]), .ZN(n11730) );
  AOI22D1BWP30P140LVT U16482 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1816]), .B1(n11760), .B2(
        inner_first_stage_data_reg[1880]), .ZN(n11729) );
  AOI22D1BWP30P140LVT U16483 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1976]), .B1(n11757), .B2(
        inner_first_stage_data_reg[1944]), .ZN(n11728) );
  AOI22D1BWP30P140LVT U16484 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[2008]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2040]), .ZN(n11727) );
  ND4D1BWP30P140LVT U16485 ( .A1(n11730), .A2(n11729), .A3(n11728), .A4(n11727), .ZN(N15371) );
  AOI22D1BWP30P140LVT U16486 ( .A1(n11760), .A2(
        inner_first_stage_data_reg[1881]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1849]), .ZN(n11734) );
  AOI22D1BWP30P140LVT U16487 ( .A1(n11757), .A2(
        inner_first_stage_data_reg[1945]), .B1(n11755), .B2(
        inner_first_stage_data_reg[1913]), .ZN(n11733) );
  AOI22D1BWP30P140LVT U16488 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1977]), .B1(n11758), .B2(
        inner_first_stage_data_reg[1817]), .ZN(n11732) );
  AOI22D1BWP30P140LVT U16489 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[2009]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2041]), .ZN(n11731) );
  ND4D1BWP30P140LVT U16490 ( .A1(n11734), .A2(n11733), .A3(n11732), .A4(n11731), .ZN(N15372) );
  AOI22D1BWP30P140LVT U16491 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1818]), .B1(n11757), .B2(
        inner_first_stage_data_reg[1946]), .ZN(n11738) );
  AOI22D1BWP30P140LVT U16492 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1978]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1850]), .ZN(n11737) );
  AOI22D1BWP30P140LVT U16493 ( .A1(n11760), .A2(
        inner_first_stage_data_reg[1882]), .B1(n11755), .B2(
        inner_first_stage_data_reg[1914]), .ZN(n11736) );
  AOI22D1BWP30P140LVT U16494 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[2010]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2042]), .ZN(n11735) );
  ND4D1BWP30P140LVT U16495 ( .A1(n11738), .A2(n11737), .A3(n11736), .A4(n11735), .ZN(N15373) );
  AOI22D1BWP30P140LVT U16496 ( .A1(n11760), .A2(
        inner_first_stage_data_reg[1883]), .B1(n11755), .B2(
        inner_first_stage_data_reg[1915]), .ZN(n11742) );
  AOI22D1BWP30P140LVT U16497 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1979]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1851]), .ZN(n11741) );
  AOI22D1BWP30P140LVT U16498 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1819]), .B1(n11757), .B2(
        inner_first_stage_data_reg[1947]), .ZN(n11740) );
  AOI22D1BWP30P140LVT U16499 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[2011]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2043]), .ZN(n11739) );
  ND4D1BWP30P140LVT U16500 ( .A1(n11742), .A2(n11741), .A3(n11740), .A4(n11739), .ZN(N15374) );
  AOI22D1BWP30P140LVT U16501 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1980]), .B1(n11758), .B2(
        inner_first_stage_data_reg[1820]), .ZN(n11746) );
  AOI22D1BWP30P140LVT U16502 ( .A1(n11757), .A2(
        inner_first_stage_data_reg[1948]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1852]), .ZN(n11745) );
  AOI22D1BWP30P140LVT U16503 ( .A1(n11760), .A2(
        inner_first_stage_data_reg[1884]), .B1(n11755), .B2(
        inner_first_stage_data_reg[1916]), .ZN(n11744) );
  AOI22D1BWP30P140LVT U16504 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[2012]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2044]), .ZN(n11743) );
  ND4D1BWP30P140LVT U16505 ( .A1(n11746), .A2(n11745), .A3(n11744), .A4(n11743), .ZN(N15375) );
  AOI22D1BWP30P140LVT U16506 ( .A1(n11757), .A2(
        inner_first_stage_data_reg[1949]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1853]), .ZN(n11750) );
  AOI22D1BWP30P140LVT U16507 ( .A1(n11760), .A2(
        inner_first_stage_data_reg[1885]), .B1(n11755), .B2(
        inner_first_stage_data_reg[1917]), .ZN(n11749) );
  AOI22D1BWP30P140LVT U16508 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1981]), .B1(n11758), .B2(
        inner_first_stage_data_reg[1821]), .ZN(n11748) );
  AOI22D1BWP30P140LVT U16509 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[2013]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2045]), .ZN(n11747) );
  ND4D1BWP30P140LVT U16510 ( .A1(n11750), .A2(n11749), .A3(n11748), .A4(n11747), .ZN(N15376) );
  AOI22D1BWP30P140LVT U16511 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1982]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1854]), .ZN(n11754) );
  AOI22D1BWP30P140LVT U16512 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1822]), .B1(n11755), .B2(
        inner_first_stage_data_reg[1918]), .ZN(n11753) );
  AOI22D1BWP30P140LVT U16513 ( .A1(n11760), .A2(
        inner_first_stage_data_reg[1886]), .B1(n11757), .B2(
        inner_first_stage_data_reg[1950]), .ZN(n11752) );
  AOI22D1BWP30P140LVT U16514 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[2014]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2046]), .ZN(n11751) );
  ND4D1BWP30P140LVT U16515 ( .A1(n11754), .A2(n11753), .A3(n11752), .A4(n11751), .ZN(N15377) );
  AOI22D1BWP30P140LVT U16516 ( .A1(n11756), .A2(
        inner_first_stage_data_reg[1983]), .B1(n11755), .B2(
        inner_first_stage_data_reg[1919]), .ZN(n11766) );
  AOI22D1BWP30P140LVT U16517 ( .A1(n11758), .A2(
        inner_first_stage_data_reg[1823]), .B1(n11757), .B2(
        inner_first_stage_data_reg[1951]), .ZN(n11765) );
  AOI22D1BWP30P140LVT U16518 ( .A1(n11760), .A2(
        inner_first_stage_data_reg[1887]), .B1(n11759), .B2(
        inner_first_stage_data_reg[1855]), .ZN(n11764) );
  AOI22D1BWP30P140LVT U16519 ( .A1(n11762), .A2(
        inner_first_stage_data_reg[2015]), .B1(n11761), .B2(
        inner_first_stage_data_reg[2047]), .ZN(n11763) );
  ND4D1BWP30P140LVT U16520 ( .A1(n11766), .A2(n11765), .A3(n11764), .A4(n11763), .ZN(N15378) );
endmodule

