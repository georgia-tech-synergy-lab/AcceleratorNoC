`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////////////////////
// Company: Gatech	
// Engineer: Mandovi Mukherjee
// 
// Create Date: 01/08/2021 
// System Name: accelerator
// Module Name: local controller
// Project Name: ARION DRBE
// Description: fetch and push data out to network; assuming the output from
// global controller comes in the form of a packet
// Dependencies:
// Additional Comments: 
/////////////////////////////////////////////////////////////////////////////////////////////////////

module global_controller(CLK, reset, boot_up, delay_matrix_N_1, from_glob_controller_delay,   from_glob_dest_addr,  from_glob_controller_valid,   write_flag, from_glob_prefetch_valid, from_glob_prefetch_start, from_glob_prefetch_stop, from_glob_prefetch_dest,  scenario_update);

    // parameter
    	parameter N_sample = 256;
	parameter datawidth = 16;
	parameter address_vector_width = 8; //can be 200 or 8: 8 for small tapeout
	parameter id_width = 4; // 16 local controllers in subscaled system
	parameter sample_address_width = 8; /// assuming 256 words: needs to change if arrangement is different
	parameter packet_width = 2*datawidth + address_vector_width;
	parameter delay_length = 12; // log(id_width*N_sample)
	

//=== IO Ports ===//


    // input
    	input CLK; // system clock, generated by VCO
	input reset;
	input boot_up;
	input [delay_length - 1:0] delay_matrx_N_1[address_vector_width - 1:0]



    // output
	output reg from_glob_controller_valid;
	output reg [address_vector_width - 1:0] from_glob_dest_addr;
	output reg [address_vector_width - 1:0] from_glob_prefetch_dest;
	output reg [sample_address_width - 1:0] from_glob_controller_delay;
	
        
	output reg write_flag;

	output reg from_glob_prefetch_valid;
	output reg [sample_address_width - 1:0] from_glob_prefetch_start;
	output reg [sample_address_width - 1:0] from_glob_prefetch_stop;
	input scenario_update;



//////////// internal status regs/signals //////////////////////////////////



///////////////////////////////////////////////////////////////////////////////    

////////// logic part ///////////////////////////////////////////////////////  




////////////sequential logic
//
//

	always @(posedge CLK) begin
	
		if (reset) begin
			from_glob_controller_delay <= 0;
			from_glob_controller_valid <= 0;
			from_glob_dest_addr <= 0;
			from_glob_prefetch_dest <= 0;
	 		from_glob_prefetch_start <= 0;
	 		from_glob_prefetch_stop <= 0;
			from_glob_prefetch_valid <= 0;
			scenario_update <= 0;
		end
		else if (boot_up) begin
			from_glob_controller_delay <= 0;
			from_glob_controller_valid <= 0;
			from_glob_dest_addr <= 0;
			from_glob_prefetch_dest <= 0;
	 		from_glob_prefetch_start <= 0;
	 		from_glob_prefetch_stop <= 0;
			from_glob_prefetch_valid <= 0;
			scenario_update <= 0;
		end
		else begin
			if (~scenario_update) begin
		
			end
			else begin
				if (busy) begin
					from_glob_prefetch_dest <= from_glob_prefetch_dest;
					from_glob_prefetch_start <= from_glob_prefetch_start;
					from_glob_prefetch_stop <= from_glob_prefetch_stop;
					from_glob_prefetch_valid <= 0;
					scenario_update <= scenario_update;
				end
				else begin
					from_glob_prefetch_dest <= calc_glob_prefetch_dest;
					from_glob_prefetch_start <= calc_glob_prefetch_start;
					from_glob_prefetch_stop <= calc_glob_prefetch_stop;
					from_glob_prefetch_valid <= 1;
					scenario_update <= scenario_update;

				end
			end
			

		end

	end
	 
	 


   
endmodule
    
