`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////////////////////
// Company: Gatech	
// Engineer: Mandovi Mukherjee
// 
// Create Date: 01/08/2021 
// System Name: accelerator
// Module Name: local controller
// Project Name: ARION DRBE
// Description: fetch and push data out to network; assuming the output from
// global controller comes in the form of a packet
// Dependencies:
// Additional Comments: 
/////////////////////////////////////////////////////////////////////////////////////////////////////

module local_controller_simple_trial(clk, reset, init, controller_id, write_flag, glob_controller_sending, from_glob_controller_delay, data_from_sram, input_boundary_flag, prev_dest_address, from_glob_dest_addr, packet_out, boundary_next, dest_address, scenario_end_flag, );
    // parameter
    parameter N_row = 1024;
	parameter datawidth = 32;
	parameter address_vector_width = 8; //can be 200 or 8: 8 for subscaled system
	parameter id_width = 11; // 1221 local controllers in subscaled system
	parameter row_address_width = 10; /// assuming 1024 rows and 64 columns: needs to change if arrangement is different
	parameter packet_width = 2*datawidth + address_vector_width;
	
	
	
        
    // input
    input clk; // system clock, generated by VCO
	input reset;
	input init;
	input glob_controller_sending; //not used
	input [2*datawidth - 1:0] data_from_sram;
	//input [2*datawidth - 1:0] prefetch_data_from_sram;
	input [id_width - 1:0] controller_id;
	input input_boundary_flag;
	input write_flag;
	input [address_vector_width - 1:0] prev_dest_address;
	input [address_vector_width - 1:0] from_glob_dest_addr;
	input [row_address_width - 1:0] from_glob_controller_delay;
	input scenario_end_flag;

    // output
    output [packet_width-1:0] packet_out; 
    //output [packet_width-1:0] prefetch_packet_out; 
    output reg boundary_next;
    output reg [address_vector_width - 1:0] dest_address;
	
	

    // internal status regs/signals
    reg [row_address_width-1:0] row_address;
	reg [id_width - 1:0] id; 
	reg [packet_width-1:0] packet_out_internal;
	//reg [packet_width-1:0] prefetch_packet_out_internal;
	reg coeff_num;
	reg [row_address_width - 1:0] delay;
    

    // logic part  
    assign packet_out = packet_out_internal;
    //assign prefetch_packet_out = prefetch_packet_out_internal;

	//sequential logic
    always @ (posedge clk) begin
        if (reset) begin
			id <= 0;
			row_address <= 0;
			//prefetch_row_address <= 0;
			packet_out_internal <= 264'bz;
			//prefetch_packet_out_internal <= 264'bz;
			dest_address <= 0;
			coeff_num <= 0;
			delay <= 0;
			//prefetch_reqd <= 0;
			//prefetch_dest_address <= 0;
			
        end
        else if (init) begin
			id <= controller_id;
			packet_out_internal <= 264'bz;
			//prefetch_packet_out_internal <= 264'bz;
			
			if (from_glob_dest_addr[0] == 1'b1 || from_glob_dest_addr[0] == 1'b0) begin
				row_address <= from_glob_controller_delay;
				//prefetch_row_address <= prefetch_row_address;
				dest_address <= from_glob_dest_addr;
				coeff_num <= 1;
				delay <= from_glob_controller_delay;
				//prefetch_reqd <= prefetch_reqd;
			end

			if (from_glob_dest_addr[0] == 1'b1 || from_glob_dest_addr[0] == 1'b0) begin
				row_address <= from_glob_controller_delay;
				//prefetch_row_address <= prefetch_row_address;
				dest_address <= from_glob_dest_addr;
				coeff_num <= 1;
				delay <= from_glob_controller_delay;
				//prefetch_reqd <= prefetch_reqd;
			end

			
			else begin
				row_address <= row_address;
				//prefetch_row_address <= prefetch_row_address;
				dest_address <= dest_address;
				coeff_num <= coeff_num;
				delay <= delay;
				//prefetch_reqd <= prefetch_reqd;
			end
			
        end
		else begin
			if (coeff_num == 1 && write_flag == 0) begin
				packet_out_internal <= {data_from_sram, dest_address};
				row_address <= row_address + 1;
				//prefetch_packet_out_internal <= 264'bz;
				//prefetch_row_address <= prefetch_row_address;
			end
			else if (coeff_num == 1 && write_flag == 1) begin
				packet_out_internal <= {64'b0, dest_address};
				row_address <= row_address + 1;	
				//prefetch_packet_out_internal <= 264'bz;
				//prefetch_row_address <= prefetch_row_address;

			end

			id <= id;
			dest_address <= dest_address;
			coeff_num <= coeff_num;
			delay <= delay;
		end  
     end
	 
	 always @ (posedge clk) begin
		if (row_address == N_row - 1) begin
			boundary_next <= 1;
		end
		else begin
			boundary_next <= 0;
		end
	 end
	 
	 
	 


   
endmodule
    
