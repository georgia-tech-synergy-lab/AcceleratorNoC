module mux_tree_128_1_seq #(
	parameter DATA_WIDTH = 32,      // could be arbitrary number
	parameter NUM_OUTPUT_DATA  = 1, // must be power of 2.
	parameter NUM_INPUT_DATA = 128   
)(
    // timeing signals
    CLK,
	rst,
	
    // data signals
	i_valid,        // valid input data signal
	i_data_bus,     // input data bus coming into distribute switch
	
	o_valid,        // output valid
    o_data_bus,     // output data 

	// control signals
	i_en,           // distribute switch enable
	i_cmd           // the input should be one-hot encoded command 
);
	//parameter
	localparam TOTAL_COMMAND = NUM_INPUT_DATA*NUM_OUTPUT_DATA;
	
	localparam WIDTH_INPUT_DATA = NUM_INPUT_DATA*DATA_WIDTH;
	localparam WIDTH_OUTPUT_DATA = NUM_OUTPUT_DATA*DATA_WIDTH;
	
    // interface
	input                                        CLK;
	input                                        rst;

	input  [NUM_INPUT_DATA-1:0]                  i_valid;             
	input  [WIDTH_INPUT_DATA-1:0]                i_data_bus;

	output [NUM_OUTPUT_DATA-1:0]                 o_valid;             
	output [WIDTH_OUTPUT_DATA-1:0]               o_data_bus; // {o_data_a, o_data_b}

	input                                        i_en;
	input  [TOTAL_COMMAND-1:0]                   i_cmd;

    reg    [NUM_OUTPUT_DATA-1:0]                 o_valid_reg;
    reg    [WIDTH_OUTPUT_DATA-1:0]               o_data_bus_reg;

    genvar i,j;
    generate
        for(i=0; i<NUM_OUTPUT_DATA; i=i+1)
        begin: o_data_output_mux
            
            // data mux
            wire [NUM_INPUT_DATA-1:0] inner_cmd_wire;
            assign inner_cmd_wire = {i_cmd[127*NUM_OUTPUT_DATA+i],i_cmd[126*NUM_OUTPUT_DATA+i],i_cmd[125*NUM_OUTPUT_DATA+i],i_cmd[124*NUM_OUTPUT_DATA+i],i_cmd[123*NUM_OUTPUT_DATA+i],i_cmd[122*NUM_OUTPUT_DATA+i],i_cmd[121*NUM_OUTPUT_DATA+i],i_cmd[120*NUM_OUTPUT_DATA+i],i_cmd[119*NUM_OUTPUT_DATA+i],i_cmd[118*NUM_OUTPUT_DATA+i],i_cmd[117*NUM_OUTPUT_DATA+i],i_cmd[116*NUM_OUTPUT_DATA+i],i_cmd[115*NUM_OUTPUT_DATA+i],i_cmd[114*NUM_OUTPUT_DATA+i],i_cmd[113*NUM_OUTPUT_DATA+i],i_cmd[112*NUM_OUTPUT_DATA+i],i_cmd[111*NUM_OUTPUT_DATA+i],i_cmd[110*NUM_OUTPUT_DATA+i],i_cmd[109*NUM_OUTPUT_DATA+i],i_cmd[108*NUM_OUTPUT_DATA+i],i_cmd[107*NUM_OUTPUT_DATA+i],i_cmd[106*NUM_OUTPUT_DATA+i],i_cmd[105*NUM_OUTPUT_DATA+i],i_cmd[104*NUM_OUTPUT_DATA+i],i_cmd[103*NUM_OUTPUT_DATA+i],i_cmd[102*NUM_OUTPUT_DATA+i],i_cmd[101*NUM_OUTPUT_DATA+i],i_cmd[100*NUM_OUTPUT_DATA+i],i_cmd[99*NUM_OUTPUT_DATA+i],i_cmd[98*NUM_OUTPUT_DATA+i],i_cmd[97*NUM_OUTPUT_DATA+i],i_cmd[96*NUM_OUTPUT_DATA+i],i_cmd[95*NUM_OUTPUT_DATA+i],i_cmd[94*NUM_OUTPUT_DATA+i],i_cmd[93*NUM_OUTPUT_DATA+i],i_cmd[92*NUM_OUTPUT_DATA+i],i_cmd[91*NUM_OUTPUT_DATA+i],i_cmd[90*NUM_OUTPUT_DATA+i],i_cmd[89*NUM_OUTPUT_DATA+i],i_cmd[88*NUM_OUTPUT_DATA+i],i_cmd[87*NUM_OUTPUT_DATA+i],i_cmd[86*NUM_OUTPUT_DATA+i],i_cmd[85*NUM_OUTPUT_DATA+i],i_cmd[84*NUM_OUTPUT_DATA+i],i_cmd[83*NUM_OUTPUT_DATA+i],i_cmd[82*NUM_OUTPUT_DATA+i],i_cmd[81*NUM_OUTPUT_DATA+i],i_cmd[80*NUM_OUTPUT_DATA+i],i_cmd[79*NUM_OUTPUT_DATA+i],i_cmd[78*NUM_OUTPUT_DATA+i],i_cmd[77*NUM_OUTPUT_DATA+i],i_cmd[76*NUM_OUTPUT_DATA+i],i_cmd[75*NUM_OUTPUT_DATA+i],i_cmd[74*NUM_OUTPUT_DATA+i],i_cmd[73*NUM_OUTPUT_DATA+i],i_cmd[72*NUM_OUTPUT_DATA+i],i_cmd[71*NUM_OUTPUT_DATA+i],i_cmd[70*NUM_OUTPUT_DATA+i],i_cmd[69*NUM_OUTPUT_DATA+i],i_cmd[68*NUM_OUTPUT_DATA+i],i_cmd[67*NUM_OUTPUT_DATA+i],i_cmd[66*NUM_OUTPUT_DATA+i],i_cmd[65*NUM_OUTPUT_DATA+i],i_cmd[64*NUM_OUTPUT_DATA+i],i_cmd[63*NUM_OUTPUT_DATA+i],i_cmd[62*NUM_OUTPUT_DATA+i],i_cmd[61*NUM_OUTPUT_DATA+i],i_cmd[60*NUM_OUTPUT_DATA+i],i_cmd[59*NUM_OUTPUT_DATA+i],i_cmd[58*NUM_OUTPUT_DATA+i],i_cmd[57*NUM_OUTPUT_DATA+i],i_cmd[56*NUM_OUTPUT_DATA+i],i_cmd[55*NUM_OUTPUT_DATA+i],i_cmd[54*NUM_OUTPUT_DATA+i],i_cmd[53*NUM_OUTPUT_DATA+i],i_cmd[52*NUM_OUTPUT_DATA+i],i_cmd[51*NUM_OUTPUT_DATA+i],i_cmd[50*NUM_OUTPUT_DATA+i],i_cmd[49*NUM_OUTPUT_DATA+i],i_cmd[48*NUM_OUTPUT_DATA+i],i_cmd[47*NUM_OUTPUT_DATA+i],i_cmd[46*NUM_OUTPUT_DATA+i],i_cmd[45*NUM_OUTPUT_DATA+i],i_cmd[44*NUM_OUTPUT_DATA+i],i_cmd[43*NUM_OUTPUT_DATA+i],i_cmd[42*NUM_OUTPUT_DATA+i],i_cmd[41*NUM_OUTPUT_DATA+i],i_cmd[40*NUM_OUTPUT_DATA+i],i_cmd[39*NUM_OUTPUT_DATA+i],i_cmd[38*NUM_OUTPUT_DATA+i],i_cmd[37*NUM_OUTPUT_DATA+i],i_cmd[36*NUM_OUTPUT_DATA+i],i_cmd[35*NUM_OUTPUT_DATA+i],i_cmd[34*NUM_OUTPUT_DATA+i],i_cmd[33*NUM_OUTPUT_DATA+i],i_cmd[32*NUM_OUTPUT_DATA+i],i_cmd[31*NUM_OUTPUT_DATA+i],i_cmd[30*NUM_OUTPUT_DATA+i],i_cmd[29*NUM_OUTPUT_DATA+i],i_cmd[28*NUM_OUTPUT_DATA+i],i_cmd[27*NUM_OUTPUT_DATA+i],i_cmd[26*NUM_OUTPUT_DATA+i],i_cmd[25*NUM_OUTPUT_DATA+i],i_cmd[24*NUM_OUTPUT_DATA+i],i_cmd[23*NUM_OUTPUT_DATA+i],i_cmd[22*NUM_OUTPUT_DATA+i],i_cmd[21*NUM_OUTPUT_DATA+i],i_cmd[20*NUM_OUTPUT_DATA+i],i_cmd[19*NUM_OUTPUT_DATA+i],i_cmd[18*NUM_OUTPUT_DATA+i],i_cmd[17*NUM_OUTPUT_DATA+i],i_cmd[16*NUM_OUTPUT_DATA+i],i_cmd[15*NUM_OUTPUT_DATA+i],i_cmd[14*NUM_OUTPUT_DATA+i],i_cmd[13*NUM_OUTPUT_DATA+i],i_cmd[12*NUM_OUTPUT_DATA+i],i_cmd[11*NUM_OUTPUT_DATA+i],i_cmd[10*NUM_OUTPUT_DATA+i],i_cmd[9*NUM_OUTPUT_DATA+i],i_cmd[8*NUM_OUTPUT_DATA+i],i_cmd[7*NUM_OUTPUT_DATA+i],i_cmd[6*NUM_OUTPUT_DATA+i],i_cmd[5*NUM_OUTPUT_DATA+i],i_cmd[4*NUM_OUTPUT_DATA+i],i_cmd[3*NUM_OUTPUT_DATA+i],i_cmd[2*NUM_OUTPUT_DATA+i],i_cmd[1*NUM_OUTPUT_DATA+i],i_cmd[0*NUM_OUTPUT_DATA+i]};
            always@(posedge CLK)
            begin
               if(i_en && (~rst))
                begin
                    case(inner_cmd_wire)
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[0])?i_data_bus[0*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[1])?i_data_bus[1*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[2])?i_data_bus[2*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[3])?i_data_bus[3*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[4])?i_data_bus[4*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[5])?i_data_bus[5*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[6])?i_data_bus[6*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[7])?i_data_bus[7*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[8])?i_data_bus[8*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[9])?i_data_bus[9*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[10])?i_data_bus[10*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[11])?i_data_bus[11*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[12])?i_data_bus[12*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[13])?i_data_bus[13*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[14])?i_data_bus[14*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[15])?i_data_bus[15*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[16])?i_data_bus[16*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[17])?i_data_bus[17*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[18])?i_data_bus[18*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[19])?i_data_bus[19*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[20])?i_data_bus[20*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[21])?i_data_bus[21*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[22])?i_data_bus[22*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[23])?i_data_bus[23*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[24])?i_data_bus[24*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[25])?i_data_bus[25*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[26])?i_data_bus[26*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[27])?i_data_bus[27*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[28])?i_data_bus[28*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[29])?i_data_bus[29*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[30])?i_data_bus[30*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[31])?i_data_bus[31*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[32])?i_data_bus[32*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[33])?i_data_bus[33*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[34])?i_data_bus[34*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[35])?i_data_bus[35*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[36])?i_data_bus[36*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[37])?i_data_bus[37*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[38])?i_data_bus[38*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[39])?i_data_bus[39*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[40])?i_data_bus[40*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[41])?i_data_bus[41*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[42])?i_data_bus[42*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[43])?i_data_bus[43*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[44])?i_data_bus[44*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[45])?i_data_bus[45*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[46])?i_data_bus[46*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[47])?i_data_bus[47*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[48])?i_data_bus[48*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[49])?i_data_bus[49*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[50])?i_data_bus[50*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[51])?i_data_bus[51*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[52])?i_data_bus[52*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[53])?i_data_bus[53*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[54])?i_data_bus[54*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[55])?i_data_bus[55*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[56])?i_data_bus[56*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[57])?i_data_bus[57*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[58])?i_data_bus[58*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[59])?i_data_bus[59*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[60])?i_data_bus[60*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[61])?i_data_bus[61*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[62])?i_data_bus[62*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[63])?i_data_bus[63*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[64])?i_data_bus[64*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[65])?i_data_bus[65*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[66])?i_data_bus[66*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[67])?i_data_bus[67*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[68])?i_data_bus[68*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[69])?i_data_bus[69*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[70])?i_data_bus[70*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[71])?i_data_bus[71*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[72])?i_data_bus[72*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[73])?i_data_bus[73*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[74])?i_data_bus[74*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[75])?i_data_bus[75*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[76])?i_data_bus[76*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[77])?i_data_bus[77*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[78])?i_data_bus[78*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[79])?i_data_bus[79*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[80])?i_data_bus[80*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[81])?i_data_bus[81*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[82])?i_data_bus[82*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[83])?i_data_bus[83*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[84])?i_data_bus[84*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[85])?i_data_bus[85*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[86])?i_data_bus[86*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[87])?i_data_bus[87*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[88])?i_data_bus[88*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[89])?i_data_bus[89*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[90])?i_data_bus[90*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[91])?i_data_bus[91*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[92])?i_data_bus[92*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[93])?i_data_bus[93*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[94])?i_data_bus[94*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[95])?i_data_bus[95*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[96])?i_data_bus[96*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[97])?i_data_bus[97*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[98])?i_data_bus[98*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[99])?i_data_bus[99*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[100])?i_data_bus[100*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[101])?i_data_bus[101*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[102])?i_data_bus[102*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[103])?i_data_bus[103*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[104])?i_data_bus[104*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[105])?i_data_bus[105*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[106])?i_data_bus[106*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[107])?i_data_bus[107*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[108])?i_data_bus[108*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[109])?i_data_bus[109*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[110])?i_data_bus[110*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[111])?i_data_bus[111*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[112])?i_data_bus[112*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[113])?i_data_bus[113*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[114])?i_data_bus[114*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[115])?i_data_bus[115*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[116])?i_data_bus[116*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[117])?i_data_bus[117*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[118])?i_data_bus[118*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[119])?i_data_bus[119*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[120])?i_data_bus[120*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[121])?i_data_bus[121*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[122])?i_data_bus[122*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[123])?i_data_bus[123*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[124])?i_data_bus[124*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[125])?i_data_bus[125*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[126])?i_data_bus[126*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        128'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= (i_valid[127])?i_data_bus[127*DATA_WIDTH+:DATA_WIDTH]:{DATA_WIDTH{1'b0}};
                        end
                        default:
                        begin
                            o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= {DATA_WIDTH{1'b0}};
                        end
                    endcase
                end
                else
                begin
                    o_data_bus_reg[i*DATA_WIDTH+:DATA_WIDTH] <= {WIDTH_OUTPUT_DATA{1'b0}};
                end
            end

            // valid mux
            wire [NUM_INPUT_DATA-1:0] inner_cmd_wire_valid;
            assign inner_cmd_wire_valid = {i_cmd[127*NUM_OUTPUT_DATA+i],i_cmd[126*NUM_OUTPUT_DATA+i],i_cmd[125*NUM_OUTPUT_DATA+i],i_cmd[124*NUM_OUTPUT_DATA+i],i_cmd[123*NUM_OUTPUT_DATA+i],i_cmd[122*NUM_OUTPUT_DATA+i],i_cmd[121*NUM_OUTPUT_DATA+i],i_cmd[120*NUM_OUTPUT_DATA+i],i_cmd[119*NUM_OUTPUT_DATA+i],i_cmd[118*NUM_OUTPUT_DATA+i],i_cmd[117*NUM_OUTPUT_DATA+i],i_cmd[116*NUM_OUTPUT_DATA+i],i_cmd[115*NUM_OUTPUT_DATA+i],i_cmd[114*NUM_OUTPUT_DATA+i],i_cmd[113*NUM_OUTPUT_DATA+i],i_cmd[112*NUM_OUTPUT_DATA+i],i_cmd[111*NUM_OUTPUT_DATA+i],i_cmd[110*NUM_OUTPUT_DATA+i],i_cmd[109*NUM_OUTPUT_DATA+i],i_cmd[108*NUM_OUTPUT_DATA+i],i_cmd[107*NUM_OUTPUT_DATA+i],i_cmd[106*NUM_OUTPUT_DATA+i],i_cmd[105*NUM_OUTPUT_DATA+i],i_cmd[104*NUM_OUTPUT_DATA+i],i_cmd[103*NUM_OUTPUT_DATA+i],i_cmd[102*NUM_OUTPUT_DATA+i],i_cmd[101*NUM_OUTPUT_DATA+i],i_cmd[100*NUM_OUTPUT_DATA+i],i_cmd[99*NUM_OUTPUT_DATA+i],i_cmd[98*NUM_OUTPUT_DATA+i],i_cmd[97*NUM_OUTPUT_DATA+i],i_cmd[96*NUM_OUTPUT_DATA+i],i_cmd[95*NUM_OUTPUT_DATA+i],i_cmd[94*NUM_OUTPUT_DATA+i],i_cmd[93*NUM_OUTPUT_DATA+i],i_cmd[92*NUM_OUTPUT_DATA+i],i_cmd[91*NUM_OUTPUT_DATA+i],i_cmd[90*NUM_OUTPUT_DATA+i],i_cmd[89*NUM_OUTPUT_DATA+i],i_cmd[88*NUM_OUTPUT_DATA+i],i_cmd[87*NUM_OUTPUT_DATA+i],i_cmd[86*NUM_OUTPUT_DATA+i],i_cmd[85*NUM_OUTPUT_DATA+i],i_cmd[84*NUM_OUTPUT_DATA+i],i_cmd[83*NUM_OUTPUT_DATA+i],i_cmd[82*NUM_OUTPUT_DATA+i],i_cmd[81*NUM_OUTPUT_DATA+i],i_cmd[80*NUM_OUTPUT_DATA+i],i_cmd[79*NUM_OUTPUT_DATA+i],i_cmd[78*NUM_OUTPUT_DATA+i],i_cmd[77*NUM_OUTPUT_DATA+i],i_cmd[76*NUM_OUTPUT_DATA+i],i_cmd[75*NUM_OUTPUT_DATA+i],i_cmd[74*NUM_OUTPUT_DATA+i],i_cmd[73*NUM_OUTPUT_DATA+i],i_cmd[72*NUM_OUTPUT_DATA+i],i_cmd[71*NUM_OUTPUT_DATA+i],i_cmd[70*NUM_OUTPUT_DATA+i],i_cmd[69*NUM_OUTPUT_DATA+i],i_cmd[68*NUM_OUTPUT_DATA+i],i_cmd[67*NUM_OUTPUT_DATA+i],i_cmd[66*NUM_OUTPUT_DATA+i],i_cmd[65*NUM_OUTPUT_DATA+i],i_cmd[64*NUM_OUTPUT_DATA+i],i_cmd[63*NUM_OUTPUT_DATA+i],i_cmd[62*NUM_OUTPUT_DATA+i],i_cmd[61*NUM_OUTPUT_DATA+i],i_cmd[60*NUM_OUTPUT_DATA+i],i_cmd[59*NUM_OUTPUT_DATA+i],i_cmd[58*NUM_OUTPUT_DATA+i],i_cmd[57*NUM_OUTPUT_DATA+i],i_cmd[56*NUM_OUTPUT_DATA+i],i_cmd[55*NUM_OUTPUT_DATA+i],i_cmd[54*NUM_OUTPUT_DATA+i],i_cmd[53*NUM_OUTPUT_DATA+i],i_cmd[52*NUM_OUTPUT_DATA+i],i_cmd[51*NUM_OUTPUT_DATA+i],i_cmd[50*NUM_OUTPUT_DATA+i],i_cmd[49*NUM_OUTPUT_DATA+i],i_cmd[48*NUM_OUTPUT_DATA+i],i_cmd[47*NUM_OUTPUT_DATA+i],i_cmd[46*NUM_OUTPUT_DATA+i],i_cmd[45*NUM_OUTPUT_DATA+i],i_cmd[44*NUM_OUTPUT_DATA+i],i_cmd[43*NUM_OUTPUT_DATA+i],i_cmd[42*NUM_OUTPUT_DATA+i],i_cmd[41*NUM_OUTPUT_DATA+i],i_cmd[40*NUM_OUTPUT_DATA+i],i_cmd[39*NUM_OUTPUT_DATA+i],i_cmd[38*NUM_OUTPUT_DATA+i],i_cmd[37*NUM_OUTPUT_DATA+i],i_cmd[36*NUM_OUTPUT_DATA+i],i_cmd[35*NUM_OUTPUT_DATA+i],i_cmd[34*NUM_OUTPUT_DATA+i],i_cmd[33*NUM_OUTPUT_DATA+i],i_cmd[32*NUM_OUTPUT_DATA+i],i_cmd[31*NUM_OUTPUT_DATA+i],i_cmd[30*NUM_OUTPUT_DATA+i],i_cmd[29*NUM_OUTPUT_DATA+i],i_cmd[28*NUM_OUTPUT_DATA+i],i_cmd[27*NUM_OUTPUT_DATA+i],i_cmd[26*NUM_OUTPUT_DATA+i],i_cmd[25*NUM_OUTPUT_DATA+i],i_cmd[24*NUM_OUTPUT_DATA+i],i_cmd[23*NUM_OUTPUT_DATA+i],i_cmd[22*NUM_OUTPUT_DATA+i],i_cmd[21*NUM_OUTPUT_DATA+i],i_cmd[20*NUM_OUTPUT_DATA+i],i_cmd[19*NUM_OUTPUT_DATA+i],i_cmd[18*NUM_OUTPUT_DATA+i],i_cmd[17*NUM_OUTPUT_DATA+i],i_cmd[16*NUM_OUTPUT_DATA+i],i_cmd[15*NUM_OUTPUT_DATA+i],i_cmd[14*NUM_OUTPUT_DATA+i],i_cmd[13*NUM_OUTPUT_DATA+i],i_cmd[12*NUM_OUTPUT_DATA+i],i_cmd[11*NUM_OUTPUT_DATA+i],i_cmd[10*NUM_OUTPUT_DATA+i],i_cmd[9*NUM_OUTPUT_DATA+i],i_cmd[8*NUM_OUTPUT_DATA+i],i_cmd[7*NUM_OUTPUT_DATA+i],i_cmd[6*NUM_OUTPUT_DATA+i],i_cmd[5*NUM_OUTPUT_DATA+i],i_cmd[4*NUM_OUTPUT_DATA+i],i_cmd[3*NUM_OUTPUT_DATA+i],i_cmd[2*NUM_OUTPUT_DATA+i],i_cmd[1*NUM_OUTPUT_DATA+i],i_cmd[0*NUM_OUTPUT_DATA+i]};
            always@(posedge CLK)
            begin
               if(i_en && (~rst))
                begin
                    case(inner_cmd_wire_valid)
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001:
                        begin
                            o_valid_reg[i] <= (i_valid[0])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010:
                        begin
                            o_valid_reg[i] <= (i_valid[1])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100:
                        begin
                            o_valid_reg[i] <= (i_valid[2])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000:
                        begin
                            o_valid_reg[i] <= (i_valid[3])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000:
                        begin
                            o_valid_reg[i] <= (i_valid[4])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000:
                        begin
                            o_valid_reg[i] <= (i_valid[5])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000:
                        begin
                            o_valid_reg[i] <= (i_valid[6])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000:
                        begin
                            o_valid_reg[i] <= (i_valid[7])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000:
                        begin
                            o_valid_reg[i] <= (i_valid[8])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[9])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[10])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[11])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[12])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[13])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[14])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[15])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[16])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[17])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[18])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[19])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[20])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[21])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[22])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[23])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[24])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[25])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[26])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[27])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[28])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[29])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[30])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[31])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[32])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[33])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[34])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[35])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[36])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[37])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[38])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[39])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[40])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[41])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[42])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[43])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[44])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[45])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[46])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[47])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[48])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[49])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[50])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[51])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[52])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[53])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[54])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[55])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[56])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[57])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[58])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[59])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[60])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[61])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[62])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[63])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[64])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[65])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[66])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[67])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[68])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[69])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[70])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[71])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[72])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[73])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[74])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[75])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[76])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[77])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[78])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[79])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[80])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[81])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[82])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[83])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[84])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[85])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[86])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[87])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[88])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[89])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[90])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[91])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[92])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[93])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[94])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[95])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[96])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[97])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[98])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[99])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[100])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[101])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[102])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[103])?1'b1:1'b0;
                        end
                        128'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[104])?1'b1:1'b0;
                        end
                        128'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[105])?1'b1:1'b0;
                        end
                        128'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[106])?1'b1:1'b0;
                        end
                        128'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[107])?1'b1:1'b0;
                        end
                        128'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[108])?1'b1:1'b0;
                        end
                        128'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[109])?1'b1:1'b0;
                        end
                        128'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[110])?1'b1:1'b0;
                        end
                        128'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[111])?1'b1:1'b0;
                        end
                        128'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[112])?1'b1:1'b0;
                        end
                        128'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[113])?1'b1:1'b0;
                        end
                        128'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[114])?1'b1:1'b0;
                        end
                        128'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[115])?1'b1:1'b0;
                        end
                        128'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[116])?1'b1:1'b0;
                        end
                        128'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[117])?1'b1:1'b0;
                        end
                        128'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[118])?1'b1:1'b0;
                        end
                        128'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[119])?1'b1:1'b0;
                        end
                        128'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[120])?1'b1:1'b0;
                        end
                        128'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[121])?1'b1:1'b0;
                        end
                        128'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[122])?1'b1:1'b0;
                        end
                        128'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[123])?1'b1:1'b0;
                        end
                        128'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[124])?1'b1:1'b0;
                        end
                        128'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[125])?1'b1:1'b0;
                        end
                        128'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[126])?1'b1:1'b0;
                        end
                        128'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
                        begin
                            o_valid_reg[i] <= (i_valid[127])?1'b1:1'b0;
                        end
                        default:
                        begin
                            o_valid_reg[i] <= 1'b0;
                        end
                    endcase
                end
                else
                begin
                    o_valid_reg[i] <= 1'b0;
                end
            end
        end
    endgenerate

    assign o_data_bus = o_data_bus_reg;
    assign o_valid = o_valid_reg;

endmodule
