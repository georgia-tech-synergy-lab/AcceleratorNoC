`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////////////////////
// Company: Gatech	
// Engineer: Mandovi Mukherjee
// 
// Create Date: 01/08/2021 
// System Name: accelerator
// Module Name: local controller
// Project Name: ARION DRBE
// Description: fetch and push data out to network; assuming the output from
// global controller comes in the form of a packet
// Dependencies:
// Additional Comments: 
/////////////////////////////////////////////////////////////////////////////////////////////////////

module local_controller_prefetch_full(CLK, reset, boot_up, start, input_boundary_flag, prev_dest_address, packet_out, boundary_next, dest_address, D, write_flag, from_glob_prefetch_valid, from_glob_prefetch_start, from_glob_prefetch_stop, from_glob_prefetch_dest,  write_boundary_next, input_write_boundary, prefetch_next_dest_addr, prefetch_next_stop_address, prefetch_boundary_prev, input_prefetch_boundary_flag, prefetch_stop_address, prefetch_dest_addr, scenario_update);

    // parameter
    	parameter N_sample = 256;
	parameter datawidth = 16;
	parameter address_vector_width = 4; //can be 200: 4 for tiny tapeout
	parameter id_width = 6; // 64 local controllers in subscaled system
	parameter sample_address_width = 8; /// assuming 1024 rows and 64 columns: needs to change if arrangement is different
	parameter packet_width = 2 + 2*datawidth + address_vector_width;  ///valid bit, real/prefetch flag, data, dest
	

//=== IO Ports ===//

     // Normal Mode Input
        input [31:0] D;
    	input CLK; // system clock, generated by VCO
	input reset;
	input boot_up;
	input start;
	
	input input_boundary_flag;
	input input_prefetch_boundary_flag;
	input input_write_boundary;
	input [address_vector_width - 1:0] prev_dest_address;
	input [address_vector_width - 1:0] prefetch_next_dest_addr;
        input [sample_address_width - 1:0] prefetch_next_stop_address;
	input [address_vector_width - 1:0] from_glob_prefetch_dest;
	
	

	input write_flag;

	input from_glob_prefetch_valid;
	input [sample_address_width - 1:0] from_glob_prefetch_start;
	input [sample_address_width - 1:0] from_glob_prefetch_stop;
	input scenario_update;

    // output
        output reg [packet_width-1:0] packet_out;   
        output reg boundary_next;
        output reg write_boundary_next;
        output reg [address_vector_width - 1:0] dest_address;
        output reg prefetch_boundary_prev;
	output reg [address_vector_width - 1:0] prefetch_dest_addr;
    	output reg [sample_address_width - 1:0] prefetch_stop_address;


//////////// internal status regs/signals //////////////////////////////////
    reg coeff_num;
    wire [2*datawidth - 1:0] data_from_sram;
    reg [2*datawidth - 1:0] packet_out_data;
    reg prefetch_reqd;
    reg [2*datawidth - 1:0] sram_D;
    wire WEBM;
    wire [31:0] DM;
    wire [31:0] BWEBM;


    wire BIST;
    wire AWT;
    wire SLP;
    wire SD;
    wire CEBM;
    reg [sample_address_width-1:0] A;	
    wire [sample_address_width-1:0] AM;
    reg sram_CEB;
    reg sram_WEB;
    reg [2*datawidth - 1:0] sram_BWEB;
    wire CLK_n;
    reg int_write_flag;
    reg internal_boundary_next;
    reg ready1;
    reg prefetch_ready1;
    reg prefetch_ready2;
    reg real_reqd;

    reg coeff_num_next;
    reg [sample_address_width - 1:0] next_scen_start_addr;
    reg scen_ready0;
    reg scen_ready1;
    reg [address_vector_width - 1:0] next_scen_prefetch_dest;

    reg prefetch_transfer;


///////////////////////////////////////////////////////////////////////////////    

////////// logic part ///////////////////////////////////////////////////////  

    assign AM = 0;
    assign WEBM = 1;
    assign CEBM = 1;
    assign BWEBM = 32'hffffffff;
    assign DM = 0;
    assign SLP = 0;
    assign SD = 0;
    assign AWT = 0;
    assign BIST = 0;
////////////sequential logic


   always @(posedge CLK_n) begin
	if (reset == 1 || scen_ready1 == 1) begin
		coeff_num_next <= 0;
		next_scen_start_addr <= 0;
		next_scen_prefetch_dest <= 0;
	end

	else if (boot_up == 0 && from_glob_prefetch_valid == 1) begin
		coeff_num_next <= 1;
		next_scen_start_addr <= from_glob_prefetch_start;
		next_scen_prefetch_dest <= from_glob_prefetch_dest;
	end
	else begin
		coeff_num_next <= coeff_num_next;
		next_scen_start_addr <= next_scen_start_addr;
		next_scen_prefetch_dest <= next_scen_prefetch_dest;
	end

   end



   always @(posedge CLK_n) begin
	if (reset == 1 || scenario_update == 1) begin
		prefetch_transfer = 0;
	end
	else if (input_prefetch_boundary_flag == 1) begin
		prefetch_transfer = 1;
	end
	else begin
		prefetch_transfer = prefetch_transfer;
	end
   end


   always @(posedge CLK_n) begin
	if (scenario_update) begin
     		scen_ready0 <= 1;
     		scen_ready1 <= 0;
	end
	else if (scen_ready0) begin
     		scen_ready0 <= 0;
     		scen_ready1 <= 1;
 	end
	else if (scen_ready1) begin
     		scen_ready0 <= 0;
     		scen_ready1 <= 0;
	end
	else    begin
     		scen_ready0 <= 0;
     		scen_ready1 <= 0;

	end

   end

   always @(posedge CLK_n) begin
	if (reset) begin
		packet_out <={1'b0,37'b0};
	end

 	else if (coeff_num == 1 && (scen_ready0 == 1 || scen_ready1 == 1 )) begin		// && write_flag == 0) begin
		packet_out <= {1'b1,1'b1,packet_out_data, dest_address};
	end
	else if (coeff_num == 1 && internal_boundary_next == 0) begin		// && write_flag == 0) begin
		packet_out <= {1'b1,1'b1,packet_out_data, dest_address};
	end
	else if (coeff_num == 1 && internal_boundary_next == 1) begin		// && write_flag == 0) begin
		packet_out <= {1'b1,1'b1,packet_out_data, dest_address};
	end
	else if (prefetch_ready2 == 1) begin
		packet_out <= {1'b1,1'b0,packet_out_data,prefetch_dest_addr};
	end
	else begin
		packet_out <= {1'b0,37'b0};
	end



   end



   always @(posedge CLK_n) begin
	if (reset) begin
		sram_CEB <= 1;
		sram_BWEB <= 32'hffffffff;
	end
	else if (write_flag == 1 || input_write_boundary == 1 || int_write_flag == 1) begin
		sram_CEB <= 0;
		sram_BWEB <= 32'h0;
	end

	else if (start == 1 || input_boundary_flag == 1) begin
		sram_CEB <= 0;
		sram_BWEB <= 32'hffffffff;
	end
        else if ( ready1 == 1 ) begin
		sram_CEB <= 0;
		sram_BWEB <= 32'hffffffff;
	end
	else if (coeff_num == 1 && internal_boundary_next == 0) begin
		if (coeff_num_next == 0 && scen_ready1 == 1) begin
			sram_CEB <= 1;
		end

		else begin
			sram_CEB <= 0;
		end
		sram_BWEB <= 32'hffffffff;
	end
	else if (coeff_num == 0) begin
		if (coeff_num_next == 1 && (scen_ready0 == 1 || scen_ready1 == 1 )) begin
			sram_CEB <= 0;
		end
		else if (input_boundary_flag == 0 && ready1 == 0  && int_write_flag==0 && input_write_boundary == 0 && prefetch_reqd == 1) begin
			if (prefetch_ready1 == 1) sram_CEB <= 0;
			else sram_CEB <= 0;
		end
		else begin
			sram_CEB <= 1;
		end
		sram_BWEB <= 32'hffffffff;
	end


	else begin 
		sram_CEB <= 1;
		sram_BWEB <= 32'hffffffff;
	end	

   end

  always @(posedge CLK_n) begin
	if (reset) begin
		A <= 8'h0;
	end
	else if (int_write_flag == 1) begin
		A <= A + 1;

	end

	else if (boot_up == 1 && from_glob_prefetch_valid == 1) begin
		A <= from_glob_prefetch_start;
	end
	else if (input_boundary_flag == 1) begin
		A <= A;
	end
	else if ( ready1 == 1 ) begin
		A <= A + 1;
	end

	else if (coeff_num == 1) begin
		if (scen_ready0 == 1) begin
			A <= next_scen_start_addr;
		end
		else if (internal_boundary_next == 1) begin
			A <= 8'h0;   //condition feasible??
		end
		else begin
			A <= A + 1;
		end
	end
	else if (coeff_num == 0 && (scen_ready0==1 || scen_ready1 == 1)) begin
		if (scen_ready0 == 1) begin
			A <= next_scen_start_addr;
		end
		else begin
			A <= A + 1;
		end
	end
	else if (coeff_num == 0 && (scen_ready0==0 && scen_ready1 == 0) && prefetch_reqd == 1) begin
		if (prefetch_ready1 == 0) begin
			if (prefetch_transfer == 1) begin
				A <= 8'hff;
			end
			else begin
				A <= next_scen_start_addr;
			end
		end
		else begin
			A <= A - 1;
		end
	end

	else begin
		A <= 8'h0;  
	end	

  end


    always @(posedge CLK_n) begin
	if (reset == 1 || write_boundary_next == 1)  begin
		int_write_flag <= 0;
		if (write_boundary_next == 1) begin
			sram_D <= D;
		end
		else begin
			sram_D <= 0;
		end

		sram_WEB <= 1;
		write_boundary_next <= 0;


	end

	else begin
		if (write_flag == 1 || input_write_boundary == 1) begin
			int_write_flag <= 1;
			sram_D <= D;
			sram_WEB <= 0;
			if (A == 8'hfe) begin
				write_boundary_next <= 1;

			end
			else begin
				write_boundary_next <= 0;

			end

		end
		else if (int_write_flag == 1) begin
			int_write_flag <= 1;
			sram_D <= D;
			sram_WEB <= 0;
			if (A == 8'hfe) begin
				write_boundary_next <= 1;

			end
			else if (A == 8'hff) begin
				write_boundary_next <= 0;

			end
			else begin
				write_boundary_next <= 0;

			end

		end

		else begin
			int_write_flag <= 0;
			sram_D <= 0;
			sram_WEB <= 1;
			write_boundary_next <= 0;

		end
	end

    end

    always @(posedge CLK_n) begin
	if (reset == 1 || scenario_update) begin
		real_reqd <= 0;
	end
	else if (boot_up == 1 && from_glob_prefetch_valid == 1) begin
		real_reqd <= 1;
	end
	else begin
		real_reqd <= real_reqd;
	end
    end

    always @ (posedge CLK_n) begin
        if (reset==1) begin
		dest_address <= 0;
		coeff_num <= 0;
		boundary_next <= 0;
		internal_boundary_next <= 0;
		ready1 <= 0;
		
        end
        else if (start==1) begin   /// start must go to 0 after 1 clock cycle
		dest_address <= dest_address;
		coeff_num <= coeff_num;
		boundary_next <= boundary_next;
		internal_boundary_next <= internal_boundary_next;
		if (real_reqd == 1) begin
			ready1 <= 1;
		end
		else begin
			ready1 <= 0;
		end
        end



        else if ((boot_up == 1 && from_glob_prefetch_valid == 1) || input_boundary_flag == 1) begin
		boundary_next <=0;
		internal_boundary_next <=0;
		if (boot_up == 1 && from_glob_prefetch_valid == 1) begin
			dest_address <= from_glob_prefetch_dest;
			ready1 <= 0;
		end
		else begin
			dest_address <= prev_dest_address;
			ready1 <= 1;
		end
		coeff_num <= 0;	
		//ready1 <= 1;
	end
        else if ( ready1 == 1 ) begin
		boundary_next <=0;
		internal_boundary_next <=0;
		dest_address <= dest_address;
		ready1 <= 0;
		coeff_num <= 1;	
	end

	else begin
		ready1 <= 0;
		if (coeff_num == 1 && scen_ready0 == 1) begin		// && write_flag == 0) begin
			boundary_next <= 0;
			internal_boundary_next <= 0;
			if (coeff_num_next == 1) begin
				dest_address <= dest_address;
				coeff_num <= 1;
			end
			else begin
				dest_address <= dest_address;
				coeff_num <= 1;
			end

		end
		else if (coeff_num == 1 && (scen_ready1 == 1)) begin 		// && write_flag == 0) begin
			boundary_next <= 0;
			internal_boundary_next <= 0;
			if (coeff_num_next == 1) begin
				dest_address <= next_scen_prefetch_dest;
				coeff_num <= 1;
			end
			else begin
				dest_address <= dest_address;
				coeff_num <= 0;
			end

		end

		else if (coeff_num == 1 && internal_boundary_next == 0) begin		// && write_flag == 0) begin
			dest_address <= dest_address;
			coeff_num <= coeff_num;
			if (A == 8'hfe) begin
				boundary_next <= 1;
				internal_boundary_next <= internal_boundary_next;
			end

			else if (A == 8'hff) begin
				boundary_next <= 0;//boundary_next;
				internal_boundary_next <= 1;
			end

			else begin
				boundary_next <= boundary_next;
				internal_boundary_next <= internal_boundary_next;
			end
		end
		else if (coeff_num == 1 && internal_boundary_next == 1) begin		// && write_flag == 0) begin
			dest_address <= dest_address;
			coeff_num <= 0;
			boundary_next <= boundary_next;
			internal_boundary_next <= 0;

		end
		else if (coeff_num == 0 && scen_ready0 == 1) begin		// && write_flag == 0) begin
			boundary_next <= 0;
			internal_boundary_next <= 0;
			if (coeff_num_next == 1) begin
				dest_address <= next_scen_prefetch_dest;
				coeff_num <= 0;
			end
			else begin
				dest_address <= 0;
				coeff_num <= 0;
			end

		end
		else if (coeff_num == 0 && scen_ready1 == 1) begin		// && write_flag == 0) begin
			boundary_next <= 0;
			internal_boundary_next <= 0;
			if (coeff_num_next == 1) begin
				dest_address <= dest_address;
				coeff_num <= 1;
			end
			else begin
				dest_address <= 0;
				coeff_num <= 0;
			end

		end
		else begin
			dest_address <= dest_address;
			coeff_num <= coeff_num;
			boundary_next <= boundary_next;
			internal_boundary_next <= internal_boundary_next;
		end

	end  
     end

     
       always @(posedge CLK_n) begin   
        if (reset == 1 || scenario_update == 1) begin
		prefetch_reqd <= 0;
		prefetch_dest_addr <= 0;
		prefetch_stop_address <= 0;
		prefetch_boundary_prev <= 0;
		prefetch_ready1 <= 0;
        end

	else if ((boot_up == 0 && from_glob_prefetch_valid == 1) || input_prefetch_boundary_flag == 1) begin
		prefetch_reqd <= 1;
		prefetch_boundary_prev <= 0;
		prefetch_ready1 <= 0;
		if (from_glob_prefetch_valid == 1) begin
			prefetch_dest_addr <= from_glob_prefetch_dest;
			prefetch_stop_address <= from_glob_prefetch_stop;
		end
		else begin
			prefetch_dest_addr <= prefetch_next_dest_addr;
			prefetch_stop_address <= prefetch_next_stop_address;
		end
	end

	else if (prefetch_boundary_prev == 1)  begin
		prefetch_dest_addr <= prefetch_dest_addr;
		prefetch_stop_address <= prefetch_stop_address;
		prefetch_reqd <= 0;
		prefetch_boundary_prev <= 0;   ////check condition
		prefetch_ready1 <= 0;
	end
	else if (coeff_num == 0 && input_boundary_flag == 0 && ready1 == 0  && int_write_flag==0 && input_write_boundary == 0 && prefetch_reqd == 1 ) begin
		prefetch_dest_addr <= prefetch_dest_addr;
		prefetch_stop_address <= prefetch_stop_address;
		if (prefetch_ready1 == 1) begin
			prefetch_boundary_prev <= prefetch_boundary_prev;   ////check condition
			if (A == prefetch_stop_address) begin
				prefetch_reqd <= 0;
				prefetch_boundary_prev <=0;
				prefetch_ready1 <= 0;
		
			end
			else if (A == 8'h0) begin
				prefetch_reqd <= 0;
				prefetch_boundary_prev <=1;
				prefetch_ready1 <= 0;

			end
			else begin
				prefetch_reqd <= prefetch_reqd;
				prefetch_boundary_prev <=prefetch_boundary_prev;
				prefetch_ready1 <= 1;
			end

		end

		else begin  ///check this branch
			prefetch_reqd <= prefetch_reqd; 
			prefetch_boundary_prev <= prefetch_boundary_prev;   ////check condition
			prefetch_ready1 <= 1;
		end
	

	end
	else begin
		prefetch_dest_addr <= prefetch_dest_addr;
		prefetch_reqd <= prefetch_reqd;
		prefetch_stop_address <= prefetch_stop_address;
		prefetch_boundary_prev <= prefetch_boundary_prev;
		prefetch_ready1 <= 0;
	end


     end

     always @(posedge CLK_n) begin
	if (reset == 1 || scenario_update == 1) begin
		prefetch_ready2 <= 0;
	end
	else if (prefetch_ready1 == 1) begin
		prefetch_ready2 <= 1;
	end
	else begin
		prefetch_ready2 <= 0;
	end
     end





     always @(posedge CLK) begin
	packet_out_data <= data_from_sram;

     end


    INVD6BWP30P140LVT UI_342 ( .I(CLK), .ZN(CLK_n) );

    TS1N28HPCPLVTB256X32M4SWBASO UI_dut_mem (.SLP(SLP), .SD(SD), .CLK(CLK), .CEB(sram_CEB), .WEB(sram_WEB), .CEBM(CEBM), .WEBM(WEBM), .AWT(AWT), .A(A[7:0]), .D(sram_D), .BWEB(sram_BWEB), .AM(AM), .DM(DM), .BWEBM(BWEBM), .BIST(BIST), .Q(data_from_sram));

	 
	 


   
endmodule
    
